
module iir_filter ( clk, rst_n, vIn, dIn, coeffs_fb, coeffs_ff, dOut, vOut );
  input [11:0] dIn;
  input [47:0] coeffs_fb;
  input [95:0] coeffs_ff;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   sw_regs_en_int, delayed_controls_0__1_, delayed_controls_1__0_,
         delayed_controls_1__1_, delayed_controls_2__0_, DP_n26, DP_n25,
         DP_n24, DP_n23, DP_n22, DP_n21, DP_n20, DP_n19, DP_n18, DP_n17,
         DP_n16, DP_n15, DP_n14, DP_n13, DP_n12, DP_n11, DP_n10, DP_n9, DP_n8,
         DP_n7, DP_n6, DP_n5, DP_n4, DP_n3, DP_n2, DP_n1, DP_fb_10_, DP_fb_11_,
         DP_fb_12_, DP_fb_13_, DP_fb_14_, DP_fb_15_, DP_fb_16_, DP_fb_17_,
         DP_fb_18_, DP_fb_19_, DP_fb_1_, DP_fb_20_, DP_fb_21_, DP_fb_22_,
         DP_fb_23_, DP_fb_2_, DP_fb_3_, DP_fb_4_, DP_fb_5_, DP_fb_6_, DP_fb_7_,
         DP_fb_8_, DP_fb_9_, DP_ff_0_, DP_ff_10_, DP_ff_11_, DP_ff_12_,
         DP_ff_13_, DP_ff_14_, DP_ff_15_, DP_ff_16_, DP_ff_17_, DP_ff_18_,
         DP_ff_19_, DP_ff_1_, DP_ff_20_, DP_ff_21_, DP_ff_22_, DP_ff_23_,
         DP_ff_2_, DP_ff_3_, DP_ff_4_, DP_ff_5_, DP_ff_6_, DP_ff_7_, DP_ff_8_,
         DP_ff_9_, DP_ff_part_0_, DP_ff_part_10_, DP_ff_part_11_,
         DP_ff_part_12_, DP_ff_part_13_, DP_ff_part_14_, DP_ff_part_15_,
         DP_ff_part_16_, DP_ff_part_17_, DP_ff_part_18_, DP_ff_part_19_,
         DP_ff_part_1_, DP_ff_part_20_, DP_ff_part_21_, DP_ff_part_22_,
         DP_ff_part_23_, DP_ff_part_2_, DP_ff_part_3_, DP_ff_part_4_,
         DP_ff_part_5_, DP_ff_part_6_, DP_ff_part_7_, DP_ff_part_8_,
         DP_ff_part_9_, DP_y_0_, DP_y_1_, DP_y_2_, DP_y_3_, DP_y_4_, DP_y_5_,
         DP_y_6_, DP_y_7_, DP_y_8_, DP_y_9_, DP_y_10_, DP_y_11_, DP_y_23,
         DP_sw1_0_, DP_sw1_1_, DP_sw1_2_, DP_sw1_3_, DP_sw1_4_, DP_sw1_5_,
         DP_sw1_6_, DP_sw1_7_, DP_sw1_8_, DP_sw1_9_, DP_sw1_10_, DP_sw1_11_,
         DP_sw1_12_, DP_sw1_13_, DP_sw1_14_, DP_sw1_15_, DP_sw1_16_,
         DP_sw1_17_, DP_sw1_18_, DP_sw1_19_, DP_sw1_20_, DP_sw1_21_,
         DP_sw1_22_, DP_sw1_23_, DP_sw0_0_, DP_sw0_1_, DP_sw0_2_, DP_sw0_3_,
         DP_sw0_4_, DP_sw0_5_, DP_sw0_6_, DP_sw0_7_, DP_sw0_8_, DP_sw0_9_,
         DP_sw0_10_, DP_sw0_11_, DP_sw0_12_, DP_sw0_13_, DP_sw0_14_,
         DP_sw0_15_, DP_sw0_16_, DP_sw0_17_, DP_sw0_18_, DP_sw0_19_,
         DP_sw0_20_, DP_sw0_21_, DP_sw0_22_, DP_sw0_23_, DP_w_0_, DP_w_1_,
         DP_w_2_, DP_w_3_, DP_w_4_, DP_w_5_, DP_w_6_, DP_w_7_, DP_w_8_,
         DP_w_9_, DP_w_10_, DP_w_11_, DP_w_12_, DP_w_13_, DP_w_14_, DP_w_15_,
         DP_w_16_, DP_w_17_, DP_w_18_, DP_w_19_, DP_w_20_, DP_w_21_, DP_w_22_,
         DP_w_23_, DP_x_0_, DP_x_1_, DP_x_2_, DP_x_3_, DP_x_4_, DP_x_5_,
         DP_x_6_, DP_x_7_, DP_x_8_, DP_x_9_, DP_x_10_, DP_x_11_, DP_reg_in_n13,
         DP_reg_in_n36, DP_reg_in_n35, DP_reg_in_n34, DP_reg_in_n33,
         DP_reg_in_n32, DP_reg_in_n31, DP_reg_in_n30, DP_reg_in_n29,
         DP_reg_in_n28, DP_reg_in_n27, DP_reg_in_n26, DP_reg_in_n25,
         DP_reg_coeff_fb_i_1_n73, DP_reg_coeff_fb_i_1_n39,
         DP_reg_coeff_fb_i_1_n28, DP_reg_coeff_fb_i_1_n26,
         DP_reg_coeff_fb_i_1_n25, DP_reg_coeff_fb_i_1_n23,
         DP_reg_coeff_fb_i_1_n21, DP_reg_coeff_fb_i_1_n18,
         DP_reg_coeff_fb_i_1_n16, DP_reg_coeff_fb_i_1_n15,
         DP_reg_coeff_fb_i_1_n14, DP_reg_coeff_fb_i_1_n13,
         DP_reg_coeff_fb_i_1_n3, DP_reg_coeff_fb_i_1_n1,
         DP_reg_coeff_fb_i_1_n72, DP_reg_coeff_fb_i_1_n71,
         DP_reg_coeff_fb_i_1_n70, DP_reg_coeff_fb_i_1_n69,
         DP_reg_coeff_fb_i_1_n68, DP_reg_coeff_fb_i_1_n67,
         DP_reg_coeff_fb_i_1_n66, DP_reg_coeff_fb_i_1_n65,
         DP_reg_coeff_fb_i_1_n64, DP_reg_coeff_fb_i_1_n63,
         DP_reg_coeff_fb_i_1_n62, DP_reg_coeff_fb_i_1_n61,
         DP_reg_coeff_fb_i_1_n60, DP_reg_coeff_fb_i_1_n59,
         DP_reg_coeff_fb_i_1_n58, DP_reg_coeff_fb_i_1_n57,
         DP_reg_coeff_fb_i_1_n56, DP_reg_coeff_fb_i_1_n55,
         DP_reg_coeff_fb_i_1_n54, DP_reg_coeff_fb_i_1_n53,
         DP_reg_coeff_fb_i_1_n52, DP_reg_coeff_fb_i_1_n51,
         DP_reg_coeff_fb_i_1_n50, DP_reg_coeff_fb_i_1_n49,
         DP_reg_coeff_fb_i_1_n48, DP_reg_coeff_fb_i_1_n47,
         DP_reg_coeff_fb_i_1_n46, DP_reg_coeff_fb_i_1_n45,
         DP_reg_coeff_fb_i_1_n44, DP_reg_coeff_fb_i_1_n43,
         DP_reg_coeff_fb_i_1_n42, DP_reg_coeff_fb_i_1_n41,
         DP_reg_coeff_fb_i_1_n40, DP_reg_coeff_fb_i_1_n38,
         DP_reg_coeff_fb_i_1_n37, DP_reg_coeff_fb_i_1_n36,
         DP_reg_coeff_fb_i_1_n34, DP_reg_coeff_fb_i_1_n32,
         DP_reg_coeff_fb_i_1_n31, DP_reg_coeff_fb_i_1_n29,
         DP_reg_coeff_fb_i_1_n83, DP_reg_coeff_fb_i_1_n82,
         DP_reg_coeff_fb_i_1_n81, DP_reg_coeff_fb_i_1_n80,
         DP_reg_coeff_fb_i_1_n79, DP_reg_coeff_fb_i_1_n78,
         DP_reg_coeff_fb_i_1_n77, DP_reg_coeff_fb_i_1_n76,
         DP_reg_coeff_fb_i_1_n75, DP_reg_coeff_fb_i_1_n74,
         DP_reg_coeff_fb_i_2_n124, DP_reg_coeff_fb_i_2_n123,
         DP_reg_coeff_fb_i_2_n122, DP_reg_coeff_fb_i_2_n121,
         DP_reg_coeff_fb_i_2_n120, DP_reg_coeff_fb_i_2_n119,
         DP_reg_coeff_fb_i_2_n118, DP_reg_coeff_fb_i_2_n117,
         DP_reg_coeff_fb_i_2_n116, DP_reg_coeff_fb_i_2_n115,
         DP_reg_coeff_fb_i_2_n114, DP_reg_coeff_fb_i_2_n113,
         DP_reg_coeff_fb_i_2_n112, DP_reg_coeff_fb_i_2_n111,
         DP_reg_coeff_fb_i_2_n110, DP_reg_coeff_fb_i_2_n109,
         DP_reg_coeff_fb_i_2_n108, DP_reg_coeff_fb_i_2_n107,
         DP_reg_coeff_fb_i_2_n106, DP_reg_coeff_fb_i_2_n105,
         DP_reg_coeff_fb_i_2_n104, DP_reg_coeff_fb_i_2_n103,
         DP_reg_coeff_fb_i_2_n102, DP_reg_coeff_fb_i_2_n101,
         DP_reg_coeff_fb_i_2_n100, DP_reg_coeff_fb_i_2_n99,
         DP_reg_coeff_fb_i_2_n98, DP_reg_coeff_fb_i_2_n97,
         DP_reg_coeff_fb_i_2_n96, DP_reg_coeff_fb_i_2_n95,
         DP_reg_coeff_fb_i_2_n94, DP_reg_coeff_fb_i_2_n93,
         DP_reg_coeff_fb_i_2_n92, DP_reg_coeff_fb_i_2_n91,
         DP_reg_coeff_fb_i_2_n90, DP_reg_coeff_fb_i_2_n89,
         DP_reg_coeff_fb_i_2_n88, DP_reg_coeff_fb_i_2_n87,
         DP_reg_coeff_fb_i_2_n86, DP_reg_coeff_fb_i_2_n85,
         DP_reg_coeff_fb_i_2_n84, DP_reg_coeff_fb_i_2_n83,
         DP_reg_coeff_fb_i_2_n82, DP_reg_coeff_fb_i_2_n81,
         DP_reg_coeff_fb_i_2_n80, DP_reg_coeff_fb_i_2_n79,
         DP_reg_coeff_fb_i_2_n78, DP_reg_coeff_fb_i_2_n77,
         DP_reg_coeff_fb_i_2_n76, DP_reg_coeff_fb_i_2_n75,
         DP_reg_coeff_fb_i_2_n73, DP_reg_coeff_fb_i_2_n42,
         DP_reg_coeff_fb_i_2_n28, DP_reg_coeff_fb_i_2_n24,
         DP_reg_coeff_fb_i_2_n22, DP_reg_coeff_fb_i_2_n21,
         DP_reg_coeff_fb_i_2_n20, DP_reg_coeff_fb_i_2_n19,
         DP_reg_coeff_fb_i_2_n18, DP_reg_coeff_fb_i_2_n17,
         DP_reg_coeff_fb_i_2_n16, DP_reg_coeff_fb_i_2_n15,
         DP_reg_coeff_fb_i_2_n14, DP_reg_coeff_fb_i_2_n12,
         DP_reg_coeff_fb_i_2_n11, DP_reg_coeff_fb_i_2_n10,
         DP_reg_coeff_fb_i_2_n9, DP_reg_coeff_fb_i_2_n8,
         DP_reg_coeff_fb_i_2_n7, DP_reg_coeff_fb_i_2_n126,
         DP_reg_coeff_fb_i_2_n125, DP_reg_b_i_0_n124, DP_reg_b_i_0_n123,
         DP_reg_b_i_0_n122, DP_reg_b_i_0_n121, DP_reg_b_i_0_n120,
         DP_reg_b_i_0_n119, DP_reg_b_i_0_n118, DP_reg_b_i_0_n117,
         DP_reg_b_i_0_n116, DP_reg_b_i_0_n115, DP_reg_b_i_0_n114,
         DP_reg_b_i_0_n113, DP_reg_b_i_0_n112, DP_reg_b_i_0_n111,
         DP_reg_b_i_0_n110, DP_reg_b_i_0_n109, DP_reg_b_i_0_n108,
         DP_reg_b_i_0_n107, DP_reg_b_i_0_n106, DP_reg_b_i_0_n105,
         DP_reg_b_i_0_n104, DP_reg_b_i_0_n103, DP_reg_b_i_0_n102,
         DP_reg_b_i_0_n101, DP_reg_b_i_0_n100, DP_reg_b_i_0_n99,
         DP_reg_b_i_0_n98, DP_reg_b_i_0_n97, DP_reg_b_i_0_n96,
         DP_reg_b_i_0_n95, DP_reg_b_i_0_n94, DP_reg_b_i_0_n93,
         DP_reg_b_i_0_n92, DP_reg_b_i_0_n91, DP_reg_b_i_0_n90,
         DP_reg_b_i_0_n89, DP_reg_b_i_0_n88, DP_reg_b_i_0_n87,
         DP_reg_b_i_0_n86, DP_reg_b_i_0_n85, DP_reg_b_i_0_n84,
         DP_reg_b_i_0_n83, DP_reg_b_i_0_n82, DP_reg_b_i_0_n81,
         DP_reg_b_i_0_n80, DP_reg_b_i_0_n79, DP_reg_b_i_0_n78,
         DP_reg_b_i_0_n77, DP_reg_b_i_0_n73, DP_reg_b_i_0_n28,
         DP_reg_b_i_0_n23, DP_reg_b_i_0_n22, DP_reg_b_i_0_n21,
         DP_reg_b_i_0_n19, DP_reg_b_i_0_n17, DP_reg_b_i_0_n15,
         DP_reg_b_i_0_n14, DP_reg_b_i_0_n13, DP_reg_b_i_0_n12,
         DP_reg_b_i_0_n11, DP_reg_b_i_0_n10, DP_reg_b_i_0_n9, DP_reg_b_i_0_n8,
         DP_reg_b_i_0_n7, DP_reg_b_i_0_n6, DP_reg_b_i_0_n5, DP_reg_b_i_0_n4,
         DP_reg_b_i_0_n3, DP_reg_b_i_0_n1, DP_reg_b_i_0_n131,
         DP_reg_b_i_0_n130, DP_reg_b_i_0_n129, DP_reg_b_i_0_n128,
         DP_reg_b_i_0_n127, DP_reg_b_i_0_n126, DP_reg_b_i_0_n125,
         DP_reg_b_i_1_n124, DP_reg_b_i_1_n123, DP_reg_b_i_1_n122,
         DP_reg_b_i_1_n121, DP_reg_b_i_1_n120, DP_reg_b_i_1_n119,
         DP_reg_b_i_1_n118, DP_reg_b_i_1_n117, DP_reg_b_i_1_n116,
         DP_reg_b_i_1_n115, DP_reg_b_i_1_n114, DP_reg_b_i_1_n113,
         DP_reg_b_i_1_n112, DP_reg_b_i_1_n111, DP_reg_b_i_1_n110,
         DP_reg_b_i_1_n109, DP_reg_b_i_1_n108, DP_reg_b_i_1_n107,
         DP_reg_b_i_1_n106, DP_reg_b_i_1_n105, DP_reg_b_i_1_n104,
         DP_reg_b_i_1_n103, DP_reg_b_i_1_n102, DP_reg_b_i_1_n101,
         DP_reg_b_i_1_n100, DP_reg_b_i_1_n99, DP_reg_b_i_1_n98,
         DP_reg_b_i_1_n97, DP_reg_b_i_1_n96, DP_reg_b_i_1_n95,
         DP_reg_b_i_1_n94, DP_reg_b_i_1_n93, DP_reg_b_i_1_n92,
         DP_reg_b_i_1_n91, DP_reg_b_i_1_n90, DP_reg_b_i_1_n89,
         DP_reg_b_i_1_n88, DP_reg_b_i_1_n87, DP_reg_b_i_1_n86,
         DP_reg_b_i_1_n85, DP_reg_b_i_1_n84, DP_reg_b_i_1_n83,
         DP_reg_b_i_1_n82, DP_reg_b_i_1_n81, DP_reg_b_i_1_n80,
         DP_reg_b_i_1_n79, DP_reg_b_i_1_n78, DP_reg_b_i_1_n77,
         DP_reg_b_i_1_n75, DP_reg_b_i_1_n74, DP_reg_b_i_1_n73,
         DP_reg_b_i_1_n42, DP_reg_b_i_1_n24, DP_reg_b_i_1_n23,
         DP_reg_b_i_1_n22, DP_reg_b_i_1_n20, DP_reg_b_i_1_n19,
         DP_reg_b_i_1_n18, DP_reg_b_i_1_n16, DP_reg_b_i_1_n15,
         DP_reg_b_i_1_n14, DP_reg_b_i_1_n13, DP_reg_b_i_1_n12,
         DP_reg_b_i_1_n11, DP_reg_b_i_1_n10, DP_reg_b_i_1_n9, DP_reg_b_i_1_n8,
         DP_reg_b_i_1_n7, DP_reg_b_i_1_n128, DP_reg_b_i_1_n127,
         DP_reg_b_i_1_n126, DP_reg_b_i_1_n125, DP_reg_b_i_2_n123,
         DP_reg_b_i_2_n122, DP_reg_b_i_2_n121, DP_reg_b_i_2_n120,
         DP_reg_b_i_2_n119, DP_reg_b_i_2_n118, DP_reg_b_i_2_n117,
         DP_reg_b_i_2_n116, DP_reg_b_i_2_n115, DP_reg_b_i_2_n114,
         DP_reg_b_i_2_n113, DP_reg_b_i_2_n112, DP_reg_b_i_2_n111,
         DP_reg_b_i_2_n110, DP_reg_b_i_2_n109, DP_reg_b_i_2_n108,
         DP_reg_b_i_2_n107, DP_reg_b_i_2_n106, DP_reg_b_i_2_n105,
         DP_reg_b_i_2_n104, DP_reg_b_i_2_n103, DP_reg_b_i_2_n102,
         DP_reg_b_i_2_n101, DP_reg_b_i_2_n100, DP_reg_b_i_2_n99,
         DP_reg_b_i_2_n98, DP_reg_b_i_2_n97, DP_reg_b_i_2_n96,
         DP_reg_b_i_2_n95, DP_reg_b_i_2_n94, DP_reg_b_i_2_n93,
         DP_reg_b_i_2_n92, DP_reg_b_i_2_n91, DP_reg_b_i_2_n90,
         DP_reg_b_i_2_n89, DP_reg_b_i_2_n88, DP_reg_b_i_2_n87,
         DP_reg_b_i_2_n86, DP_reg_b_i_2_n85, DP_reg_b_i_2_n84,
         DP_reg_b_i_2_n83, DP_reg_b_i_2_n82, DP_reg_b_i_2_n81,
         DP_reg_b_i_2_n80, DP_reg_b_i_2_n79, DP_reg_b_i_2_n78,
         DP_reg_b_i_2_n77, DP_reg_b_i_2_n76, DP_reg_b_i_2_n75,
         DP_reg_b_i_2_n74, DP_reg_b_i_2_n73, DP_reg_b_i_2_n44,
         DP_reg_b_i_2_n23, DP_reg_b_i_2_n22, DP_reg_b_i_2_n21,
         DP_reg_b_i_2_n19, DP_reg_b_i_2_n18, DP_reg_b_i_2_n17,
         DP_reg_b_i_2_n15, DP_reg_b_i_2_n13, DP_reg_b_i_2_n11, DP_reg_b_i_2_n9,
         DP_reg_b_i_2_n8, DP_reg_b_i_2_n7, DP_reg_b_i_2_n6, DP_reg_b_i_2_n5,
         DP_reg_b_i_2_n4, DP_reg_b_i_2_n3, DP_reg_b_i_2_n1, DP_reg_b_i_2_n130,
         DP_reg_b_i_2_n129, DP_reg_b_i_2_n128, DP_reg_b_i_2_n127,
         DP_reg_b_i_2_n126, DP_reg_b_i_2_n125, DP_reg_b_i_2_n124,
         DP_reg_b_i_3_n125, DP_reg_b_i_3_n124, DP_reg_b_i_3_n123,
         DP_reg_b_i_3_n122, DP_reg_b_i_3_n121, DP_reg_b_i_3_n120,
         DP_reg_b_i_3_n119, DP_reg_b_i_3_n118, DP_reg_b_i_3_n117,
         DP_reg_b_i_3_n116, DP_reg_b_i_3_n115, DP_reg_b_i_3_n114,
         DP_reg_b_i_3_n113, DP_reg_b_i_3_n112, DP_reg_b_i_3_n111,
         DP_reg_b_i_3_n110, DP_reg_b_i_3_n109, DP_reg_b_i_3_n108,
         DP_reg_b_i_3_n107, DP_reg_b_i_3_n106, DP_reg_b_i_3_n105,
         DP_reg_b_i_3_n104, DP_reg_b_i_3_n103, DP_reg_b_i_3_n102,
         DP_reg_b_i_3_n101, DP_reg_b_i_3_n100, DP_reg_b_i_3_n99,
         DP_reg_b_i_3_n98, DP_reg_b_i_3_n97, DP_reg_b_i_3_n96,
         DP_reg_b_i_3_n95, DP_reg_b_i_3_n94, DP_reg_b_i_3_n93,
         DP_reg_b_i_3_n92, DP_reg_b_i_3_n91, DP_reg_b_i_3_n90,
         DP_reg_b_i_3_n89, DP_reg_b_i_3_n88, DP_reg_b_i_3_n87,
         DP_reg_b_i_3_n86, DP_reg_b_i_3_n85, DP_reg_b_i_3_n84,
         DP_reg_b_i_3_n83, DP_reg_b_i_3_n82, DP_reg_b_i_3_n81,
         DP_reg_b_i_3_n80, DP_reg_b_i_3_n79, DP_reg_b_i_3_n78,
         DP_reg_b_i_3_n77, DP_reg_b_i_3_n73, DP_reg_b_i_3_n24,
         DP_reg_b_i_3_n23, DP_reg_b_i_3_n22, DP_reg_b_i_3_n20,
         DP_reg_b_i_3_n18, DP_reg_b_i_3_n16, DP_reg_b_i_3_n14,
         DP_reg_b_i_3_n12, DP_reg_b_i_3_n10, DP_reg_b_i_3_n9, DP_reg_b_i_3_n8,
         DP_reg_b_i_3_n7, DP_reg_b_i_3_n6, DP_reg_b_i_3_n5, DP_reg_b_i_3_n2,
         DP_reg_b_i_3_n1, DP_reg_b_i_3_n134, DP_reg_b_i_3_n133,
         DP_reg_b_i_3_n132, DP_reg_b_i_3_n131, DP_reg_b_i_3_n130,
         DP_reg_b_i_3_n129, DP_reg_b_i_3_n128, DP_reg_b_i_3_n127,
         DP_reg_b_i_3_n126, DP_reg_sw0_n87, DP_reg_sw0_n86, DP_reg_sw0_n85,
         DP_reg_sw0_n84, DP_reg_sw0_n83, DP_reg_sw0_n82, DP_reg_sw0_n81,
         DP_reg_sw0_n80, DP_reg_sw0_n79, DP_reg_sw0_n78, DP_reg_sw0_n77,
         DP_reg_sw0_n76, DP_reg_sw0_n75, DP_reg_sw0_n74, DP_reg_sw0_n73,
         DP_reg_sw0_n72, DP_reg_sw0_n71, DP_reg_sw0_n70, DP_reg_sw0_n69,
         DP_reg_sw0_n68, DP_reg_sw0_n67, DP_reg_sw0_n66, DP_reg_sw0_n65,
         DP_reg_sw0_n48, DP_reg_sw0_n47, DP_reg_sw0_n46, DP_reg_sw0_n45,
         DP_reg_sw0_n44, DP_reg_sw0_n43, DP_reg_sw0_n42, DP_reg_sw0_n41,
         DP_reg_sw0_n22, DP_reg_sw0_n21, DP_reg_sw0_n19, DP_reg_sw0_n17,
         DP_reg_sw0_n15, DP_reg_sw0_n14, DP_reg_sw0_n12, DP_reg_sw0_n10,
         DP_reg_sw0_n9, DP_reg_sw0_n8, DP_reg_sw0_n7, DP_reg_sw0_n6,
         DP_reg_sw0_n3, DP_reg_sw1_n114, DP_reg_sw1_n113, DP_reg_sw1_n112,
         DP_reg_sw1_n111, DP_reg_sw1_n110, DP_reg_sw1_n109, DP_reg_sw1_n108,
         DP_reg_sw1_n107, DP_reg_sw1_n106, DP_reg_sw1_n105, DP_reg_sw1_n104,
         DP_reg_sw1_n103, DP_reg_sw1_n102, DP_reg_sw1_n101, DP_reg_sw1_n100,
         DP_reg_sw1_n99, DP_reg_sw1_n98, DP_reg_sw1_n97, DP_reg_sw1_n96,
         DP_reg_sw1_n95, DP_reg_sw1_n94, DP_reg_sw1_n93, DP_reg_sw1_n92,
         DP_reg_sw1_n91, DP_reg_sw1_n90, DP_reg_sw1_n89, DP_reg_sw1_n88,
         DP_reg_sw1_n87, DP_reg_sw1_n86, DP_reg_sw1_n85, DP_reg_sw1_n84,
         DP_reg_sw1_n83, DP_reg_sw1_n82, DP_reg_sw1_n81, DP_reg_sw1_n80,
         DP_reg_sw1_n79, DP_reg_sw1_n78, DP_reg_sw1_n77, DP_reg_sw1_n76,
         DP_reg_sw1_n75, DP_reg_sw1_n74, DP_reg_sw1_n73, DP_reg_sw1_n45,
         DP_reg_sw1_n33, DP_reg_sw1_n31, DP_reg_sw1_n27, DP_reg_sw1_n25,
         DP_reg_sw1_n24, DP_reg_sw1_n23, DP_reg_sw1_n22, DP_reg_sw1_n21,
         DP_reg_sw1_n20, DP_reg_sw1_n19, DP_reg_sw1_n18, DP_reg_sw1_n17,
         DP_reg_sw1_n16, DP_reg_sw1_n14, DP_reg_sw1_n12, DP_reg_sw1_n10,
         DP_reg_sw1_n8, DP_reg_sw1_n7, DP_reg_sw1_n6, DP_reg_sw1_n5,
         DP_reg_sw1_n4, DP_reg_sw1_n3, DP_reg_sw1_n1, DP_reg_sw2_n52,
         DP_reg_sw2_n51, DP_reg_sw2_n48, DP_reg_sw2_n47, DP_reg_sw2_n46,
         DP_reg_sw2_n45, DP_reg_sw2_n44, DP_reg_sw2_n43, DP_reg_sw2_n42,
         DP_reg_sw2_n41, DP_reg_sw2_n40, DP_reg_sw2_n39, DP_reg_sw2_n38,
         DP_reg_sw2_n37, DP_reg_sw2_n36, DP_reg_sw2_n35, DP_reg_sw2_n34,
         DP_reg_sw2_n33, DP_reg_sw2_n32, DP_reg_sw2_n31, DP_reg_sw2_n30,
         DP_reg_sw2_n29, DP_reg_sw2_n28, DP_reg_sw2_n27, DP_reg_sw2_n26,
         DP_reg_sw2_n25, DP_reg_ret0_n100, DP_reg_ret0_n99, DP_reg_ret0_n98,
         DP_reg_ret0_n97, DP_reg_ret0_n96, DP_reg_ret0_n95, DP_reg_ret0_n94,
         DP_reg_ret0_n93, DP_reg_ret0_n92, DP_reg_ret0_n91, DP_reg_ret0_n90,
         DP_reg_ret0_n89, DP_reg_ret0_n88, DP_reg_ret0_n87, DP_reg_ret0_n86,
         DP_reg_ret0_n85, DP_reg_ret0_n84, DP_reg_ret0_n83, DP_reg_ret0_n82,
         DP_reg_ret0_n81, DP_reg_ret0_n80, DP_reg_ret0_n79, DP_reg_ret0_n78,
         DP_reg_ret0_n77, DP_reg_ret0_n76, DP_reg_ret0_n75, DP_reg_ret0_n73,
         DP_reg_ret0_n48, DP_reg_ret0_n47, DP_reg_ret0_n45, DP_reg_ret0_n44,
         DP_reg_ret0_n42, DP_reg_ret0_n41, DP_reg_ret0_n39, DP_reg_ret0_n38,
         DP_reg_ret0_n36, DP_reg_ret0_n35, DP_reg_ret0_n33, DP_reg_ret0_n32,
         DP_reg_ret0_n30, DP_reg_ret0_n29, DP_reg_ret0_n27, DP_reg_ret0_n26,
         DP_reg_ret0_n24, DP_reg_ret0_n23, DP_reg_ret0_n21, DP_reg_ret0_n20,
         DP_reg_ret0_n18, DP_reg_ret0_n17, DP_reg_ret0_n6, DP_reg_ret0_n5,
         DP_reg_ret1_n103, DP_reg_ret1_n102, DP_reg_ret1_n101,
         DP_reg_ret1_n100, DP_reg_ret1_n99, DP_reg_ret1_n98, DP_reg_ret1_n97,
         DP_reg_ret1_n96, DP_reg_ret1_n95, DP_reg_ret1_n94, DP_reg_ret1_n93,
         DP_reg_ret1_n92, DP_reg_ret1_n91, DP_reg_ret1_n90, DP_reg_ret1_n89,
         DP_reg_ret1_n88, DP_reg_ret1_n87, DP_reg_ret1_n86, DP_reg_ret1_n85,
         DP_reg_ret1_n84, DP_reg_ret1_n83, DP_reg_ret1_n82, DP_reg_ret1_n81,
         DP_reg_ret1_n80, DP_reg_ret1_n79, DP_reg_ret1_n78, DP_reg_ret1_n76,
         DP_reg_ret1_n75, DP_reg_ret1_n74, DP_reg_ret1_n48, DP_reg_ret1_n47,
         DP_reg_ret1_n45, DP_reg_ret1_n44, DP_reg_ret1_n42, DP_reg_ret1_n41,
         DP_reg_ret1_n39, DP_reg_ret1_n38, DP_reg_ret1_n36, DP_reg_ret1_n35,
         DP_reg_ret1_n33, DP_reg_ret1_n32, DP_reg_ret1_n30, DP_reg_ret1_n29,
         DP_reg_ret1_n27, DP_reg_ret1_n26, DP_reg_ret1_n24, DP_reg_ret1_n23,
         DP_reg_ret1_n21, DP_reg_ret1_n20, DP_reg_ret1_n6, DP_reg_ret1_n5,
         DP_reg_pipe00_n78, DP_reg_pipe00_n77, DP_reg_pipe00_n76,
         DP_reg_pipe00_n75, DP_reg_pipe00_n74, DP_reg_pipe00_n73,
         DP_reg_pipe00_n72, DP_reg_pipe00_n71, DP_reg_pipe00_n70,
         DP_reg_pipe00_n69, DP_reg_pipe00_n68, DP_reg_pipe00_n67,
         DP_reg_pipe00_n66, DP_reg_pipe00_n65, DP_reg_pipe00_n64,
         DP_reg_pipe00_n63, DP_reg_pipe00_n62, DP_reg_pipe00_n61,
         DP_reg_pipe00_n60, DP_reg_pipe00_n48, DP_reg_pipe00_n47,
         DP_reg_pipe00_n46, DP_reg_pipe00_n45, DP_reg_pipe00_n44,
         DP_reg_pipe00_n43, DP_reg_pipe00_n42, DP_reg_pipe00_n41,
         DP_reg_pipe00_n40, DP_reg_pipe00_n39, DP_reg_pipe00_n38,
         DP_reg_pipe00_n37, DP_reg_pipe00_n36, DP_reg_pipe00_n14,
         DP_reg_pipe00_n13, DP_reg_pipe00_n12, DP_reg_pipe00_n11,
         DP_reg_pipe00_n10, DP_reg_pipe00_n9, DP_reg_pipe00_n8,
         DP_reg_pipe00_n7, DP_reg_pipe00_n5, DP_reg_pipe00_n4,
         DP_reg_pipe01_n111, DP_reg_pipe01_n110, DP_reg_pipe01_n109,
         DP_reg_pipe01_n108, DP_reg_pipe01_n107, DP_reg_pipe01_n106,
         DP_reg_pipe01_n105, DP_reg_pipe01_n104, DP_reg_pipe01_n103,
         DP_reg_pipe01_n102, DP_reg_pipe01_n101, DP_reg_pipe01_n100,
         DP_reg_pipe01_n99, DP_reg_pipe01_n98, DP_reg_pipe01_n97,
         DP_reg_pipe01_n96, DP_reg_pipe01_n95, DP_reg_pipe01_n94,
         DP_reg_pipe01_n93, DP_reg_pipe01_n92, DP_reg_pipe01_n91,
         DP_reg_pipe01_n90, DP_reg_pipe01_n89, DP_reg_pipe01_n88,
         DP_reg_pipe01_n87, DP_reg_pipe01_n86, DP_reg_pipe01_n85,
         DP_reg_pipe01_n84, DP_reg_pipe01_n83, DP_reg_pipe01_n82,
         DP_reg_pipe01_n81, DP_reg_pipe01_n80, DP_reg_pipe01_n79,
         DP_reg_pipe01_n78, DP_reg_pipe01_n77, DP_reg_pipe01_n76,
         DP_reg_pipe01_n75, DP_reg_pipe01_n74, DP_reg_pipe01_n73,
         DP_reg_pipe01_n72, DP_reg_pipe01_n71, DP_reg_pipe01_n38,
         DP_reg_pipe01_n36, DP_reg_pipe01_n29, DP_reg_pipe01_n27,
         DP_reg_pipe01_n25, DP_reg_pipe01_n24, DP_reg_pipe01_n23,
         DP_reg_pipe01_n22, DP_reg_pipe01_n21, DP_reg_pipe01_n20,
         DP_reg_pipe01_n19, DP_reg_pipe01_n18, DP_reg_pipe01_n17,
         DP_reg_pipe01_n16, DP_reg_pipe01_n15, DP_reg_pipe01_n14,
         DP_reg_pipe01_n13, DP_reg_pipe01_n12, DP_reg_pipe01_n11,
         DP_reg_pipe01_n9, DP_reg_pipe01_n7, DP_reg_pipe01_n5,
         DP_reg_pipe01_n4, DP_reg_pipe02_n114, DP_reg_pipe02_n113,
         DP_reg_pipe02_n112, DP_reg_pipe02_n111, DP_reg_pipe02_n110,
         DP_reg_pipe02_n109, DP_reg_pipe02_n108, DP_reg_pipe02_n107,
         DP_reg_pipe02_n106, DP_reg_pipe02_n105, DP_reg_pipe02_n104,
         DP_reg_pipe02_n103, DP_reg_pipe02_n102, DP_reg_pipe02_n101,
         DP_reg_pipe02_n100, DP_reg_pipe02_n99, DP_reg_pipe02_n98,
         DP_reg_pipe02_n97, DP_reg_pipe02_n96, DP_reg_pipe02_n95,
         DP_reg_pipe02_n94, DP_reg_pipe02_n93, DP_reg_pipe02_n92,
         DP_reg_pipe02_n91, DP_reg_pipe02_n90, DP_reg_pipe02_n89,
         DP_reg_pipe02_n88, DP_reg_pipe02_n87, DP_reg_pipe02_n86,
         DP_reg_pipe02_n85, DP_reg_pipe02_n84, DP_reg_pipe02_n83,
         DP_reg_pipe02_n82, DP_reg_pipe02_n81, DP_reg_pipe02_n80,
         DP_reg_pipe02_n79, DP_reg_pipe02_n78, DP_reg_pipe02_n77,
         DP_reg_pipe02_n76, DP_reg_pipe02_n75, DP_reg_pipe02_n74,
         DP_reg_pipe02_n73, DP_reg_pipe02_n72, DP_reg_pipe02_n39,
         DP_reg_pipe02_n32, DP_reg_pipe02_n27, DP_reg_pipe02_n25,
         DP_reg_pipe02_n24, DP_reg_pipe02_n23, DP_reg_pipe02_n22,
         DP_reg_pipe02_n21, DP_reg_pipe02_n20, DP_reg_pipe02_n19,
         DP_reg_pipe02_n17, DP_reg_pipe02_n16, DP_reg_pipe02_n15,
         DP_reg_pipe02_n14, DP_reg_pipe02_n13, DP_reg_pipe02_n12,
         DP_reg_pipe02_n10, DP_reg_pipe02_n9, DP_reg_pipe02_n8,
         DP_reg_pipe02_n7, DP_reg_pipe02_n5, DP_reg_pipe02_n3,
         DP_reg_pipe02_n2, DP_reg_pipe03_n113, DP_reg_pipe03_n112,
         DP_reg_pipe03_n111, DP_reg_pipe03_n110, DP_reg_pipe03_n109,
         DP_reg_pipe03_n108, DP_reg_pipe03_n107, DP_reg_pipe03_n106,
         DP_reg_pipe03_n105, DP_reg_pipe03_n104, DP_reg_pipe03_n103,
         DP_reg_pipe03_n102, DP_reg_pipe03_n101, DP_reg_pipe03_n100,
         DP_reg_pipe03_n99, DP_reg_pipe03_n98, DP_reg_pipe03_n97,
         DP_reg_pipe03_n96, DP_reg_pipe03_n95, DP_reg_pipe03_n94,
         DP_reg_pipe03_n93, DP_reg_pipe03_n92, DP_reg_pipe03_n91,
         DP_reg_pipe03_n90, DP_reg_pipe03_n89, DP_reg_pipe03_n88,
         DP_reg_pipe03_n87, DP_reg_pipe03_n86, DP_reg_pipe03_n85,
         DP_reg_pipe03_n84, DP_reg_pipe03_n83, DP_reg_pipe03_n82,
         DP_reg_pipe03_n81, DP_reg_pipe03_n80, DP_reg_pipe03_n79,
         DP_reg_pipe03_n78, DP_reg_pipe03_n77, DP_reg_pipe03_n76,
         DP_reg_pipe03_n75, DP_reg_pipe03_n74, DP_reg_pipe03_n73,
         DP_reg_pipe03_n72, DP_reg_pipe03_n39, DP_reg_pipe03_n34,
         DP_reg_pipe03_n33, DP_reg_pipe03_n27, DP_reg_pipe03_n25,
         DP_reg_pipe03_n24, DP_reg_pipe03_n23, DP_reg_pipe03_n22,
         DP_reg_pipe03_n21, DP_reg_pipe03_n20, DP_reg_pipe03_n18,
         DP_reg_pipe03_n17, DP_reg_pipe03_n16, DP_reg_pipe03_n15,
         DP_reg_pipe03_n12, DP_reg_pipe03_n11, DP_reg_pipe03_n10,
         DP_reg_pipe03_n9, DP_reg_pipe03_n8, DP_reg_pipe03_n6,
         DP_reg_pipe03_n5, DP_reg_pipe03_n4, DP_reg_pipe03_n3,
         DP_reg_pipe03_n1, DP_reg_pipe10_n107, DP_reg_pipe10_n106,
         DP_reg_pipe10_n105, DP_reg_pipe10_n104, DP_reg_pipe10_n103,
         DP_reg_pipe10_n102, DP_reg_pipe10_n101, DP_reg_pipe10_n100,
         DP_reg_pipe10_n99, DP_reg_pipe10_n98, DP_reg_pipe10_n97,
         DP_reg_pipe10_n96, DP_reg_pipe10_n95, DP_reg_pipe10_n94,
         DP_reg_pipe10_n93, DP_reg_pipe10_n92, DP_reg_pipe10_n91,
         DP_reg_pipe10_n90, DP_reg_pipe10_n89, DP_reg_pipe10_n88,
         DP_reg_pipe10_n87, DP_reg_pipe10_n86, DP_reg_pipe10_n85,
         DP_reg_pipe10_n84, DP_reg_pipe10_n82, DP_reg_pipe10_n81,
         DP_reg_pipe10_n79, DP_reg_pipe10_n78, DP_reg_pipe10_n77,
         DP_reg_pipe10_n75, DP_reg_pipe10_n74, DP_reg_pipe10_n48,
         DP_reg_pipe10_n47, DP_reg_pipe10_n45, DP_reg_pipe10_n44,
         DP_reg_pipe10_n42, DP_reg_pipe10_n41, DP_reg_pipe10_n39,
         DP_reg_pipe10_n38, DP_reg_pipe10_n36, DP_reg_pipe10_n35,
         DP_reg_pipe10_n33, DP_reg_pipe10_n32, DP_reg_pipe10_n30,
         DP_reg_pipe10_n29, DP_reg_pipe10_n27, DP_reg_pipe10_n26,
         DP_reg_pipe10_n13, DP_reg_pipe10_n12, DP_reg_pipe11_n97,
         DP_reg_pipe11_n96, DP_reg_pipe11_n95, DP_reg_pipe11_n94,
         DP_reg_pipe11_n93, DP_reg_pipe11_n92, DP_reg_pipe11_n91,
         DP_reg_pipe11_n90, DP_reg_pipe11_n89, DP_reg_pipe11_n88,
         DP_reg_pipe11_n87, DP_reg_pipe11_n86, DP_reg_pipe11_n85,
         DP_reg_pipe11_n84, DP_reg_pipe11_n83, DP_reg_pipe11_n82,
         DP_reg_pipe11_n81, DP_reg_pipe11_n80, DP_reg_pipe11_n79,
         DP_reg_pipe11_n78, DP_reg_pipe11_n77, DP_reg_pipe11_n76,
         DP_reg_pipe11_n75, DP_reg_pipe11_n74, DP_reg_pipe11_n73,
         DP_reg_pipe11_n48, DP_reg_pipe11_n47, DP_reg_pipe11_n46,
         DP_reg_pipe11_n45, DP_reg_pipe11_n44, DP_reg_pipe11_n43,
         DP_reg_pipe11_n42, DP_reg_pipe11_n41, DP_reg_pipe11_n40,
         DP_reg_pipe11_n39, DP_reg_pipe11_n38, DP_reg_pipe11_n37,
         DP_reg_pipe11_n36, DP_reg_pipe11_n35, DP_reg_pipe11_n34,
         DP_reg_pipe11_n33, DP_reg_pipe11_n32, DP_reg_pipe11_n31,
         DP_reg_pipe11_n30, DP_reg_pipe11_n29, DP_reg_pipe11_n28,
         DP_reg_pipe11_n27, DP_reg_pipe11_n26, DP_reg_pipe11_n3,
         DP_reg_pipe12_n101, DP_reg_pipe12_n100, DP_reg_pipe12_n99,
         DP_reg_pipe12_n98, DP_reg_pipe12_n97, DP_reg_pipe12_n96,
         DP_reg_pipe12_n95, DP_reg_pipe12_n94, DP_reg_pipe12_n93,
         DP_reg_pipe12_n92, DP_reg_pipe12_n91, DP_reg_pipe12_n90,
         DP_reg_pipe12_n89, DP_reg_pipe12_n88, DP_reg_pipe12_n87,
         DP_reg_pipe12_n86, DP_reg_pipe12_n85, DP_reg_pipe12_n84,
         DP_reg_pipe12_n83, DP_reg_pipe12_n82, DP_reg_pipe12_n81,
         DP_reg_pipe12_n80, DP_reg_pipe12_n79, DP_reg_pipe12_n78,
         DP_reg_pipe12_n76, DP_reg_pipe12_n75, DP_reg_pipe12_n73,
         DP_reg_pipe12_n48, DP_reg_pipe12_n47, DP_reg_pipe12_n45,
         DP_reg_pipe12_n44, DP_reg_pipe12_n42, DP_reg_pipe12_n41,
         DP_reg_pipe12_n39, DP_reg_pipe12_n38, DP_reg_pipe12_n36,
         DP_reg_pipe12_n35, DP_reg_pipe12_n33, DP_reg_pipe12_n32,
         DP_reg_pipe12_n30, DP_reg_pipe12_n29, DP_reg_pipe12_n27,
         DP_reg_pipe12_n26, DP_reg_pipe12_n24, DP_reg_pipe12_n23,
         DP_reg_pipe12_n21, DP_reg_pipe12_n20, DP_reg_pipe12_n8,
         DP_reg_pipe12_n7, DP_reg_pipe13_n106, DP_reg_pipe13_n105,
         DP_reg_pipe13_n104, DP_reg_pipe13_n103, DP_reg_pipe13_n102,
         DP_reg_pipe13_n101, DP_reg_pipe13_n100, DP_reg_pipe13_n99,
         DP_reg_pipe13_n98, DP_reg_pipe13_n97, DP_reg_pipe13_n96,
         DP_reg_pipe13_n95, DP_reg_pipe13_n94, DP_reg_pipe13_n93,
         DP_reg_pipe13_n92, DP_reg_pipe13_n91, DP_reg_pipe13_n90,
         DP_reg_pipe13_n89, DP_reg_pipe13_n88, DP_reg_pipe13_n87,
         DP_reg_pipe13_n86, DP_reg_pipe13_n85, DP_reg_pipe13_n84,
         DP_reg_pipe13_n83, DP_reg_pipe13_n81, DP_reg_pipe13_n80,
         DP_reg_pipe13_n78, DP_reg_pipe13_n77, DP_reg_pipe13_n76,
         DP_reg_pipe13_n74, DP_reg_pipe13_n73, DP_reg_pipe13_n47,
         DP_reg_pipe13_n46, DP_reg_pipe13_n44, DP_reg_pipe13_n43,
         DP_reg_pipe13_n41, DP_reg_pipe13_n40, DP_reg_pipe13_n38,
         DP_reg_pipe13_n37, DP_reg_pipe13_n35, DP_reg_pipe13_n34,
         DP_reg_pipe13_n32, DP_reg_pipe13_n31, DP_reg_pipe13_n29,
         DP_reg_pipe13_n28, DP_reg_pipe13_n26, DP_reg_pipe13_n25,
         DP_reg_pipe13_n14, DP_reg_pipe13_n13, DP_reg_out_n26, DP_reg_out_n24,
         DP_reg_out_n23, DP_reg_out_n22, DP_reg_out_n21, DP_reg_out_n20,
         DP_reg_out_n19, DP_reg_out_n18, DP_reg_out_n17, DP_reg_out_n16,
         DP_reg_out_n15, DP_reg_out_n14, DP_reg_out_n1,
         DP_add_2_root_add_0_root_add_223_n296,
         DP_add_2_root_add_0_root_add_223_n295,
         DP_add_2_root_add_0_root_add_223_n294,
         DP_add_2_root_add_0_root_add_223_n213,
         DP_add_2_root_add_0_root_add_223_n212,
         DP_add_2_root_add_0_root_add_223_n211,
         DP_add_2_root_add_0_root_add_223_n209,
         DP_add_2_root_add_0_root_add_223_n208,
         DP_add_2_root_add_0_root_add_223_n207,
         DP_add_2_root_add_0_root_add_223_n206,
         DP_add_2_root_add_0_root_add_223_n205,
         DP_add_2_root_add_0_root_add_223_n203,
         DP_add_2_root_add_0_root_add_223_n201,
         DP_add_2_root_add_0_root_add_223_n199,
         DP_add_2_root_add_0_root_add_223_n198,
         DP_add_2_root_add_0_root_add_223_n197,
         DP_add_2_root_add_0_root_add_223_n195,
         DP_add_2_root_add_0_root_add_223_n193,
         DP_add_2_root_add_0_root_add_223_n192,
         DP_add_2_root_add_0_root_add_223_n190,
         DP_add_2_root_add_0_root_add_223_n188,
         DP_add_2_root_add_0_root_add_223_n187,
         DP_add_2_root_add_0_root_add_223_n186,
         DP_add_2_root_add_0_root_add_223_n185,
         DP_add_2_root_add_0_root_add_223_n184,
         DP_add_2_root_add_0_root_add_223_n183,
         DP_add_2_root_add_0_root_add_223_n182,
         DP_add_2_root_add_0_root_add_223_n181,
         DP_add_2_root_add_0_root_add_223_n180,
         DP_add_2_root_add_0_root_add_223_n179,
         DP_add_2_root_add_0_root_add_223_n178,
         DP_add_2_root_add_0_root_add_223_n177,
         DP_add_2_root_add_0_root_add_223_n176,
         DP_add_2_root_add_0_root_add_223_n175,
         DP_add_2_root_add_0_root_add_223_n174,
         DP_add_2_root_add_0_root_add_223_n173,
         DP_add_2_root_add_0_root_add_223_n172,
         DP_add_2_root_add_0_root_add_223_n171,
         DP_add_2_root_add_0_root_add_223_n170,
         DP_add_2_root_add_0_root_add_223_n169,
         DP_add_2_root_add_0_root_add_223_n168,
         DP_add_2_root_add_0_root_add_223_n167,
         DP_add_2_root_add_0_root_add_223_n166,
         DP_add_2_root_add_0_root_add_223_n165,
         DP_add_2_root_add_0_root_add_223_n164,
         DP_add_2_root_add_0_root_add_223_n163,
         DP_add_2_root_add_0_root_add_223_n162,
         DP_add_2_root_add_0_root_add_223_n161,
         DP_add_2_root_add_0_root_add_223_n160,
         DP_add_2_root_add_0_root_add_223_n159,
         DP_add_2_root_add_0_root_add_223_n158,
         DP_add_2_root_add_0_root_add_223_n157,
         DP_add_2_root_add_0_root_add_223_n156,
         DP_add_2_root_add_0_root_add_223_n155,
         DP_add_2_root_add_0_root_add_223_n154,
         DP_add_2_root_add_0_root_add_223_n153,
         DP_add_2_root_add_0_root_add_223_n152,
         DP_add_2_root_add_0_root_add_223_n151,
         DP_add_2_root_add_0_root_add_223_n150,
         DP_add_2_root_add_0_root_add_223_n149,
         DP_add_2_root_add_0_root_add_223_n148,
         DP_add_2_root_add_0_root_add_223_n147,
         DP_add_2_root_add_0_root_add_223_n145,
         DP_add_2_root_add_0_root_add_223_n143,
         DP_add_2_root_add_0_root_add_223_n142,
         DP_add_2_root_add_0_root_add_223_n141,
         DP_add_2_root_add_0_root_add_223_n140,
         DP_add_2_root_add_0_root_add_223_n139,
         DP_add_2_root_add_0_root_add_223_n138,
         DP_add_2_root_add_0_root_add_223_n137,
         DP_add_2_root_add_0_root_add_223_n136,
         DP_add_2_root_add_0_root_add_223_n135,
         DP_add_2_root_add_0_root_add_223_n134,
         DP_add_2_root_add_0_root_add_223_n133,
         DP_add_2_root_add_0_root_add_223_n132,
         DP_add_2_root_add_0_root_add_223_n131,
         DP_add_2_root_add_0_root_add_223_n130,
         DP_add_2_root_add_0_root_add_223_n129,
         DP_add_2_root_add_0_root_add_223_n128,
         DP_add_2_root_add_0_root_add_223_n127,
         DP_add_2_root_add_0_root_add_223_n126,
         DP_add_2_root_add_0_root_add_223_n125,
         DP_add_2_root_add_0_root_add_223_n124,
         DP_add_2_root_add_0_root_add_223_n123,
         DP_add_2_root_add_0_root_add_223_n122,
         DP_add_2_root_add_0_root_add_223_n121,
         DP_add_2_root_add_0_root_add_223_n120,
         DP_add_2_root_add_0_root_add_223_n119,
         DP_add_2_root_add_0_root_add_223_n118,
         DP_add_2_root_add_0_root_add_223_n117,
         DP_add_2_root_add_0_root_add_223_n116,
         DP_add_2_root_add_0_root_add_223_n115,
         DP_add_2_root_add_0_root_add_223_n114,
         DP_add_2_root_add_0_root_add_223_n113,
         DP_add_2_root_add_0_root_add_223_n112,
         DP_add_2_root_add_0_root_add_223_n111,
         DP_add_2_root_add_0_root_add_223_n110,
         DP_add_2_root_add_0_root_add_223_n109,
         DP_add_2_root_add_0_root_add_223_n108,
         DP_add_2_root_add_0_root_add_223_n107,
         DP_add_2_root_add_0_root_add_223_n106,
         DP_add_2_root_add_0_root_add_223_n105,
         DP_add_2_root_add_0_root_add_223_n104,
         DP_add_2_root_add_0_root_add_223_n103,
         DP_add_2_root_add_0_root_add_223_n102,
         DP_add_2_root_add_0_root_add_223_n101,
         DP_add_2_root_add_0_root_add_223_n100,
         DP_add_2_root_add_0_root_add_223_n99,
         DP_add_2_root_add_0_root_add_223_n98,
         DP_add_2_root_add_0_root_add_223_n97,
         DP_add_2_root_add_0_root_add_223_n96,
         DP_add_2_root_add_0_root_add_223_n95,
         DP_add_2_root_add_0_root_add_223_n94,
         DP_add_2_root_add_0_root_add_223_n93,
         DP_add_2_root_add_0_root_add_223_n92,
         DP_add_2_root_add_0_root_add_223_n91,
         DP_add_2_root_add_0_root_add_223_n90,
         DP_add_2_root_add_0_root_add_223_n89,
         DP_add_2_root_add_0_root_add_223_n88,
         DP_add_2_root_add_0_root_add_223_n87,
         DP_add_2_root_add_0_root_add_223_n86,
         DP_add_2_root_add_0_root_add_223_n85,
         DP_add_2_root_add_0_root_add_223_n84,
         DP_add_2_root_add_0_root_add_223_n83,
         DP_add_2_root_add_0_root_add_223_n82,
         DP_add_2_root_add_0_root_add_223_n81,
         DP_add_2_root_add_0_root_add_223_n80,
         DP_add_2_root_add_0_root_add_223_n79,
         DP_add_2_root_add_0_root_add_223_n78,
         DP_add_2_root_add_0_root_add_223_n77,
         DP_add_2_root_add_0_root_add_223_n76,
         DP_add_2_root_add_0_root_add_223_n75,
         DP_add_2_root_add_0_root_add_223_n74,
         DP_add_2_root_add_0_root_add_223_n73,
         DP_add_2_root_add_0_root_add_223_n72,
         DP_add_2_root_add_0_root_add_223_n71,
         DP_add_2_root_add_0_root_add_223_n70,
         DP_add_2_root_add_0_root_add_223_n69,
         DP_add_2_root_add_0_root_add_223_n68,
         DP_add_2_root_add_0_root_add_223_n67,
         DP_add_2_root_add_0_root_add_223_n66,
         DP_add_2_root_add_0_root_add_223_n65,
         DP_add_2_root_add_0_root_add_223_n64,
         DP_add_2_root_add_0_root_add_223_n63,
         DP_add_2_root_add_0_root_add_223_n62,
         DP_add_2_root_add_0_root_add_223_n61,
         DP_add_2_root_add_0_root_add_223_n60,
         DP_add_2_root_add_0_root_add_223_n59,
         DP_add_2_root_add_0_root_add_223_n58,
         DP_add_2_root_add_0_root_add_223_n57,
         DP_add_2_root_add_0_root_add_223_n56,
         DP_add_2_root_add_0_root_add_223_n55,
         DP_add_2_root_add_0_root_add_223_n54,
         DP_add_2_root_add_0_root_add_223_n53,
         DP_add_2_root_add_0_root_add_223_n52,
         DP_add_2_root_add_0_root_add_223_n51,
         DP_add_2_root_add_0_root_add_223_n50,
         DP_add_2_root_add_0_root_add_223_n49,
         DP_add_2_root_add_0_root_add_223_n48,
         DP_add_2_root_add_0_root_add_223_n47,
         DP_add_2_root_add_0_root_add_223_n46,
         DP_add_2_root_add_0_root_add_223_n45,
         DP_add_2_root_add_0_root_add_223_n44,
         DP_add_2_root_add_0_root_add_223_n43,
         DP_add_2_root_add_0_root_add_223_n42,
         DP_add_2_root_add_0_root_add_223_n41,
         DP_add_2_root_add_0_root_add_223_n40,
         DP_add_2_root_add_0_root_add_223_n39,
         DP_add_2_root_add_0_root_add_223_n38,
         DP_add_2_root_add_0_root_add_223_n37,
         DP_add_2_root_add_0_root_add_223_n36,
         DP_add_2_root_add_0_root_add_223_n35,
         DP_add_2_root_add_0_root_add_223_n34,
         DP_add_2_root_add_0_root_add_223_n33,
         DP_add_2_root_add_0_root_add_223_n32,
         DP_add_2_root_add_0_root_add_223_n30,
         DP_add_2_root_add_0_root_add_223_n28,
         DP_add_2_root_add_0_root_add_223_n27,
         DP_add_2_root_add_0_root_add_223_n24,
         DP_add_2_root_add_0_root_add_223_n23,
         DP_add_2_root_add_0_root_add_223_n22,
         DP_add_2_root_add_0_root_add_223_n21,
         DP_add_2_root_add_0_root_add_223_n20,
         DP_add_2_root_add_0_root_add_223_n19,
         DP_add_2_root_add_0_root_add_223_n18,
         DP_add_2_root_add_0_root_add_223_n17,
         DP_add_2_root_add_0_root_add_223_n16,
         DP_add_2_root_add_0_root_add_223_n15,
         DP_add_2_root_add_0_root_add_223_n14,
         DP_add_2_root_add_0_root_add_223_n13,
         DP_add_2_root_add_0_root_add_223_n12,
         DP_add_2_root_add_0_root_add_223_n11,
         DP_add_2_root_add_0_root_add_223_n10,
         DP_add_2_root_add_0_root_add_223_n9,
         DP_add_2_root_add_0_root_add_223_n8,
         DP_add_2_root_add_0_root_add_223_n7,
         DP_add_2_root_add_0_root_add_223_n6,
         DP_add_2_root_add_0_root_add_223_n5,
         DP_add_2_root_add_0_root_add_223_n4,
         DP_add_2_root_add_0_root_add_223_n3,
         DP_add_2_root_add_0_root_add_223_n2,
         DP_add_2_root_add_0_root_add_223_n1,
         DP_add_1_root_add_0_root_add_223_n296,
         DP_add_1_root_add_0_root_add_223_n295,
         DP_add_1_root_add_0_root_add_223_n294,
         DP_add_1_root_add_0_root_add_223_n213,
         DP_add_1_root_add_0_root_add_223_n212,
         DP_add_1_root_add_0_root_add_223_n211,
         DP_add_1_root_add_0_root_add_223_n209,
         DP_add_1_root_add_0_root_add_223_n208,
         DP_add_1_root_add_0_root_add_223_n207,
         DP_add_1_root_add_0_root_add_223_n206,
         DP_add_1_root_add_0_root_add_223_n205,
         DP_add_1_root_add_0_root_add_223_n203,
         DP_add_1_root_add_0_root_add_223_n201,
         DP_add_1_root_add_0_root_add_223_n199,
         DP_add_1_root_add_0_root_add_223_n198,
         DP_add_1_root_add_0_root_add_223_n197,
         DP_add_1_root_add_0_root_add_223_n195,
         DP_add_1_root_add_0_root_add_223_n193,
         DP_add_1_root_add_0_root_add_223_n192,
         DP_add_1_root_add_0_root_add_223_n190,
         DP_add_1_root_add_0_root_add_223_n188,
         DP_add_1_root_add_0_root_add_223_n187,
         DP_add_1_root_add_0_root_add_223_n186,
         DP_add_1_root_add_0_root_add_223_n185,
         DP_add_1_root_add_0_root_add_223_n184,
         DP_add_1_root_add_0_root_add_223_n183,
         DP_add_1_root_add_0_root_add_223_n182,
         DP_add_1_root_add_0_root_add_223_n181,
         DP_add_1_root_add_0_root_add_223_n180,
         DP_add_1_root_add_0_root_add_223_n179,
         DP_add_1_root_add_0_root_add_223_n178,
         DP_add_1_root_add_0_root_add_223_n177,
         DP_add_1_root_add_0_root_add_223_n176,
         DP_add_1_root_add_0_root_add_223_n175,
         DP_add_1_root_add_0_root_add_223_n174,
         DP_add_1_root_add_0_root_add_223_n173,
         DP_add_1_root_add_0_root_add_223_n172,
         DP_add_1_root_add_0_root_add_223_n171,
         DP_add_1_root_add_0_root_add_223_n170,
         DP_add_1_root_add_0_root_add_223_n169,
         DP_add_1_root_add_0_root_add_223_n168,
         DP_add_1_root_add_0_root_add_223_n167,
         DP_add_1_root_add_0_root_add_223_n166,
         DP_add_1_root_add_0_root_add_223_n165,
         DP_add_1_root_add_0_root_add_223_n164,
         DP_add_1_root_add_0_root_add_223_n163,
         DP_add_1_root_add_0_root_add_223_n162,
         DP_add_1_root_add_0_root_add_223_n161,
         DP_add_1_root_add_0_root_add_223_n160,
         DP_add_1_root_add_0_root_add_223_n159,
         DP_add_1_root_add_0_root_add_223_n158,
         DP_add_1_root_add_0_root_add_223_n157,
         DP_add_1_root_add_0_root_add_223_n156,
         DP_add_1_root_add_0_root_add_223_n155,
         DP_add_1_root_add_0_root_add_223_n154,
         DP_add_1_root_add_0_root_add_223_n153,
         DP_add_1_root_add_0_root_add_223_n152,
         DP_add_1_root_add_0_root_add_223_n151,
         DP_add_1_root_add_0_root_add_223_n150,
         DP_add_1_root_add_0_root_add_223_n149,
         DP_add_1_root_add_0_root_add_223_n148,
         DP_add_1_root_add_0_root_add_223_n147,
         DP_add_1_root_add_0_root_add_223_n145,
         DP_add_1_root_add_0_root_add_223_n143,
         DP_add_1_root_add_0_root_add_223_n142,
         DP_add_1_root_add_0_root_add_223_n141,
         DP_add_1_root_add_0_root_add_223_n140,
         DP_add_1_root_add_0_root_add_223_n139,
         DP_add_1_root_add_0_root_add_223_n138,
         DP_add_1_root_add_0_root_add_223_n137,
         DP_add_1_root_add_0_root_add_223_n136,
         DP_add_1_root_add_0_root_add_223_n135,
         DP_add_1_root_add_0_root_add_223_n134,
         DP_add_1_root_add_0_root_add_223_n133,
         DP_add_1_root_add_0_root_add_223_n132,
         DP_add_1_root_add_0_root_add_223_n131,
         DP_add_1_root_add_0_root_add_223_n130,
         DP_add_1_root_add_0_root_add_223_n129,
         DP_add_1_root_add_0_root_add_223_n128,
         DP_add_1_root_add_0_root_add_223_n127,
         DP_add_1_root_add_0_root_add_223_n126,
         DP_add_1_root_add_0_root_add_223_n125,
         DP_add_1_root_add_0_root_add_223_n124,
         DP_add_1_root_add_0_root_add_223_n123,
         DP_add_1_root_add_0_root_add_223_n122,
         DP_add_1_root_add_0_root_add_223_n121,
         DP_add_1_root_add_0_root_add_223_n120,
         DP_add_1_root_add_0_root_add_223_n119,
         DP_add_1_root_add_0_root_add_223_n118,
         DP_add_1_root_add_0_root_add_223_n117,
         DP_add_1_root_add_0_root_add_223_n116,
         DP_add_1_root_add_0_root_add_223_n115,
         DP_add_1_root_add_0_root_add_223_n114,
         DP_add_1_root_add_0_root_add_223_n113,
         DP_add_1_root_add_0_root_add_223_n112,
         DP_add_1_root_add_0_root_add_223_n111,
         DP_add_1_root_add_0_root_add_223_n110,
         DP_add_1_root_add_0_root_add_223_n109,
         DP_add_1_root_add_0_root_add_223_n108,
         DP_add_1_root_add_0_root_add_223_n107,
         DP_add_1_root_add_0_root_add_223_n106,
         DP_add_1_root_add_0_root_add_223_n105,
         DP_add_1_root_add_0_root_add_223_n104,
         DP_add_1_root_add_0_root_add_223_n103,
         DP_add_1_root_add_0_root_add_223_n102,
         DP_add_1_root_add_0_root_add_223_n101,
         DP_add_1_root_add_0_root_add_223_n100,
         DP_add_1_root_add_0_root_add_223_n99,
         DP_add_1_root_add_0_root_add_223_n98,
         DP_add_1_root_add_0_root_add_223_n97,
         DP_add_1_root_add_0_root_add_223_n96,
         DP_add_1_root_add_0_root_add_223_n95,
         DP_add_1_root_add_0_root_add_223_n94,
         DP_add_1_root_add_0_root_add_223_n93,
         DP_add_1_root_add_0_root_add_223_n92,
         DP_add_1_root_add_0_root_add_223_n91,
         DP_add_1_root_add_0_root_add_223_n90,
         DP_add_1_root_add_0_root_add_223_n89,
         DP_add_1_root_add_0_root_add_223_n88,
         DP_add_1_root_add_0_root_add_223_n87,
         DP_add_1_root_add_0_root_add_223_n86,
         DP_add_1_root_add_0_root_add_223_n85,
         DP_add_1_root_add_0_root_add_223_n84,
         DP_add_1_root_add_0_root_add_223_n83,
         DP_add_1_root_add_0_root_add_223_n82,
         DP_add_1_root_add_0_root_add_223_n81,
         DP_add_1_root_add_0_root_add_223_n80,
         DP_add_1_root_add_0_root_add_223_n79,
         DP_add_1_root_add_0_root_add_223_n77,
         DP_add_1_root_add_0_root_add_223_n75,
         DP_add_1_root_add_0_root_add_223_n74,
         DP_add_1_root_add_0_root_add_223_n73,
         DP_add_1_root_add_0_root_add_223_n72,
         DP_add_1_root_add_0_root_add_223_n71,
         DP_add_1_root_add_0_root_add_223_n70,
         DP_add_1_root_add_0_root_add_223_n69,
         DP_add_1_root_add_0_root_add_223_n68,
         DP_add_1_root_add_0_root_add_223_n67,
         DP_add_1_root_add_0_root_add_223_n66,
         DP_add_1_root_add_0_root_add_223_n65,
         DP_add_1_root_add_0_root_add_223_n64,
         DP_add_1_root_add_0_root_add_223_n63,
         DP_add_1_root_add_0_root_add_223_n62,
         DP_add_1_root_add_0_root_add_223_n61,
         DP_add_1_root_add_0_root_add_223_n60,
         DP_add_1_root_add_0_root_add_223_n59,
         DP_add_1_root_add_0_root_add_223_n58,
         DP_add_1_root_add_0_root_add_223_n57,
         DP_add_1_root_add_0_root_add_223_n56,
         DP_add_1_root_add_0_root_add_223_n55,
         DP_add_1_root_add_0_root_add_223_n54,
         DP_add_1_root_add_0_root_add_223_n53,
         DP_add_1_root_add_0_root_add_223_n52,
         DP_add_1_root_add_0_root_add_223_n51,
         DP_add_1_root_add_0_root_add_223_n50,
         DP_add_1_root_add_0_root_add_223_n49,
         DP_add_1_root_add_0_root_add_223_n48,
         DP_add_1_root_add_0_root_add_223_n47,
         DP_add_1_root_add_0_root_add_223_n46,
         DP_add_1_root_add_0_root_add_223_n45,
         DP_add_1_root_add_0_root_add_223_n44,
         DP_add_1_root_add_0_root_add_223_n43,
         DP_add_1_root_add_0_root_add_223_n42,
         DP_add_1_root_add_0_root_add_223_n41,
         DP_add_1_root_add_0_root_add_223_n40,
         DP_add_1_root_add_0_root_add_223_n39,
         DP_add_1_root_add_0_root_add_223_n38,
         DP_add_1_root_add_0_root_add_223_n37,
         DP_add_1_root_add_0_root_add_223_n36,
         DP_add_1_root_add_0_root_add_223_n35,
         DP_add_1_root_add_0_root_add_223_n34,
         DP_add_1_root_add_0_root_add_223_n33,
         DP_add_1_root_add_0_root_add_223_n32,
         DP_add_1_root_add_0_root_add_223_n30,
         DP_add_1_root_add_0_root_add_223_n28,
         DP_add_1_root_add_0_root_add_223_n27,
         DP_add_1_root_add_0_root_add_223_n24,
         DP_add_1_root_add_0_root_add_223_n23,
         DP_add_1_root_add_0_root_add_223_n22,
         DP_add_1_root_add_0_root_add_223_n21,
         DP_add_1_root_add_0_root_add_223_n20,
         DP_add_1_root_add_0_root_add_223_n19,
         DP_add_1_root_add_0_root_add_223_n18,
         DP_add_1_root_add_0_root_add_223_n17,
         DP_add_1_root_add_0_root_add_223_n16,
         DP_add_1_root_add_0_root_add_223_n15,
         DP_add_1_root_add_0_root_add_223_n14,
         DP_add_1_root_add_0_root_add_223_n13,
         DP_add_1_root_add_0_root_add_223_n12,
         DP_add_1_root_add_0_root_add_223_n11,
         DP_add_1_root_add_0_root_add_223_n10,
         DP_add_1_root_add_0_root_add_223_n9,
         DP_add_1_root_add_0_root_add_223_n8,
         DP_add_1_root_add_0_root_add_223_n7,
         DP_add_1_root_add_0_root_add_223_n6,
         DP_add_1_root_add_0_root_add_223_n5,
         DP_add_1_root_add_0_root_add_223_n4,
         DP_add_1_root_add_0_root_add_223_n3,
         DP_add_1_root_add_0_root_add_223_n2,
         DP_add_1_root_add_0_root_add_223_n1,
         DP_add_1_root_sub_0_root_sub_217_n297,
         DP_add_1_root_sub_0_root_sub_217_n296,
         DP_add_1_root_sub_0_root_sub_217_n295,
         DP_add_1_root_sub_0_root_sub_217_n293,
         DP_add_1_root_sub_0_root_sub_217_n213,
         DP_add_1_root_sub_0_root_sub_217_n212,
         DP_add_1_root_sub_0_root_sub_217_n211,
         DP_add_1_root_sub_0_root_sub_217_n209,
         DP_add_1_root_sub_0_root_sub_217_n208,
         DP_add_1_root_sub_0_root_sub_217_n207,
         DP_add_1_root_sub_0_root_sub_217_n206,
         DP_add_1_root_sub_0_root_sub_217_n205,
         DP_add_1_root_sub_0_root_sub_217_n203,
         DP_add_1_root_sub_0_root_sub_217_n201,
         DP_add_1_root_sub_0_root_sub_217_n199,
         DP_add_1_root_sub_0_root_sub_217_n198,
         DP_add_1_root_sub_0_root_sub_217_n197,
         DP_add_1_root_sub_0_root_sub_217_n195,
         DP_add_1_root_sub_0_root_sub_217_n193,
         DP_add_1_root_sub_0_root_sub_217_n190,
         DP_add_1_root_sub_0_root_sub_217_n188,
         DP_add_1_root_sub_0_root_sub_217_n187,
         DP_add_1_root_sub_0_root_sub_217_n186,
         DP_add_1_root_sub_0_root_sub_217_n185,
         DP_add_1_root_sub_0_root_sub_217_n184,
         DP_add_1_root_sub_0_root_sub_217_n183,
         DP_add_1_root_sub_0_root_sub_217_n182,
         DP_add_1_root_sub_0_root_sub_217_n181,
         DP_add_1_root_sub_0_root_sub_217_n180,
         DP_add_1_root_sub_0_root_sub_217_n179,
         DP_add_1_root_sub_0_root_sub_217_n178,
         DP_add_1_root_sub_0_root_sub_217_n177,
         DP_add_1_root_sub_0_root_sub_217_n176,
         DP_add_1_root_sub_0_root_sub_217_n175,
         DP_add_1_root_sub_0_root_sub_217_n174,
         DP_add_1_root_sub_0_root_sub_217_n173,
         DP_add_1_root_sub_0_root_sub_217_n172,
         DP_add_1_root_sub_0_root_sub_217_n171,
         DP_add_1_root_sub_0_root_sub_217_n170,
         DP_add_1_root_sub_0_root_sub_217_n169,
         DP_add_1_root_sub_0_root_sub_217_n168,
         DP_add_1_root_sub_0_root_sub_217_n167,
         DP_add_1_root_sub_0_root_sub_217_n166,
         DP_add_1_root_sub_0_root_sub_217_n165,
         DP_add_1_root_sub_0_root_sub_217_n164,
         DP_add_1_root_sub_0_root_sub_217_n163,
         DP_add_1_root_sub_0_root_sub_217_n162,
         DP_add_1_root_sub_0_root_sub_217_n161,
         DP_add_1_root_sub_0_root_sub_217_n160,
         DP_add_1_root_sub_0_root_sub_217_n159,
         DP_add_1_root_sub_0_root_sub_217_n158,
         DP_add_1_root_sub_0_root_sub_217_n157,
         DP_add_1_root_sub_0_root_sub_217_n156,
         DP_add_1_root_sub_0_root_sub_217_n155,
         DP_add_1_root_sub_0_root_sub_217_n154,
         DP_add_1_root_sub_0_root_sub_217_n153,
         DP_add_1_root_sub_0_root_sub_217_n152,
         DP_add_1_root_sub_0_root_sub_217_n151,
         DP_add_1_root_sub_0_root_sub_217_n150,
         DP_add_1_root_sub_0_root_sub_217_n149,
         DP_add_1_root_sub_0_root_sub_217_n148,
         DP_add_1_root_sub_0_root_sub_217_n147,
         DP_add_1_root_sub_0_root_sub_217_n145,
         DP_add_1_root_sub_0_root_sub_217_n143,
         DP_add_1_root_sub_0_root_sub_217_n142,
         DP_add_1_root_sub_0_root_sub_217_n141,
         DP_add_1_root_sub_0_root_sub_217_n140,
         DP_add_1_root_sub_0_root_sub_217_n139,
         DP_add_1_root_sub_0_root_sub_217_n138,
         DP_add_1_root_sub_0_root_sub_217_n137,
         DP_add_1_root_sub_0_root_sub_217_n136,
         DP_add_1_root_sub_0_root_sub_217_n135,
         DP_add_1_root_sub_0_root_sub_217_n134,
         DP_add_1_root_sub_0_root_sub_217_n133,
         DP_add_1_root_sub_0_root_sub_217_n132,
         DP_add_1_root_sub_0_root_sub_217_n131,
         DP_add_1_root_sub_0_root_sub_217_n130,
         DP_add_1_root_sub_0_root_sub_217_n129,
         DP_add_1_root_sub_0_root_sub_217_n128,
         DP_add_1_root_sub_0_root_sub_217_n127,
         DP_add_1_root_sub_0_root_sub_217_n126,
         DP_add_1_root_sub_0_root_sub_217_n125,
         DP_add_1_root_sub_0_root_sub_217_n124,
         DP_add_1_root_sub_0_root_sub_217_n123,
         DP_add_1_root_sub_0_root_sub_217_n122,
         DP_add_1_root_sub_0_root_sub_217_n121,
         DP_add_1_root_sub_0_root_sub_217_n120,
         DP_add_1_root_sub_0_root_sub_217_n119,
         DP_add_1_root_sub_0_root_sub_217_n118,
         DP_add_1_root_sub_0_root_sub_217_n117,
         DP_add_1_root_sub_0_root_sub_217_n116,
         DP_add_1_root_sub_0_root_sub_217_n115,
         DP_add_1_root_sub_0_root_sub_217_n114,
         DP_add_1_root_sub_0_root_sub_217_n113,
         DP_add_1_root_sub_0_root_sub_217_n112,
         DP_add_1_root_sub_0_root_sub_217_n111,
         DP_add_1_root_sub_0_root_sub_217_n110,
         DP_add_1_root_sub_0_root_sub_217_n109,
         DP_add_1_root_sub_0_root_sub_217_n108,
         DP_add_1_root_sub_0_root_sub_217_n107,
         DP_add_1_root_sub_0_root_sub_217_n106,
         DP_add_1_root_sub_0_root_sub_217_n105,
         DP_add_1_root_sub_0_root_sub_217_n104,
         DP_add_1_root_sub_0_root_sub_217_n103,
         DP_add_1_root_sub_0_root_sub_217_n102,
         DP_add_1_root_sub_0_root_sub_217_n101,
         DP_add_1_root_sub_0_root_sub_217_n100,
         DP_add_1_root_sub_0_root_sub_217_n99,
         DP_add_1_root_sub_0_root_sub_217_n98,
         DP_add_1_root_sub_0_root_sub_217_n97,
         DP_add_1_root_sub_0_root_sub_217_n96,
         DP_add_1_root_sub_0_root_sub_217_n95,
         DP_add_1_root_sub_0_root_sub_217_n94,
         DP_add_1_root_sub_0_root_sub_217_n93,
         DP_add_1_root_sub_0_root_sub_217_n92,
         DP_add_1_root_sub_0_root_sub_217_n91,
         DP_add_1_root_sub_0_root_sub_217_n90,
         DP_add_1_root_sub_0_root_sub_217_n89,
         DP_add_1_root_sub_0_root_sub_217_n88,
         DP_add_1_root_sub_0_root_sub_217_n87,
         DP_add_1_root_sub_0_root_sub_217_n86,
         DP_add_1_root_sub_0_root_sub_217_n85,
         DP_add_1_root_sub_0_root_sub_217_n84,
         DP_add_1_root_sub_0_root_sub_217_n83,
         DP_add_1_root_sub_0_root_sub_217_n82,
         DP_add_1_root_sub_0_root_sub_217_n81,
         DP_add_1_root_sub_0_root_sub_217_n80,
         DP_add_1_root_sub_0_root_sub_217_n79,
         DP_add_1_root_sub_0_root_sub_217_n78,
         DP_add_1_root_sub_0_root_sub_217_n77,
         DP_add_1_root_sub_0_root_sub_217_n76,
         DP_add_1_root_sub_0_root_sub_217_n75,
         DP_add_1_root_sub_0_root_sub_217_n74,
         DP_add_1_root_sub_0_root_sub_217_n73,
         DP_add_1_root_sub_0_root_sub_217_n72,
         DP_add_1_root_sub_0_root_sub_217_n71,
         DP_add_1_root_sub_0_root_sub_217_n70,
         DP_add_1_root_sub_0_root_sub_217_n69,
         DP_add_1_root_sub_0_root_sub_217_n68,
         DP_add_1_root_sub_0_root_sub_217_n67,
         DP_add_1_root_sub_0_root_sub_217_n66,
         DP_add_1_root_sub_0_root_sub_217_n65,
         DP_add_1_root_sub_0_root_sub_217_n64,
         DP_add_1_root_sub_0_root_sub_217_n63,
         DP_add_1_root_sub_0_root_sub_217_n62,
         DP_add_1_root_sub_0_root_sub_217_n61,
         DP_add_1_root_sub_0_root_sub_217_n60,
         DP_add_1_root_sub_0_root_sub_217_n59,
         DP_add_1_root_sub_0_root_sub_217_n58,
         DP_add_1_root_sub_0_root_sub_217_n57,
         DP_add_1_root_sub_0_root_sub_217_n56,
         DP_add_1_root_sub_0_root_sub_217_n55,
         DP_add_1_root_sub_0_root_sub_217_n54,
         DP_add_1_root_sub_0_root_sub_217_n53,
         DP_add_1_root_sub_0_root_sub_217_n52,
         DP_add_1_root_sub_0_root_sub_217_n51,
         DP_add_1_root_sub_0_root_sub_217_n50,
         DP_add_1_root_sub_0_root_sub_217_n49,
         DP_add_1_root_sub_0_root_sub_217_n48,
         DP_add_1_root_sub_0_root_sub_217_n47,
         DP_add_1_root_sub_0_root_sub_217_n46,
         DP_add_1_root_sub_0_root_sub_217_n45,
         DP_add_1_root_sub_0_root_sub_217_n44,
         DP_add_1_root_sub_0_root_sub_217_n43,
         DP_add_1_root_sub_0_root_sub_217_n42,
         DP_add_1_root_sub_0_root_sub_217_n41,
         DP_add_1_root_sub_0_root_sub_217_n40,
         DP_add_1_root_sub_0_root_sub_217_n39,
         DP_add_1_root_sub_0_root_sub_217_n38,
         DP_add_1_root_sub_0_root_sub_217_n36,
         DP_add_1_root_sub_0_root_sub_217_n34,
         DP_add_1_root_sub_0_root_sub_217_n33,
         DP_add_1_root_sub_0_root_sub_217_n32,
         DP_add_1_root_sub_0_root_sub_217_n30,
         DP_add_1_root_sub_0_root_sub_217_n28,
         DP_add_1_root_sub_0_root_sub_217_n27,
         DP_add_1_root_sub_0_root_sub_217_n24,
         DP_add_1_root_sub_0_root_sub_217_n23,
         DP_add_1_root_sub_0_root_sub_217_n22,
         DP_add_1_root_sub_0_root_sub_217_n21,
         DP_add_1_root_sub_0_root_sub_217_n20,
         DP_add_1_root_sub_0_root_sub_217_n19,
         DP_add_1_root_sub_0_root_sub_217_n18,
         DP_add_1_root_sub_0_root_sub_217_n17,
         DP_add_1_root_sub_0_root_sub_217_n16,
         DP_add_1_root_sub_0_root_sub_217_n15,
         DP_add_1_root_sub_0_root_sub_217_n14,
         DP_add_1_root_sub_0_root_sub_217_n13,
         DP_add_1_root_sub_0_root_sub_217_n12,
         DP_add_1_root_sub_0_root_sub_217_n11,
         DP_add_1_root_sub_0_root_sub_217_n10,
         DP_add_1_root_sub_0_root_sub_217_n9,
         DP_add_1_root_sub_0_root_sub_217_n8,
         DP_add_1_root_sub_0_root_sub_217_n7,
         DP_add_1_root_sub_0_root_sub_217_n6,
         DP_add_1_root_sub_0_root_sub_217_n5,
         DP_add_1_root_sub_0_root_sub_217_n4,
         DP_add_1_root_sub_0_root_sub_217_n3,
         DP_add_1_root_sub_0_root_sub_217_n2,
         DP_add_1_root_sub_0_root_sub_217_n1,
         DP_sub_0_root_sub_0_root_sub_217_n239,
         DP_sub_0_root_sub_0_root_sub_217_n238,
         DP_sub_0_root_sub_0_root_sub_217_n161,
         DP_sub_0_root_sub_0_root_sub_217_n160,
         DP_sub_0_root_sub_0_root_sub_217_n159,
         DP_sub_0_root_sub_0_root_sub_217_n158,
         DP_sub_0_root_sub_0_root_sub_217_n157,
         DP_sub_0_root_sub_0_root_sub_217_n156,
         DP_sub_0_root_sub_0_root_sub_217_n155,
         DP_sub_0_root_sub_0_root_sub_217_n154,
         DP_sub_0_root_sub_0_root_sub_217_n153,
         DP_sub_0_root_sub_0_root_sub_217_n152,
         DP_sub_0_root_sub_0_root_sub_217_n151,
         DP_sub_0_root_sub_0_root_sub_217_n150,
         DP_sub_0_root_sub_0_root_sub_217_n149,
         DP_sub_0_root_sub_0_root_sub_217_n148,
         DP_sub_0_root_sub_0_root_sub_217_n147,
         DP_sub_0_root_sub_0_root_sub_217_n146,
         DP_sub_0_root_sub_0_root_sub_217_n145,
         DP_sub_0_root_sub_0_root_sub_217_n143,
         DP_sub_0_root_sub_0_root_sub_217_n141,
         DP_sub_0_root_sub_0_root_sub_217_n139,
         DP_sub_0_root_sub_0_root_sub_217_n138,
         DP_sub_0_root_sub_0_root_sub_217_n137,
         DP_sub_0_root_sub_0_root_sub_217_n135,
         DP_sub_0_root_sub_0_root_sub_217_n134,
         DP_sub_0_root_sub_0_root_sub_217_n133,
         DP_sub_0_root_sub_0_root_sub_217_n132,
         DP_sub_0_root_sub_0_root_sub_217_n131,
         DP_sub_0_root_sub_0_root_sub_217_n130,
         DP_sub_0_root_sub_0_root_sub_217_n129,
         DP_sub_0_root_sub_0_root_sub_217_n128,
         DP_sub_0_root_sub_0_root_sub_217_n127,
         DP_sub_0_root_sub_0_root_sub_217_n126,
         DP_sub_0_root_sub_0_root_sub_217_n125,
         DP_sub_0_root_sub_0_root_sub_217_n124,
         DP_sub_0_root_sub_0_root_sub_217_n123,
         DP_sub_0_root_sub_0_root_sub_217_n122,
         DP_sub_0_root_sub_0_root_sub_217_n121,
         DP_sub_0_root_sub_0_root_sub_217_n120,
         DP_sub_0_root_sub_0_root_sub_217_n119,
         DP_sub_0_root_sub_0_root_sub_217_n118,
         DP_sub_0_root_sub_0_root_sub_217_n117,
         DP_sub_0_root_sub_0_root_sub_217_n116,
         DP_sub_0_root_sub_0_root_sub_217_n115,
         DP_sub_0_root_sub_0_root_sub_217_n114,
         DP_sub_0_root_sub_0_root_sub_217_n113,
         DP_sub_0_root_sub_0_root_sub_217_n112,
         DP_sub_0_root_sub_0_root_sub_217_n111,
         DP_sub_0_root_sub_0_root_sub_217_n110,
         DP_sub_0_root_sub_0_root_sub_217_n109,
         DP_sub_0_root_sub_0_root_sub_217_n108,
         DP_sub_0_root_sub_0_root_sub_217_n107,
         DP_sub_0_root_sub_0_root_sub_217_n106,
         DP_sub_0_root_sub_0_root_sub_217_n105,
         DP_sub_0_root_sub_0_root_sub_217_n104,
         DP_sub_0_root_sub_0_root_sub_217_n103,
         DP_sub_0_root_sub_0_root_sub_217_n102,
         DP_sub_0_root_sub_0_root_sub_217_n101,
         DP_sub_0_root_sub_0_root_sub_217_n100,
         DP_sub_0_root_sub_0_root_sub_217_n99,
         DP_sub_0_root_sub_0_root_sub_217_n98,
         DP_sub_0_root_sub_0_root_sub_217_n97,
         DP_sub_0_root_sub_0_root_sub_217_n96,
         DP_sub_0_root_sub_0_root_sub_217_n95,
         DP_sub_0_root_sub_0_root_sub_217_n94,
         DP_sub_0_root_sub_0_root_sub_217_n93,
         DP_sub_0_root_sub_0_root_sub_217_n92,
         DP_sub_0_root_sub_0_root_sub_217_n91,
         DP_sub_0_root_sub_0_root_sub_217_n90,
         DP_sub_0_root_sub_0_root_sub_217_n89,
         DP_sub_0_root_sub_0_root_sub_217_n88,
         DP_sub_0_root_sub_0_root_sub_217_n87,
         DP_sub_0_root_sub_0_root_sub_217_n86,
         DP_sub_0_root_sub_0_root_sub_217_n84,
         DP_sub_0_root_sub_0_root_sub_217_n82,
         DP_sub_0_root_sub_0_root_sub_217_n81,
         DP_sub_0_root_sub_0_root_sub_217_n80,
         DP_sub_0_root_sub_0_root_sub_217_n79,
         DP_sub_0_root_sub_0_root_sub_217_n78,
         DP_sub_0_root_sub_0_root_sub_217_n77,
         DP_sub_0_root_sub_0_root_sub_217_n76,
         DP_sub_0_root_sub_0_root_sub_217_n75,
         DP_sub_0_root_sub_0_root_sub_217_n74,
         DP_sub_0_root_sub_0_root_sub_217_n73,
         DP_sub_0_root_sub_0_root_sub_217_n72,
         DP_sub_0_root_sub_0_root_sub_217_n71,
         DP_sub_0_root_sub_0_root_sub_217_n70,
         DP_sub_0_root_sub_0_root_sub_217_n69,
         DP_sub_0_root_sub_0_root_sub_217_n68,
         DP_sub_0_root_sub_0_root_sub_217_n67,
         DP_sub_0_root_sub_0_root_sub_217_n66,
         DP_sub_0_root_sub_0_root_sub_217_n65,
         DP_sub_0_root_sub_0_root_sub_217_n64,
         DP_sub_0_root_sub_0_root_sub_217_n63,
         DP_sub_0_root_sub_0_root_sub_217_n62,
         DP_sub_0_root_sub_0_root_sub_217_n61,
         DP_sub_0_root_sub_0_root_sub_217_n60,
         DP_sub_0_root_sub_0_root_sub_217_n59,
         DP_sub_0_root_sub_0_root_sub_217_n58,
         DP_sub_0_root_sub_0_root_sub_217_n57,
         DP_sub_0_root_sub_0_root_sub_217_n56,
         DP_sub_0_root_sub_0_root_sub_217_n55,
         DP_sub_0_root_sub_0_root_sub_217_n54,
         DP_sub_0_root_sub_0_root_sub_217_n53,
         DP_sub_0_root_sub_0_root_sub_217_n52,
         DP_sub_0_root_sub_0_root_sub_217_n51,
         DP_sub_0_root_sub_0_root_sub_217_n50,
         DP_sub_0_root_sub_0_root_sub_217_n49,
         DP_sub_0_root_sub_0_root_sub_217_n48,
         DP_sub_0_root_sub_0_root_sub_217_n47,
         DP_sub_0_root_sub_0_root_sub_217_n46,
         DP_sub_0_root_sub_0_root_sub_217_n45,
         DP_sub_0_root_sub_0_root_sub_217_n44,
         DP_sub_0_root_sub_0_root_sub_217_n43,
         DP_sub_0_root_sub_0_root_sub_217_n42,
         DP_sub_0_root_sub_0_root_sub_217_n41,
         DP_sub_0_root_sub_0_root_sub_217_n40,
         DP_sub_0_root_sub_0_root_sub_217_n39,
         DP_sub_0_root_sub_0_root_sub_217_n38,
         DP_sub_0_root_sub_0_root_sub_217_n37,
         DP_sub_0_root_sub_0_root_sub_217_n36,
         DP_sub_0_root_sub_0_root_sub_217_n35,
         DP_sub_0_root_sub_0_root_sub_217_n34,
         DP_sub_0_root_sub_0_root_sub_217_n33,
         DP_sub_0_root_sub_0_root_sub_217_n32,
         DP_sub_0_root_sub_0_root_sub_217_n31,
         DP_sub_0_root_sub_0_root_sub_217_n30,
         DP_sub_0_root_sub_0_root_sub_217_n29,
         DP_sub_0_root_sub_0_root_sub_217_n28,
         DP_sub_0_root_sub_0_root_sub_217_n27,
         DP_sub_0_root_sub_0_root_sub_217_n26,
         DP_sub_0_root_sub_0_root_sub_217_n25,
         DP_sub_0_root_sub_0_root_sub_217_n24,
         DP_sub_0_root_sub_0_root_sub_217_n23,
         DP_sub_0_root_sub_0_root_sub_217_n22,
         DP_sub_0_root_sub_0_root_sub_217_n21,
         DP_sub_0_root_sub_0_root_sub_217_n19,
         DP_sub_0_root_sub_0_root_sub_217_n17,
         DP_sub_0_root_sub_0_root_sub_217_n16,
         DP_sub_0_root_sub_0_root_sub_217_n14,
         DP_sub_0_root_sub_0_root_sub_217_n13,
         DP_sub_0_root_sub_0_root_sub_217_n12,
         DP_sub_0_root_sub_0_root_sub_217_n11,
         DP_sub_0_root_sub_0_root_sub_217_n10,
         DP_sub_0_root_sub_0_root_sub_217_n9,
         DP_sub_0_root_sub_0_root_sub_217_n8,
         DP_sub_0_root_sub_0_root_sub_217_n7,
         DP_sub_0_root_sub_0_root_sub_217_n6,
         DP_sub_0_root_sub_0_root_sub_217_n5,
         DP_sub_0_root_sub_0_root_sub_217_n4,
         DP_sub_0_root_sub_0_root_sub_217_n3,
         DP_sub_0_root_sub_0_root_sub_217_n2,
         DP_sub_0_root_sub_0_root_sub_217_n1,
         DP_add_0_root_add_0_root_add_223_n245,
         DP_add_0_root_add_0_root_add_223_n244,
         DP_add_0_root_add_0_root_add_223_n243,
         DP_add_0_root_add_0_root_add_223_n175,
         DP_add_0_root_add_0_root_add_223_n173,
         DP_add_0_root_add_0_root_add_223_n171,
         DP_add_0_root_add_0_root_add_223_n170,
         DP_add_0_root_add_0_root_add_223_n169,
         DP_add_0_root_add_0_root_add_223_n167,
         DP_add_0_root_add_0_root_add_223_n166,
         DP_add_0_root_add_0_root_add_223_n165,
         DP_add_0_root_add_0_root_add_223_n162,
         DP_add_0_root_add_0_root_add_223_n161,
         DP_add_0_root_add_0_root_add_223_n160,
         DP_add_0_root_add_0_root_add_223_n159,
         DP_add_0_root_add_0_root_add_223_n158,
         DP_add_0_root_add_0_root_add_223_n157,
         DP_add_0_root_add_0_root_add_223_n156,
         DP_add_0_root_add_0_root_add_223_n155,
         DP_add_0_root_add_0_root_add_223_n154,
         DP_add_0_root_add_0_root_add_223_n153,
         DP_add_0_root_add_0_root_add_223_n152,
         DP_add_0_root_add_0_root_add_223_n151,
         DP_add_0_root_add_0_root_add_223_n150,
         DP_add_0_root_add_0_root_add_223_n149,
         DP_add_0_root_add_0_root_add_223_n148,
         DP_add_0_root_add_0_root_add_223_n147,
         DP_add_0_root_add_0_root_add_223_n146,
         DP_add_0_root_add_0_root_add_223_n145,
         DP_add_0_root_add_0_root_add_223_n144,
         DP_add_0_root_add_0_root_add_223_n143,
         DP_add_0_root_add_0_root_add_223_n142,
         DP_add_0_root_add_0_root_add_223_n141,
         DP_add_0_root_add_0_root_add_223_n140,
         DP_add_0_root_add_0_root_add_223_n139,
         DP_add_0_root_add_0_root_add_223_n138,
         DP_add_0_root_add_0_root_add_223_n137,
         DP_add_0_root_add_0_root_add_223_n136,
         DP_add_0_root_add_0_root_add_223_n135,
         DP_add_0_root_add_0_root_add_223_n134,
         DP_add_0_root_add_0_root_add_223_n133,
         DP_add_0_root_add_0_root_add_223_n132,
         DP_add_0_root_add_0_root_add_223_n131,
         DP_add_0_root_add_0_root_add_223_n130,
         DP_add_0_root_add_0_root_add_223_n129,
         DP_add_0_root_add_0_root_add_223_n128,
         DP_add_0_root_add_0_root_add_223_n127,
         DP_add_0_root_add_0_root_add_223_n126,
         DP_add_0_root_add_0_root_add_223_n125,
         DP_add_0_root_add_0_root_add_223_n124,
         DP_add_0_root_add_0_root_add_223_n123,
         DP_add_0_root_add_0_root_add_223_n122,
         DP_add_0_root_add_0_root_add_223_n121,
         DP_add_0_root_add_0_root_add_223_n120,
         DP_add_0_root_add_0_root_add_223_n119,
         DP_add_0_root_add_0_root_add_223_n118,
         DP_add_0_root_add_0_root_add_223_n117,
         DP_add_0_root_add_0_root_add_223_n116,
         DP_add_0_root_add_0_root_add_223_n115,
         DP_add_0_root_add_0_root_add_223_n114,
         DP_add_0_root_add_0_root_add_223_n113,
         DP_add_0_root_add_0_root_add_223_n112,
         DP_add_0_root_add_0_root_add_223_n111,
         DP_add_0_root_add_0_root_add_223_n110,
         DP_add_0_root_add_0_root_add_223_n109,
         DP_add_0_root_add_0_root_add_223_n108,
         DP_add_0_root_add_0_root_add_223_n107,
         DP_add_0_root_add_0_root_add_223_n106,
         DP_add_0_root_add_0_root_add_223_n105,
         DP_add_0_root_add_0_root_add_223_n104,
         DP_add_0_root_add_0_root_add_223_n103,
         DP_add_0_root_add_0_root_add_223_n102,
         DP_add_0_root_add_0_root_add_223_n101,
         DP_add_0_root_add_0_root_add_223_n100,
         DP_add_0_root_add_0_root_add_223_n99,
         DP_add_0_root_add_0_root_add_223_n98,
         DP_add_0_root_add_0_root_add_223_n97,
         DP_add_0_root_add_0_root_add_223_n96,
         DP_add_0_root_add_0_root_add_223_n95,
         DP_add_0_root_add_0_root_add_223_n94,
         DP_add_0_root_add_0_root_add_223_n93,
         DP_add_0_root_add_0_root_add_223_n92,
         DP_add_0_root_add_0_root_add_223_n91,
         DP_add_0_root_add_0_root_add_223_n90,
         DP_add_0_root_add_0_root_add_223_n89,
         DP_add_0_root_add_0_root_add_223_n88,
         DP_add_0_root_add_0_root_add_223_n87,
         DP_add_0_root_add_0_root_add_223_n86,
         DP_add_0_root_add_0_root_add_223_n85,
         DP_add_0_root_add_0_root_add_223_n84,
         DP_add_0_root_add_0_root_add_223_n83,
         DP_add_0_root_add_0_root_add_223_n82,
         DP_add_0_root_add_0_root_add_223_n81,
         DP_add_0_root_add_0_root_add_223_n80,
         DP_add_0_root_add_0_root_add_223_n79,
         DP_add_0_root_add_0_root_add_223_n78,
         DP_add_0_root_add_0_root_add_223_n77,
         DP_add_0_root_add_0_root_add_223_n76,
         DP_add_0_root_add_0_root_add_223_n75,
         DP_add_0_root_add_0_root_add_223_n74,
         DP_add_0_root_add_0_root_add_223_n73,
         DP_add_0_root_add_0_root_add_223_n72,
         DP_add_0_root_add_0_root_add_223_n71,
         DP_add_0_root_add_0_root_add_223_n70,
         DP_add_0_root_add_0_root_add_223_n69,
         DP_add_0_root_add_0_root_add_223_n68,
         DP_add_0_root_add_0_root_add_223_n66,
         DP_add_0_root_add_0_root_add_223_n64,
         DP_add_0_root_add_0_root_add_223_n63,
         DP_add_0_root_add_0_root_add_223_n62,
         DP_add_0_root_add_0_root_add_223_n61,
         DP_add_0_root_add_0_root_add_223_n60,
         DP_add_0_root_add_0_root_add_223_n59,
         DP_add_0_root_add_0_root_add_223_n58,
         DP_add_0_root_add_0_root_add_223_n57,
         DP_add_0_root_add_0_root_add_223_n56,
         DP_add_0_root_add_0_root_add_223_n55,
         DP_add_0_root_add_0_root_add_223_n54,
         DP_add_0_root_add_0_root_add_223_n53,
         DP_add_0_root_add_0_root_add_223_n52,
         DP_add_0_root_add_0_root_add_223_n51,
         DP_add_0_root_add_0_root_add_223_n50,
         DP_add_0_root_add_0_root_add_223_n49,
         DP_add_0_root_add_0_root_add_223_n48,
         DP_add_0_root_add_0_root_add_223_n47,
         DP_add_0_root_add_0_root_add_223_n46,
         DP_add_0_root_add_0_root_add_223_n45,
         DP_add_0_root_add_0_root_add_223_n44,
         DP_add_0_root_add_0_root_add_223_n43,
         DP_add_0_root_add_0_root_add_223_n42,
         DP_add_0_root_add_0_root_add_223_n41,
         DP_add_0_root_add_0_root_add_223_n39,
         DP_add_0_root_add_0_root_add_223_n38,
         DP_add_0_root_add_0_root_add_223_n37,
         DP_add_0_root_add_0_root_add_223_n36,
         DP_add_0_root_add_0_root_add_223_n35,
         DP_add_0_root_add_0_root_add_223_n34,
         DP_add_0_root_add_0_root_add_223_n33,
         DP_add_0_root_add_0_root_add_223_n32,
         DP_add_0_root_add_0_root_add_223_n31,
         DP_add_0_root_add_0_root_add_223_n30,
         DP_add_0_root_add_0_root_add_223_n29,
         DP_add_0_root_add_0_root_add_223_n28,
         DP_add_0_root_add_0_root_add_223_n27,
         DP_add_0_root_add_0_root_add_223_n25,
         DP_add_0_root_add_0_root_add_223_n23,
         DP_add_0_root_add_0_root_add_223_n22,
         DP_add_0_root_add_0_root_add_223_n21,
         DP_add_0_root_add_0_root_add_223_n19,
         DP_add_0_root_add_0_root_add_223_n17,
         DP_add_0_root_add_0_root_add_223_n16,
         DP_add_0_root_add_0_root_add_223_n14,
         DP_add_0_root_add_0_root_add_223_n13,
         DP_add_0_root_add_0_root_add_223_n12,
         DP_add_0_root_add_0_root_add_223_n11,
         DP_add_0_root_add_0_root_add_223_n10,
         DP_add_0_root_add_0_root_add_223_n9,
         DP_add_0_root_add_0_root_add_223_n8,
         DP_add_0_root_add_0_root_add_223_n7,
         DP_add_0_root_add_0_root_add_223_n6,
         DP_add_0_root_add_0_root_add_223_n5,
         DP_add_0_root_add_0_root_add_223_n4,
         DP_add_0_root_add_0_root_add_223_n3,
         DP_add_0_root_add_0_root_add_223_n2,
         DP_add_0_root_add_0_root_add_223_n1, DP_mult_205_n2341,
         DP_mult_205_n2340, DP_mult_205_n2339, DP_mult_205_n2338,
         DP_mult_205_n2337, DP_mult_205_n2336, DP_mult_205_n2335,
         DP_mult_205_n2334, DP_mult_205_n2333, DP_mult_205_n2332,
         DP_mult_205_n2331, DP_mult_205_n2330, DP_mult_205_n2329,
         DP_mult_205_n2328, DP_mult_205_n2327, DP_mult_205_n2326,
         DP_mult_205_n2325, DP_mult_205_n2324, DP_mult_205_n2323,
         DP_mult_205_n2322, DP_mult_205_n2321, DP_mult_205_n2320,
         DP_mult_205_n2319, DP_mult_205_n2318, DP_mult_205_n2317,
         DP_mult_205_n2316, DP_mult_205_n2315, DP_mult_205_n2314,
         DP_mult_205_n2313, DP_mult_205_n2312, DP_mult_205_n2311,
         DP_mult_205_n2310, DP_mult_205_n2309, DP_mult_205_n2308,
         DP_mult_205_n2307, DP_mult_205_n2306, DP_mult_205_n2305,
         DP_mult_205_n2304, DP_mult_205_n2303, DP_mult_205_n2302,
         DP_mult_205_n2301, DP_mult_205_n2300, DP_mult_205_n2299,
         DP_mult_205_n2298, DP_mult_205_n2297, DP_mult_205_n2296,
         DP_mult_205_n2295, DP_mult_205_n2294, DP_mult_205_n2293,
         DP_mult_205_n2292, DP_mult_205_n2291, DP_mult_205_n2290,
         DP_mult_205_n2289, DP_mult_205_n2288, DP_mult_205_n2287,
         DP_mult_205_n2286, DP_mult_205_n2285, DP_mult_205_n2284,
         DP_mult_205_n2283, DP_mult_205_n2282, DP_mult_205_n2281,
         DP_mult_205_n2280, DP_mult_205_n2279, DP_mult_205_n2278,
         DP_mult_205_n2277, DP_mult_205_n2276, DP_mult_205_n2275,
         DP_mult_205_n2274, DP_mult_205_n2273, DP_mult_205_n2272,
         DP_mult_205_n2271, DP_mult_205_n2270, DP_mult_205_n2269,
         DP_mult_205_n2268, DP_mult_205_n2267, DP_mult_205_n2266,
         DP_mult_205_n2265, DP_mult_205_n2264, DP_mult_205_n2263,
         DP_mult_205_n2262, DP_mult_205_n2261, DP_mult_205_n2260,
         DP_mult_205_n2259, DP_mult_205_n2258, DP_mult_205_n2257,
         DP_mult_205_n2256, DP_mult_205_n2255, DP_mult_205_n2254,
         DP_mult_205_n2253, DP_mult_205_n2252, DP_mult_205_n2251,
         DP_mult_205_n2250, DP_mult_205_n2249, DP_mult_205_n2248,
         DP_mult_205_n2247, DP_mult_205_n2246, DP_mult_205_n2245,
         DP_mult_205_n2244, DP_mult_205_n2243, DP_mult_205_n2242,
         DP_mult_205_n2241, DP_mult_205_n2240, DP_mult_205_n2239,
         DP_mult_205_n2238, DP_mult_205_n2237, DP_mult_205_n2236,
         DP_mult_205_n2235, DP_mult_205_n2234, DP_mult_205_n2233,
         DP_mult_205_n2232, DP_mult_205_n2231, DP_mult_205_n2230,
         DP_mult_205_n2229, DP_mult_205_n2228, DP_mult_205_n2227,
         DP_mult_205_n2226, DP_mult_205_n2225, DP_mult_205_n2224,
         DP_mult_205_n2223, DP_mult_205_n2222, DP_mult_205_n2221,
         DP_mult_205_n2220, DP_mult_205_n2219, DP_mult_205_n2218,
         DP_mult_205_n2217, DP_mult_205_n2216, DP_mult_205_n2215,
         DP_mult_205_n2214, DP_mult_205_n2213, DP_mult_205_n2212,
         DP_mult_205_n2211, DP_mult_205_n2210, DP_mult_205_n2209,
         DP_mult_205_n2208, DP_mult_205_n2207, DP_mult_205_n2206,
         DP_mult_205_n2205, DP_mult_205_n2204, DP_mult_205_n2203,
         DP_mult_205_n2202, DP_mult_205_n2201, DP_mult_205_n2200,
         DP_mult_205_n2199, DP_mult_205_n2198, DP_mult_205_n2197,
         DP_mult_205_n2196, DP_mult_205_n2195, DP_mult_205_n2194,
         DP_mult_205_n2193, DP_mult_205_n2192, DP_mult_205_n2191,
         DP_mult_205_n2190, DP_mult_205_n2189, DP_mult_205_n2188,
         DP_mult_205_n2187, DP_mult_205_n2186, DP_mult_205_n2185,
         DP_mult_205_n2184, DP_mult_205_n2183, DP_mult_205_n2182,
         DP_mult_205_n2181, DP_mult_205_n2180, DP_mult_205_n2179,
         DP_mult_205_n2178, DP_mult_205_n2177, DP_mult_205_n2176,
         DP_mult_205_n2175, DP_mult_205_n2174, DP_mult_205_n2173,
         DP_mult_205_n2172, DP_mult_205_n2171, DP_mult_205_n2170,
         DP_mult_205_n2169, DP_mult_205_n2168, DP_mult_205_n2167,
         DP_mult_205_n2166, DP_mult_205_n2165, DP_mult_205_n2164,
         DP_mult_205_n2163, DP_mult_205_n2162, DP_mult_205_n2161,
         DP_mult_205_n2160, DP_mult_205_n2159, DP_mult_205_n2158,
         DP_mult_205_n2157, DP_mult_205_n2156, DP_mult_205_n2155,
         DP_mult_205_n2154, DP_mult_205_n2153, DP_mult_205_n2152,
         DP_mult_205_n2151, DP_mult_205_n2150, DP_mult_205_n2149,
         DP_mult_205_n2148, DP_mult_205_n2147, DP_mult_205_n2146,
         DP_mult_205_n2145, DP_mult_205_n2144, DP_mult_205_n2143,
         DP_mult_205_n2142, DP_mult_205_n2141, DP_mult_205_n2140,
         DP_mult_205_n2139, DP_mult_205_n2138, DP_mult_205_n2137,
         DP_mult_205_n2136, DP_mult_205_n2135, DP_mult_205_n2134,
         DP_mult_205_n2133, DP_mult_205_n2132, DP_mult_205_n2131,
         DP_mult_205_n2130, DP_mult_205_n2129, DP_mult_205_n2128,
         DP_mult_205_n2127, DP_mult_205_n2126, DP_mult_205_n2125,
         DP_mult_205_n2124, DP_mult_205_n2123, DP_mult_205_n2122,
         DP_mult_205_n2121, DP_mult_205_n2120, DP_mult_205_n2119,
         DP_mult_205_n2118, DP_mult_205_n2117, DP_mult_205_n2116,
         DP_mult_205_n2115, DP_mult_205_n2114, DP_mult_205_n2113,
         DP_mult_205_n2112, DP_mult_205_n2111, DP_mult_205_n2110,
         DP_mult_205_n2109, DP_mult_205_n2108, DP_mult_205_n2107,
         DP_mult_205_n2106, DP_mult_205_n2105, DP_mult_205_n2104,
         DP_mult_205_n2103, DP_mult_205_n2102, DP_mult_205_n2101,
         DP_mult_205_n2100, DP_mult_205_n2099, DP_mult_205_n2098,
         DP_mult_205_n2097, DP_mult_205_n2096, DP_mult_205_n2095,
         DP_mult_205_n2094, DP_mult_205_n2093, DP_mult_205_n2092,
         DP_mult_205_n2091, DP_mult_205_n2090, DP_mult_205_n2089,
         DP_mult_205_n2088, DP_mult_205_n2087, DP_mult_205_n2086,
         DP_mult_205_n2085, DP_mult_205_n2084, DP_mult_205_n2083,
         DP_mult_205_n2082, DP_mult_205_n2081, DP_mult_205_n2080,
         DP_mult_205_n2079, DP_mult_205_n2078, DP_mult_205_n2077,
         DP_mult_205_n2076, DP_mult_205_n2075, DP_mult_205_n2074,
         DP_mult_205_n2073, DP_mult_205_n2072, DP_mult_205_n2071,
         DP_mult_205_n2070, DP_mult_205_n2069, DP_mult_205_n2068,
         DP_mult_205_n2067, DP_mult_205_n2066, DP_mult_205_n2065,
         DP_mult_205_n2064, DP_mult_205_n2063, DP_mult_205_n2062,
         DP_mult_205_n2061, DP_mult_205_n2060, DP_mult_205_n2059,
         DP_mult_205_n2058, DP_mult_205_n2057, DP_mult_205_n2056,
         DP_mult_205_n2055, DP_mult_205_n2054, DP_mult_205_n2053,
         DP_mult_205_n2052, DP_mult_205_n2051, DP_mult_205_n2050,
         DP_mult_205_n2049, DP_mult_205_n2048, DP_mult_205_n2047,
         DP_mult_205_n2046, DP_mult_205_n2045, DP_mult_205_n2044,
         DP_mult_205_n2043, DP_mult_205_n2042, DP_mult_205_n2041,
         DP_mult_205_n2040, DP_mult_205_n2039, DP_mult_205_n2038,
         DP_mult_205_n2037, DP_mult_205_n2036, DP_mult_205_n2035,
         DP_mult_205_n2034, DP_mult_205_n2033, DP_mult_205_n2032,
         DP_mult_205_n2031, DP_mult_205_n2030, DP_mult_205_n2029,
         DP_mult_205_n2028, DP_mult_205_n2027, DP_mult_205_n2026,
         DP_mult_205_n2025, DP_mult_205_n2024, DP_mult_205_n2023,
         DP_mult_205_n2022, DP_mult_205_n2021, DP_mult_205_n2020,
         DP_mult_205_n2019, DP_mult_205_n2018, DP_mult_205_n2017,
         DP_mult_205_n2016, DP_mult_205_n2015, DP_mult_205_n2014,
         DP_mult_205_n2013, DP_mult_205_n2012, DP_mult_205_n2011,
         DP_mult_205_n2010, DP_mult_205_n2009, DP_mult_205_n2008,
         DP_mult_205_n2007, DP_mult_205_n2006, DP_mult_205_n2005,
         DP_mult_205_n2004, DP_mult_205_n2003, DP_mult_205_n2002,
         DP_mult_205_n2001, DP_mult_205_n2000, DP_mult_205_n1999,
         DP_mult_205_n1998, DP_mult_205_n1997, DP_mult_205_n1996,
         DP_mult_205_n1995, DP_mult_205_n1994, DP_mult_205_n1993,
         DP_mult_205_n1992, DP_mult_205_n1991, DP_mult_205_n1990,
         DP_mult_205_n1989, DP_mult_205_n1988, DP_mult_205_n1987,
         DP_mult_205_n1986, DP_mult_205_n1985, DP_mult_205_n1984,
         DP_mult_205_n1983, DP_mult_205_n1982, DP_mult_205_n1981,
         DP_mult_205_n1980, DP_mult_205_n1979, DP_mult_205_n1978,
         DP_mult_205_n1977, DP_mult_205_n1976, DP_mult_205_n1975,
         DP_mult_205_n1974, DP_mult_205_n1973, DP_mult_205_n1972,
         DP_mult_205_n1971, DP_mult_205_n1970, DP_mult_205_n1969,
         DP_mult_205_n1968, DP_mult_205_n1967, DP_mult_205_n1966,
         DP_mult_205_n1965, DP_mult_205_n1964, DP_mult_205_n1963,
         DP_mult_205_n1962, DP_mult_205_n1961, DP_mult_205_n1960,
         DP_mult_205_n1959, DP_mult_205_n1958, DP_mult_205_n1957,
         DP_mult_205_n1956, DP_mult_205_n1955, DP_mult_205_n1954,
         DP_mult_205_n1953, DP_mult_205_n1952, DP_mult_205_n1951,
         DP_mult_205_n1950, DP_mult_205_n1949, DP_mult_205_n1948,
         DP_mult_205_n1947, DP_mult_205_n1946, DP_mult_205_n1945,
         DP_mult_205_n1944, DP_mult_205_n1943, DP_mult_205_n1942,
         DP_mult_205_n1941, DP_mult_205_n1940, DP_mult_205_n1939,
         DP_mult_205_n1938, DP_mult_205_n1937, DP_mult_205_n1936,
         DP_mult_205_n1935, DP_mult_205_n1934, DP_mult_205_n1933,
         DP_mult_205_n1932, DP_mult_205_n1931, DP_mult_205_n1930,
         DP_mult_205_n1929, DP_mult_205_n1817, DP_mult_205_n1816,
         DP_mult_205_n1815, DP_mult_205_n1814, DP_mult_205_n1813,
         DP_mult_205_n1812, DP_mult_205_n1811, DP_mult_205_n1810,
         DP_mult_205_n1809, DP_mult_205_n1808, DP_mult_205_n1781,
         DP_mult_205_n1780, DP_mult_205_n1779, DP_mult_205_n1778,
         DP_mult_205_n1777, DP_mult_205_n1776, DP_mult_205_n1775,
         DP_mult_205_n1774, DP_mult_205_n1773, DP_mult_205_n1772,
         DP_mult_205_n1771, DP_mult_205_n1770, DP_mult_205_n1769,
         DP_mult_205_n1768, DP_mult_205_n1767, DP_mult_205_n1766,
         DP_mult_205_n1765, DP_mult_205_n1764, DP_mult_205_n1763,
         DP_mult_205_n1762, DP_mult_205_n1761, DP_mult_205_n1760,
         DP_mult_205_n1759, DP_mult_205_n1758, DP_mult_205_n1757,
         DP_mult_205_n1756, DP_mult_205_n1755, DP_mult_205_n1754,
         DP_mult_205_n1753, DP_mult_205_n1752, DP_mult_205_n1751,
         DP_mult_205_n1750, DP_mult_205_n1749, DP_mult_205_n1748,
         DP_mult_205_n1747, DP_mult_205_n1746, DP_mult_205_n1745,
         DP_mult_205_n1744, DP_mult_205_n1743, DP_mult_205_n1742,
         DP_mult_205_n1741, DP_mult_205_n1740, DP_mult_205_n1739,
         DP_mult_205_n1738, DP_mult_205_n1737, DP_mult_205_n1736,
         DP_mult_205_n1735, DP_mult_205_n1734, DP_mult_205_n1733,
         DP_mult_205_n1732, DP_mult_205_n1731, DP_mult_205_n1730,
         DP_mult_205_n1729, DP_mult_205_n1728, DP_mult_205_n1727,
         DP_mult_205_n1726, DP_mult_205_n1725, DP_mult_205_n1724,
         DP_mult_205_n1723, DP_mult_205_n1722, DP_mult_205_n1721,
         DP_mult_205_n1720, DP_mult_205_n1719, DP_mult_205_n1718,
         DP_mult_205_n1717, DP_mult_205_n1716, DP_mult_205_n1715,
         DP_mult_205_n1714, DP_mult_205_n1713, DP_mult_205_n1712,
         DP_mult_205_n1711, DP_mult_205_n1710, DP_mult_205_n1709,
         DP_mult_205_n1708, DP_mult_205_n1707, DP_mult_205_n1706,
         DP_mult_205_n1705, DP_mult_205_n1704, DP_mult_205_n1703,
         DP_mult_205_n1702, DP_mult_205_n1701, DP_mult_205_n1700,
         DP_mult_205_n1699, DP_mult_205_n1698, DP_mult_205_n1697,
         DP_mult_205_n1696, DP_mult_205_n1695, DP_mult_205_n1694,
         DP_mult_205_n1693, DP_mult_205_n1692, DP_mult_205_n1691,
         DP_mult_205_n1690, DP_mult_205_n1689, DP_mult_205_n1688,
         DP_mult_205_n1687, DP_mult_205_n1686, DP_mult_205_n1685,
         DP_mult_205_n1684, DP_mult_205_n1683, DP_mult_205_n1682,
         DP_mult_205_n1681, DP_mult_205_n1680, DP_mult_205_n1679,
         DP_mult_205_n1678, DP_mult_205_n1677, DP_mult_205_n1676,
         DP_mult_205_n1675, DP_mult_205_n1674, DP_mult_205_n1673,
         DP_mult_205_n1672, DP_mult_205_n1671, DP_mult_205_n1670,
         DP_mult_205_n1669, DP_mult_205_n1668, DP_mult_205_n1667,
         DP_mult_205_n1666, DP_mult_205_n1665, DP_mult_205_n1664,
         DP_mult_205_n1663, DP_mult_205_n1662, DP_mult_205_n1661,
         DP_mult_205_n1660, DP_mult_205_n1659, DP_mult_205_n1658,
         DP_mult_205_n1657, DP_mult_205_n1656, DP_mult_205_n1655,
         DP_mult_205_n1654, DP_mult_205_n1653, DP_mult_205_n1652,
         DP_mult_205_n1651, DP_mult_205_n1650, DP_mult_205_n1649,
         DP_mult_205_n1648, DP_mult_205_n1647, DP_mult_205_n1646,
         DP_mult_205_n1645, DP_mult_205_n1644, DP_mult_205_n1643,
         DP_mult_205_n1642, DP_mult_205_n1641, DP_mult_205_n1640,
         DP_mult_205_n1639, DP_mult_205_n1638, DP_mult_205_n1637,
         DP_mult_205_n1636, DP_mult_205_n1635, DP_mult_205_n1634,
         DP_mult_205_n1633, DP_mult_205_n1632, DP_mult_205_n1631,
         DP_mult_205_n1630, DP_mult_205_n1629, DP_mult_205_n1628,
         DP_mult_205_n1627, DP_mult_205_n1626, DP_mult_205_n1625,
         DP_mult_205_n1624, DP_mult_205_n1623, DP_mult_205_n1622,
         DP_mult_205_n1621, DP_mult_205_n1620, DP_mult_205_n1619,
         DP_mult_205_n1618, DP_mult_205_n1617, DP_mult_205_n1616,
         DP_mult_205_n1615, DP_mult_205_n1614, DP_mult_205_n1613,
         DP_mult_205_n1612, DP_mult_205_n1611, DP_mult_205_n1610,
         DP_mult_205_n1609, DP_mult_205_n1608, DP_mult_205_n1607,
         DP_mult_205_n1606, DP_mult_205_n1605, DP_mult_205_n1604,
         DP_mult_205_n1603, DP_mult_205_n1602, DP_mult_205_n1601,
         DP_mult_205_n1600, DP_mult_205_n1599, DP_mult_205_n1598,
         DP_mult_205_n1597, DP_mult_205_n1596, DP_mult_205_n1595,
         DP_mult_205_n1594, DP_mult_205_n1593, DP_mult_205_n1592,
         DP_mult_205_n1591, DP_mult_205_n1590, DP_mult_205_n1589,
         DP_mult_205_n1588, DP_mult_205_n1587, DP_mult_205_n1586,
         DP_mult_205_n1585, DP_mult_205_n1584, DP_mult_205_n1583,
         DP_mult_205_n1582, DP_mult_205_n1581, DP_mult_205_n1580,
         DP_mult_205_n1579, DP_mult_205_n1578, DP_mult_205_n1577,
         DP_mult_205_n1576, DP_mult_205_n1575, DP_mult_205_n1574,
         DP_mult_205_n1573, DP_mult_205_n1572, DP_mult_205_n1571,
         DP_mult_205_n1570, DP_mult_205_n1569, DP_mult_205_n1568,
         DP_mult_205_n1567, DP_mult_205_n1566, DP_mult_205_n1565,
         DP_mult_205_n1564, DP_mult_205_n1563, DP_mult_205_n1562,
         DP_mult_205_n1561, DP_mult_205_n1560, DP_mult_205_n1559,
         DP_mult_205_n1558, DP_mult_205_n1557, DP_mult_205_n1556,
         DP_mult_205_n1555, DP_mult_205_n1554, DP_mult_205_n1553,
         DP_mult_205_n1552, DP_mult_205_n1551, DP_mult_205_n1550,
         DP_mult_205_n1549, DP_mult_205_n1548, DP_mult_205_n1547,
         DP_mult_205_n1546, DP_mult_205_n1545, DP_mult_205_n1544,
         DP_mult_205_n1543, DP_mult_205_n1542, DP_mult_205_n1541,
         DP_mult_205_n1540, DP_mult_205_n1539, DP_mult_205_n1538,
         DP_mult_205_n1537, DP_mult_205_n1536, DP_mult_205_n1535,
         DP_mult_205_n1534, DP_mult_205_n1533, DP_mult_205_n1532,
         DP_mult_205_n1531, DP_mult_205_n1530, DP_mult_205_n1529,
         DP_mult_205_n1528, DP_mult_205_n1527, DP_mult_205_n1526,
         DP_mult_205_n1525, DP_mult_205_n1524, DP_mult_205_n1523,
         DP_mult_205_n1522, DP_mult_205_n1521, DP_mult_205_n1520,
         DP_mult_205_n1519, DP_mult_205_n1518, DP_mult_205_n1517,
         DP_mult_205_n1516, DP_mult_205_n1515, DP_mult_205_n1514,
         DP_mult_205_n1513, DP_mult_205_n1512, DP_mult_205_n1511,
         DP_mult_205_n1510, DP_mult_205_n1509, DP_mult_205_n1508,
         DP_mult_205_n1507, DP_mult_205_n1506, DP_mult_205_n1505,
         DP_mult_205_n1504, DP_mult_205_n1503, DP_mult_205_n1502,
         DP_mult_205_n1501, DP_mult_205_n1500, DP_mult_205_n1499,
         DP_mult_205_n1498, DP_mult_205_n1497, DP_mult_205_n1496,
         DP_mult_205_n1495, DP_mult_205_n1494, DP_mult_205_n1493,
         DP_mult_205_n1492, DP_mult_205_n1491, DP_mult_205_n1490,
         DP_mult_205_n1489, DP_mult_205_n1488, DP_mult_205_n1487,
         DP_mult_205_n1486, DP_mult_205_n1485, DP_mult_205_n1484,
         DP_mult_205_n1483, DP_mult_205_n1482, DP_mult_205_n1481,
         DP_mult_205_n1480, DP_mult_205_n1479, DP_mult_205_n1478,
         DP_mult_205_n1477, DP_mult_205_n1476, DP_mult_205_n1475,
         DP_mult_205_n1474, DP_mult_205_n1473, DP_mult_205_n1472,
         DP_mult_205_n1471, DP_mult_205_n1470, DP_mult_205_n1469,
         DP_mult_205_n1468, DP_mult_205_n1467, DP_mult_205_n1466,
         DP_mult_205_n1465, DP_mult_205_n1464, DP_mult_205_n1463,
         DP_mult_205_n1462, DP_mult_205_n1461, DP_mult_205_n1460,
         DP_mult_205_n1459, DP_mult_205_n1458, DP_mult_205_n1457,
         DP_mult_205_n1456, DP_mult_205_n1455, DP_mult_205_n1454,
         DP_mult_205_n1453, DP_mult_205_n1452, DP_mult_205_n1451,
         DP_mult_205_n1450, DP_mult_205_n1449, DP_mult_205_n1448,
         DP_mult_205_n1447, DP_mult_205_n1446, DP_mult_205_n1445,
         DP_mult_205_n1444, DP_mult_205_n1443, DP_mult_205_n1442,
         DP_mult_205_n1441, DP_mult_205_n1440, DP_mult_205_n1439,
         DP_mult_205_n1438, DP_mult_205_n1437, DP_mult_205_n1436,
         DP_mult_205_n1435, DP_mult_205_n1434, DP_mult_205_n1433,
         DP_mult_205_n1432, DP_mult_205_n1431, DP_mult_205_n1430,
         DP_mult_205_n1429, DP_mult_205_n1428, DP_mult_205_n1427,
         DP_mult_205_n1426, DP_mult_205_n1425, DP_mult_205_n1424,
         DP_mult_205_n1423, DP_mult_205_n1422, DP_mult_205_n1421,
         DP_mult_205_n1420, DP_mult_205_n1419, DP_mult_205_n1418,
         DP_mult_205_n1417, DP_mult_205_n1416, DP_mult_205_n1415,
         DP_mult_205_n1414, DP_mult_205_n1413, DP_mult_205_n1412,
         DP_mult_205_n1411, DP_mult_205_n1410, DP_mult_205_n1409,
         DP_mult_205_n1408, DP_mult_205_n1407, DP_mult_205_n1406,
         DP_mult_205_n1405, DP_mult_205_n1404, DP_mult_205_n1403,
         DP_mult_205_n1402, DP_mult_205_n1401, DP_mult_205_n1400,
         DP_mult_205_n1399, DP_mult_205_n1398, DP_mult_205_n1397,
         DP_mult_205_n1396, DP_mult_205_n1395, DP_mult_205_n1394,
         DP_mult_205_n1393, DP_mult_205_n1392, DP_mult_205_n1391,
         DP_mult_205_n1390, DP_mult_205_n1389, DP_mult_205_n1388,
         DP_mult_205_n1387, DP_mult_205_n1386, DP_mult_205_n1385,
         DP_mult_205_n1384, DP_mult_205_n1383, DP_mult_205_n1382,
         DP_mult_205_n1381, DP_mult_205_n1380, DP_mult_205_n1379,
         DP_mult_205_n1378, DP_mult_205_n1377, DP_mult_205_n1376,
         DP_mult_205_n1375, DP_mult_205_n1374, DP_mult_205_n1373,
         DP_mult_205_n1372, DP_mult_205_n1371, DP_mult_205_n1370,
         DP_mult_205_n1369, DP_mult_205_n1368, DP_mult_205_n1367,
         DP_mult_205_n1366, DP_mult_205_n1365, DP_mult_205_n1364,
         DP_mult_205_n1363, DP_mult_205_n1362, DP_mult_205_n1361,
         DP_mult_205_n1360, DP_mult_205_n1359, DP_mult_205_n1358,
         DP_mult_205_n1357, DP_mult_205_n1356, DP_mult_205_n1355,
         DP_mult_205_n1354, DP_mult_205_n1353, DP_mult_205_n1352,
         DP_mult_205_n1351, DP_mult_205_n1350, DP_mult_205_n1349,
         DP_mult_205_n1348, DP_mult_205_n1347, DP_mult_205_n1346,
         DP_mult_205_n1345, DP_mult_205_n1344, DP_mult_205_n1343,
         DP_mult_205_n1342, DP_mult_205_n1341, DP_mult_205_n1340,
         DP_mult_205_n1339, DP_mult_205_n1338, DP_mult_205_n1337,
         DP_mult_205_n1336, DP_mult_205_n1335, DP_mult_205_n1334,
         DP_mult_205_n1333, DP_mult_205_n1332, DP_mult_205_n1331,
         DP_mult_205_n1330, DP_mult_205_n1329, DP_mult_205_n1328,
         DP_mult_205_n1327, DP_mult_205_n1326, DP_mult_205_n1325,
         DP_mult_205_n1324, DP_mult_205_n1323, DP_mult_205_n1322,
         DP_mult_205_n1321, DP_mult_205_n1320, DP_mult_205_n1319,
         DP_mult_205_n1318, DP_mult_205_n1317, DP_mult_205_n1316,
         DP_mult_205_n1315, DP_mult_205_n1314, DP_mult_205_n1313,
         DP_mult_205_n1312, DP_mult_205_n1311, DP_mult_205_n1310,
         DP_mult_205_n1309, DP_mult_205_n1308, DP_mult_205_n1307,
         DP_mult_205_n1306, DP_mult_205_n1305, DP_mult_205_n1304,
         DP_mult_205_n1303, DP_mult_205_n1302, DP_mult_205_n1301,
         DP_mult_205_n1300, DP_mult_205_n1299, DP_mult_205_n1298,
         DP_mult_205_n1297, DP_mult_205_n1296, DP_mult_205_n1295,
         DP_mult_205_n1294, DP_mult_205_n1293, DP_mult_205_n1292,
         DP_mult_205_n1291, DP_mult_205_n1290, DP_mult_205_n1289,
         DP_mult_205_n1288, DP_mult_205_n1287, DP_mult_205_n1286,
         DP_mult_205_n1285, DP_mult_205_n1284, DP_mult_205_n1283,
         DP_mult_205_n1282, DP_mult_205_n1281, DP_mult_205_n1280,
         DP_mult_205_n1279, DP_mult_205_n1278, DP_mult_205_n1277,
         DP_mult_205_n1276, DP_mult_205_n1275, DP_mult_205_n1274,
         DP_mult_205_n1273, DP_mult_205_n1272, DP_mult_205_n1271,
         DP_mult_205_n1270, DP_mult_205_n1269, DP_mult_205_n1268,
         DP_mult_205_n1267, DP_mult_205_n1266, DP_mult_205_n1265,
         DP_mult_205_n1264, DP_mult_205_n1263, DP_mult_205_n1262,
         DP_mult_205_n1261, DP_mult_205_n1260, DP_mult_205_n1259,
         DP_mult_205_n1258, DP_mult_205_n1257, DP_mult_205_n1256,
         DP_mult_205_n1255, DP_mult_205_n1254, DP_mult_205_n1253,
         DP_mult_205_n1252, DP_mult_205_n1251, DP_mult_205_n1250,
         DP_mult_205_n1249, DP_mult_205_n1248, DP_mult_205_n1247,
         DP_mult_205_n1246, DP_mult_205_n1245, DP_mult_205_n1244,
         DP_mult_205_n1243, DP_mult_205_n1242, DP_mult_205_n1241,
         DP_mult_205_n1240, DP_mult_205_n1239, DP_mult_205_n1238,
         DP_mult_205_n1237, DP_mult_205_n1236, DP_mult_205_n1235,
         DP_mult_205_n1234, DP_mult_205_n1233, DP_mult_205_n1232,
         DP_mult_205_n1231, DP_mult_205_n1230, DP_mult_205_n1229,
         DP_mult_205_n1228, DP_mult_205_n1227, DP_mult_205_n1226,
         DP_mult_205_n1225, DP_mult_205_n1224, DP_mult_205_n1223,
         DP_mult_205_n1222, DP_mult_205_n1221, DP_mult_205_n1220,
         DP_mult_205_n1219, DP_mult_205_n1218, DP_mult_205_n1217,
         DP_mult_205_n1216, DP_mult_205_n1215, DP_mult_205_n1214,
         DP_mult_205_n1213, DP_mult_205_n1212, DP_mult_205_n1211,
         DP_mult_205_n1210, DP_mult_205_n1209, DP_mult_205_n1208,
         DP_mult_205_n1207, DP_mult_205_n1206, DP_mult_205_n1205,
         DP_mult_205_n1204, DP_mult_205_n1203, DP_mult_205_n1202,
         DP_mult_205_n1201, DP_mult_205_n1200, DP_mult_205_n1199,
         DP_mult_205_n1198, DP_mult_205_n1197, DP_mult_205_n1196,
         DP_mult_205_n1195, DP_mult_205_n1194, DP_mult_205_n1193,
         DP_mult_205_n1192, DP_mult_205_n1191, DP_mult_205_n1190,
         DP_mult_205_n1189, DP_mult_205_n1188, DP_mult_205_n1187,
         DP_mult_205_n1186, DP_mult_205_n1185, DP_mult_205_n1184,
         DP_mult_205_n1183, DP_mult_205_n1182, DP_mult_205_n1181,
         DP_mult_205_n1180, DP_mult_205_n1179, DP_mult_205_n1178,
         DP_mult_205_n1177, DP_mult_205_n1176, DP_mult_205_n1175,
         DP_mult_205_n1174, DP_mult_205_n1173, DP_mult_205_n1172,
         DP_mult_205_n1171, DP_mult_205_n1170, DP_mult_205_n1169,
         DP_mult_205_n1168, DP_mult_205_n1167, DP_mult_205_n1166,
         DP_mult_205_n1165, DP_mult_205_n1164, DP_mult_205_n1163,
         DP_mult_205_n1162, DP_mult_205_n1161, DP_mult_205_n1160,
         DP_mult_205_n1159, DP_mult_205_n1158, DP_mult_205_n1157,
         DP_mult_205_n1156, DP_mult_205_n1155, DP_mult_205_n1154,
         DP_mult_205_n1153, DP_mult_205_n1152, DP_mult_205_n1151,
         DP_mult_205_n1150, DP_mult_205_n1149, DP_mult_205_n1148,
         DP_mult_205_n1147, DP_mult_205_n1146, DP_mult_205_n1145,
         DP_mult_205_n1144, DP_mult_205_n1143, DP_mult_205_n1142,
         DP_mult_205_n1141, DP_mult_205_n1140, DP_mult_205_n1139,
         DP_mult_205_n1138, DP_mult_205_n1137, DP_mult_205_n1136,
         DP_mult_205_n1135, DP_mult_205_n1134, DP_mult_205_n1133,
         DP_mult_205_n1132, DP_mult_205_n1131, DP_mult_205_n1130,
         DP_mult_205_n1129, DP_mult_205_n1128, DP_mult_205_n1127,
         DP_mult_205_n1126, DP_mult_205_n1125, DP_mult_205_n1124,
         DP_mult_205_n1123, DP_mult_205_n1122, DP_mult_205_n1121,
         DP_mult_205_n1120, DP_mult_205_n1119, DP_mult_205_n1118,
         DP_mult_205_n1117, DP_mult_205_n1116, DP_mult_205_n1115,
         DP_mult_205_n1114, DP_mult_205_n1113, DP_mult_205_n1112,
         DP_mult_205_n1111, DP_mult_205_n1110, DP_mult_205_n1109,
         DP_mult_205_n1108, DP_mult_205_n1107, DP_mult_205_n1106,
         DP_mult_205_n1105, DP_mult_205_n1104, DP_mult_205_n1103,
         DP_mult_205_n1102, DP_mult_205_n1101, DP_mult_205_n1100,
         DP_mult_205_n1099, DP_mult_205_n1098, DP_mult_205_n1097,
         DP_mult_205_n1096, DP_mult_205_n1095, DP_mult_205_n1094,
         DP_mult_205_n1093, DP_mult_205_n1092, DP_mult_205_n1091,
         DP_mult_205_n1090, DP_mult_205_n1089, DP_mult_205_n1088,
         DP_mult_205_n1087, DP_mult_205_n1086, DP_mult_205_n1085,
         DP_mult_205_n1084, DP_mult_205_n1083, DP_mult_205_n1082,
         DP_mult_205_n1081, DP_mult_205_n1080, DP_mult_205_n1079,
         DP_mult_205_n1078, DP_mult_205_n1077, DP_mult_205_n1076,
         DP_mult_205_n1075, DP_mult_205_n1074, DP_mult_205_n1073,
         DP_mult_205_n1072, DP_mult_205_n1071, DP_mult_205_n1070,
         DP_mult_205_n1069, DP_mult_205_n1068, DP_mult_205_n1067,
         DP_mult_205_n1066, DP_mult_205_n1065, DP_mult_205_n1064,
         DP_mult_205_n1063, DP_mult_205_n1062, DP_mult_205_n1061,
         DP_mult_205_n1060, DP_mult_205_n1059, DP_mult_205_n1058,
         DP_mult_205_n1057, DP_mult_205_n1056, DP_mult_205_n1055,
         DP_mult_205_n1054, DP_mult_205_n1053, DP_mult_205_n1052,
         DP_mult_205_n1051, DP_mult_205_n1050, DP_mult_205_n1049,
         DP_mult_205_n1048, DP_mult_205_n1047, DP_mult_205_n1046,
         DP_mult_205_n1045, DP_mult_205_n1044, DP_mult_205_n1043,
         DP_mult_205_n1042, DP_mult_205_n1041, DP_mult_205_n1040,
         DP_mult_205_n1039, DP_mult_205_n1038, DP_mult_205_n1037,
         DP_mult_205_n1036, DP_mult_205_n1035, DP_mult_205_n1034,
         DP_mult_205_n1033, DP_mult_205_n1032, DP_mult_205_n1031,
         DP_mult_205_n1030, DP_mult_205_n1029, DP_mult_205_n1028,
         DP_mult_205_n1027, DP_mult_205_n1026, DP_mult_205_n1025,
         DP_mult_205_n1024, DP_mult_205_n1023, DP_mult_205_n1022,
         DP_mult_205_n1021, DP_mult_205_n1020, DP_mult_205_n1019,
         DP_mult_205_n1018, DP_mult_205_n1017, DP_mult_205_n1016,
         DP_mult_205_n1015, DP_mult_205_n1014, DP_mult_205_n1013,
         DP_mult_205_n1012, DP_mult_205_n1011, DP_mult_205_n1010,
         DP_mult_205_n1009, DP_mult_205_n1008, DP_mult_205_n1007,
         DP_mult_205_n1006, DP_mult_205_n1005, DP_mult_205_n1004,
         DP_mult_205_n1003, DP_mult_205_n1002, DP_mult_205_n1001,
         DP_mult_205_n1000, DP_mult_205_n999, DP_mult_205_n998,
         DP_mult_205_n997, DP_mult_205_n996, DP_mult_205_n995,
         DP_mult_205_n994, DP_mult_205_n993, DP_mult_205_n992,
         DP_mult_205_n991, DP_mult_205_n990, DP_mult_205_n989,
         DP_mult_205_n988, DP_mult_205_n987, DP_mult_205_n986,
         DP_mult_205_n985, DP_mult_205_n984, DP_mult_205_n983,
         DP_mult_205_n982, DP_mult_205_n981, DP_mult_205_n980,
         DP_mult_205_n979, DP_mult_205_n978, DP_mult_205_n977,
         DP_mult_205_n976, DP_mult_205_n975, DP_mult_205_n974,
         DP_mult_205_n973, DP_mult_205_n972, DP_mult_205_n971,
         DP_mult_205_n970, DP_mult_205_n969, DP_mult_205_n968,
         DP_mult_205_n967, DP_mult_205_n966, DP_mult_205_n965,
         DP_mult_205_n964, DP_mult_205_n963, DP_mult_205_n962,
         DP_mult_205_n961, DP_mult_205_n959, DP_mult_205_n958,
         DP_mult_205_n957, DP_mult_205_n956, DP_mult_205_n955,
         DP_mult_205_n954, DP_mult_205_n953, DP_mult_205_n952,
         DP_mult_205_n951, DP_mult_205_n950, DP_mult_205_n949,
         DP_mult_205_n948, DP_mult_205_n947, DP_mult_205_n946,
         DP_mult_205_n945, DP_mult_205_n944, DP_mult_205_n943,
         DP_mult_205_n942, DP_mult_205_n941, DP_mult_205_n940,
         DP_mult_205_n939, DP_mult_205_n938, DP_mult_205_n937,
         DP_mult_205_n936, DP_mult_205_n935, DP_mult_205_n934,
         DP_mult_205_n933, DP_mult_205_n932, DP_mult_205_n931,
         DP_mult_205_n930, DP_mult_205_n929, DP_mult_205_n928,
         DP_mult_205_n927, DP_mult_205_n926, DP_mult_205_n925,
         DP_mult_205_n924, DP_mult_205_n923, DP_mult_205_n922,
         DP_mult_205_n921, DP_mult_205_n920, DP_mult_205_n919,
         DP_mult_205_n918, DP_mult_205_n917, DP_mult_205_n916,
         DP_mult_205_n915, DP_mult_205_n914, DP_mult_205_n913,
         DP_mult_205_n912, DP_mult_205_n911, DP_mult_205_n910,
         DP_mult_205_n909, DP_mult_205_n908, DP_mult_205_n907,
         DP_mult_205_n906, DP_mult_205_n905, DP_mult_205_n904,
         DP_mult_205_n903, DP_mult_205_n902, DP_mult_205_n901,
         DP_mult_205_n900, DP_mult_205_n899, DP_mult_205_n898,
         DP_mult_205_n897, DP_mult_205_n896, DP_mult_205_n895,
         DP_mult_205_n894, DP_mult_205_n893, DP_mult_205_n892,
         DP_mult_205_n891, DP_mult_205_n890, DP_mult_205_n889,
         DP_mult_205_n888, DP_mult_205_n887, DP_mult_205_n886,
         DP_mult_205_n885, DP_mult_205_n884, DP_mult_205_n883,
         DP_mult_205_n882, DP_mult_205_n881, DP_mult_205_n880,
         DP_mult_205_n879, DP_mult_205_n878, DP_mult_205_n877,
         DP_mult_205_n876, DP_mult_205_n875, DP_mult_205_n874,
         DP_mult_205_n873, DP_mult_205_n872, DP_mult_205_n871,
         DP_mult_205_n870, DP_mult_205_n869, DP_mult_205_n868,
         DP_mult_205_n867, DP_mult_205_n866, DP_mult_205_n865,
         DP_mult_205_n864, DP_mult_205_n863, DP_mult_205_n862,
         DP_mult_205_n861, DP_mult_205_n860, DP_mult_205_n859,
         DP_mult_205_n858, DP_mult_205_n857, DP_mult_205_n856,
         DP_mult_205_n855, DP_mult_205_n854, DP_mult_205_n853,
         DP_mult_205_n852, DP_mult_205_n851, DP_mult_205_n850,
         DP_mult_205_n849, DP_mult_205_n848, DP_mult_205_n847,
         DP_mult_205_n846, DP_mult_205_n845, DP_mult_205_n844,
         DP_mult_205_n843, DP_mult_205_n842, DP_mult_205_n841,
         DP_mult_205_n840, DP_mult_205_n839, DP_mult_205_n838,
         DP_mult_205_n837, DP_mult_205_n836, DP_mult_205_n835,
         DP_mult_205_n834, DP_mult_205_n833, DP_mult_205_n832,
         DP_mult_205_n831, DP_mult_205_n830, DP_mult_205_n829,
         DP_mult_205_n828, DP_mult_205_n827, DP_mult_205_n826,
         DP_mult_205_n825, DP_mult_205_n824, DP_mult_205_n823,
         DP_mult_205_n822, DP_mult_205_n821, DP_mult_205_n820,
         DP_mult_205_n819, DP_mult_205_n818, DP_mult_205_n817,
         DP_mult_205_n816, DP_mult_205_n815, DP_mult_205_n814,
         DP_mult_205_n813, DP_mult_205_n812, DP_mult_205_n811,
         DP_mult_205_n810, DP_mult_205_n809, DP_mult_205_n808,
         DP_mult_205_n807, DP_mult_205_n806, DP_mult_205_n805,
         DP_mult_205_n804, DP_mult_205_n803, DP_mult_205_n802,
         DP_mult_205_n801, DP_mult_205_n800, DP_mult_205_n799,
         DP_mult_205_n798, DP_mult_205_n797, DP_mult_205_n796,
         DP_mult_205_n795, DP_mult_205_n794, DP_mult_205_n793,
         DP_mult_205_n792, DP_mult_205_n791, DP_mult_205_n790,
         DP_mult_205_n789, DP_mult_205_n788, DP_mult_205_n787,
         DP_mult_205_n786, DP_mult_205_n785, DP_mult_205_n784,
         DP_mult_205_n783, DP_mult_205_n782, DP_mult_205_n781,
         DP_mult_205_n780, DP_mult_205_n779, DP_mult_205_n778,
         DP_mult_205_n777, DP_mult_205_n776, DP_mult_205_n775,
         DP_mult_205_n774, DP_mult_205_n773, DP_mult_205_n772,
         DP_mult_205_n771, DP_mult_205_n770, DP_mult_205_n769,
         DP_mult_205_n768, DP_mult_205_n767, DP_mult_205_n766,
         DP_mult_205_n765, DP_mult_205_n764, DP_mult_205_n763,
         DP_mult_205_n762, DP_mult_205_n761, DP_mult_205_n760,
         DP_mult_205_n759, DP_mult_205_n758, DP_mult_205_n757,
         DP_mult_205_n756, DP_mult_205_n755, DP_mult_205_n754,
         DP_mult_205_n753, DP_mult_205_n752, DP_mult_205_n751,
         DP_mult_205_n750, DP_mult_205_n749, DP_mult_205_n748,
         DP_mult_205_n747, DP_mult_205_n746, DP_mult_205_n745,
         DP_mult_205_n744, DP_mult_205_n743, DP_mult_205_n742,
         DP_mult_205_n741, DP_mult_205_n740, DP_mult_205_n739,
         DP_mult_205_n738, DP_mult_205_n737, DP_mult_205_n736,
         DP_mult_205_n735, DP_mult_205_n734, DP_mult_205_n733,
         DP_mult_205_n732, DP_mult_205_n731, DP_mult_205_n730,
         DP_mult_205_n729, DP_mult_205_n728, DP_mult_205_n727,
         DP_mult_205_n726, DP_mult_205_n725, DP_mult_205_n724,
         DP_mult_205_n723, DP_mult_205_n722, DP_mult_205_n721,
         DP_mult_205_n720, DP_mult_205_n719, DP_mult_205_n718,
         DP_mult_205_n717, DP_mult_205_n716, DP_mult_205_n715,
         DP_mult_205_n714, DP_mult_205_n713, DP_mult_205_n712,
         DP_mult_205_n711, DP_mult_205_n710, DP_mult_205_n709,
         DP_mult_205_n708, DP_mult_205_n707, DP_mult_205_n706,
         DP_mult_205_n705, DP_mult_205_n704, DP_mult_205_n703,
         DP_mult_205_n702, DP_mult_205_n701, DP_mult_205_n700,
         DP_mult_205_n699, DP_mult_205_n698, DP_mult_205_n697,
         DP_mult_205_n696, DP_mult_205_n695, DP_mult_205_n694,
         DP_mult_205_n693, DP_mult_205_n692, DP_mult_205_n691,
         DP_mult_205_n690, DP_mult_205_n689, DP_mult_205_n688,
         DP_mult_205_n687, DP_mult_205_n686, DP_mult_205_n685,
         DP_mult_205_n684, DP_mult_205_n683, DP_mult_205_n682,
         DP_mult_205_n681, DP_mult_205_n680, DP_mult_205_n679,
         DP_mult_205_n678, DP_mult_205_n677, DP_mult_205_n676,
         DP_mult_205_n675, DP_mult_205_n668, DP_mult_205_n666,
         DP_mult_205_n663, DP_mult_205_n662, DP_mult_205_n657,
         DP_mult_205_n646, DP_mult_205_n645, DP_mult_205_n644,
         DP_mult_205_n643, DP_mult_205_n638, DP_mult_205_n637,
         DP_mult_205_n636, DP_mult_205_n635, DP_mult_205_n634,
         DP_mult_205_n633, DP_mult_205_n632, DP_mult_205_n631,
         DP_mult_205_n630, DP_mult_205_n629, DP_mult_205_n628,
         DP_mult_205_n627, DP_mult_205_n626, DP_mult_205_n625,
         DP_mult_205_n620, DP_mult_205_n611, DP_mult_205_n610,
         DP_mult_205_n609, DP_mult_205_n600, DP_mult_205_n599,
         DP_mult_205_n598, DP_mult_205_n597, DP_mult_205_n596,
         DP_mult_205_n595, DP_mult_205_n594, DP_mult_205_n593,
         DP_mult_205_n592, DP_mult_205_n591, DP_mult_205_n590,
         DP_mult_205_n589, DP_mult_205_n588, DP_mult_205_n583,
         DP_mult_205_n582, DP_mult_205_n581, DP_mult_205_n572,
         DP_mult_205_n571, DP_mult_205_n570, DP_mult_205_n569,
         DP_mult_205_n568, DP_mult_205_n567, DP_mult_205_n565,
         DP_mult_205_n564, DP_mult_205_n563, DP_mult_205_n562,
         DP_mult_205_n561, DP_mult_205_n560, DP_mult_205_n559,
         DP_mult_205_n558, DP_mult_205_n555, DP_mult_205_n554,
         DP_mult_205_n553, DP_mult_205_n552, DP_mult_205_n551,
         DP_mult_205_n550, DP_mult_205_n547, DP_mult_205_n546,
         DP_mult_205_n545, DP_mult_205_n544, DP_mult_205_n543,
         DP_mult_205_n542, DP_mult_205_n541, DP_mult_205_n540,
         DP_mult_205_n539, DP_mult_205_n538, DP_mult_205_n537,
         DP_mult_205_n536, DP_mult_205_n535, DP_mult_205_n534,
         DP_mult_205_n533, DP_mult_205_n532, DP_mult_205_n531,
         DP_mult_205_n526, DP_mult_205_n525, DP_mult_205_n524,
         DP_mult_205_n522, DP_mult_205_n521, DP_mult_205_n520,
         DP_mult_205_n517, DP_mult_205_n516, DP_mult_205_n515,
         DP_mult_205_n514, DP_mult_205_n513, DP_mult_205_n512,
         DP_mult_205_n511, DP_mult_205_n508, DP_mult_205_n507,
         DP_mult_205_n506, DP_mult_205_n505, DP_mult_205_n504,
         DP_mult_205_n503, DP_mult_205_n502, DP_mult_205_n501,
         DP_mult_205_n499, DP_mult_205_n498, DP_mult_205_n497,
         DP_mult_205_n496, DP_mult_205_n495, DP_mult_205_n492,
         DP_mult_205_n491, DP_mult_205_n490, DP_mult_205_n489,
         DP_mult_205_n488, DP_mult_205_n487, DP_mult_205_n486,
         DP_mult_205_n483, DP_mult_205_n481, DP_mult_205_n480,
         DP_mult_205_n479, DP_mult_205_n478, DP_mult_205_n477,
         DP_mult_205_n476, DP_mult_205_n475, DP_mult_205_n474,
         DP_mult_205_n472, DP_mult_205_n468, DP_mult_205_n467,
         DP_mult_205_n466, DP_mult_205_n465, DP_mult_205_n464,
         DP_mult_205_n463, DP_mult_205_n462, DP_mult_205_n461,
         DP_mult_205_n459, DP_mult_205_n457, DP_mult_205_n456,
         DP_mult_205_n455, DP_mult_205_n454, DP_mult_205_n453,
         DP_mult_205_n452, DP_mult_205_n451, DP_mult_205_n450,
         DP_mult_205_n448, DP_mult_205_n445, DP_mult_205_n439,
         DP_mult_205_n438, DP_mult_205_n437, DP_mult_205_n436,
         DP_mult_205_n435, DP_mult_205_n434, DP_mult_205_n432,
         DP_mult_205_n431, DP_mult_205_n430, DP_mult_205_n429,
         DP_mult_205_n428, DP_mult_205_n427, DP_mult_205_n426,
         DP_mult_205_n423, DP_mult_205_n422, DP_mult_205_n421,
         DP_mult_205_n420, DP_mult_205_n419, DP_mult_205_n418,
         DP_mult_205_n416, DP_mult_205_n412, DP_mult_205_n411,
         DP_mult_205_n410, DP_mult_205_n409, DP_mult_205_n407,
         DP_mult_205_n405, DP_mult_205_n402, DP_mult_205_n401,
         DP_mult_205_n400, DP_mult_205_n399, DP_mult_205_n398,
         DP_mult_205_n397, DP_mult_205_n396, DP_mult_205_n394,
         DP_mult_205_n390, DP_mult_205_n389, DP_mult_205_n388,
         DP_mult_205_n387, DP_mult_205_n384, DP_mult_205_n383,
         DP_mult_205_n382, DP_mult_205_n381, DP_mult_205_n380,
         DP_mult_205_n379, DP_mult_205_n378, DP_mult_205_n376,
         DP_mult_205_n372, DP_mult_205_n371, DP_mult_205_n370,
         DP_mult_205_n369, DP_mult_205_n367, DP_mult_205_n365,
         DP_mult_205_n364, DP_mult_205_n363, DP_mult_205_n362,
         DP_mult_205_n361, DP_mult_205_n360, DP_mult_205_n359,
         DP_mult_205_n356, DP_mult_205_n355, DP_mult_205_n354,
         DP_mult_205_n353, DP_mult_205_n352, DP_mult_205_n350,
         DP_mult_205_n348, DP_mult_205_n347, DP_mult_205_n346,
         DP_mult_205_n345, DP_mult_205_n344, DP_mult_205_n343,
         DP_mult_205_n342, DP_mult_205_n341, DP_mult_205_n339,
         DP_mult_205_n337, DP_mult_205_n336, DP_mult_205_n335,
         DP_mult_205_n334, DP_mult_205_n333, DP_mult_205_n332,
         DP_mult_205_n327, DP_mult_205_n326, DP_mult_205_n325,
         DP_mult_205_n320, DP_mult_205_n319, DP_mult_205_n318,
         DP_mult_205_n317, DP_mult_205_n316, DP_mult_205_n315,
         DP_mult_205_n314, DP_mult_205_n313, DP_mult_205_n312,
         DP_mult_205_n311, DP_mult_205_n310, DP_mult_205_n309,
         DP_mult_205_n308, DP_mult_205_n307, DP_mult_205_n306,
         DP_mult_205_n305, DP_mult_205_n304, DP_mult_205_n303,
         DP_mult_205_n302, DP_mult_205_n301, DP_mult_205_n293,
         DP_mult_205_n289, DP_mult_205_n287, DP_mult_205_n283,
         DP_mult_205_n279, DP_mult_205_n277, DP_mult_205_n259,
         DP_mult_205_n251, DP_mult_204_n2395, DP_mult_204_n2394,
         DP_mult_204_n2393, DP_mult_204_n2392, DP_mult_204_n2391,
         DP_mult_204_n2390, DP_mult_204_n2389, DP_mult_204_n2388,
         DP_mult_204_n2387, DP_mult_204_n2386, DP_mult_204_n2385,
         DP_mult_204_n2384, DP_mult_204_n2383, DP_mult_204_n2382,
         DP_mult_204_n2381, DP_mult_204_n2380, DP_mult_204_n2379,
         DP_mult_204_n2378, DP_mult_204_n2377, DP_mult_204_n2376,
         DP_mult_204_n2375, DP_mult_204_n2374, DP_mult_204_n2373,
         DP_mult_204_n2372, DP_mult_204_n2371, DP_mult_204_n2370,
         DP_mult_204_n2369, DP_mult_204_n2368, DP_mult_204_n2367,
         DP_mult_204_n2366, DP_mult_204_n2365, DP_mult_204_n2364,
         DP_mult_204_n2363, DP_mult_204_n2362, DP_mult_204_n2361,
         DP_mult_204_n2360, DP_mult_204_n2359, DP_mult_204_n2358,
         DP_mult_204_n2357, DP_mult_204_n2356, DP_mult_204_n2355,
         DP_mult_204_n2354, DP_mult_204_n2353, DP_mult_204_n2352,
         DP_mult_204_n2351, DP_mult_204_n2350, DP_mult_204_n2349,
         DP_mult_204_n2348, DP_mult_204_n2347, DP_mult_204_n2346,
         DP_mult_204_n2345, DP_mult_204_n2344, DP_mult_204_n2343,
         DP_mult_204_n2342, DP_mult_204_n2341, DP_mult_204_n2340,
         DP_mult_204_n2339, DP_mult_204_n2338, DP_mult_204_n2337,
         DP_mult_204_n2336, DP_mult_204_n2335, DP_mult_204_n2334,
         DP_mult_204_n2333, DP_mult_204_n2332, DP_mult_204_n2331,
         DP_mult_204_n2330, DP_mult_204_n2329, DP_mult_204_n2328,
         DP_mult_204_n2327, DP_mult_204_n2326, DP_mult_204_n2325,
         DP_mult_204_n2324, DP_mult_204_n2323, DP_mult_204_n2322,
         DP_mult_204_n2321, DP_mult_204_n2320, DP_mult_204_n2319,
         DP_mult_204_n2318, DP_mult_204_n2317, DP_mult_204_n2316,
         DP_mult_204_n2315, DP_mult_204_n2314, DP_mult_204_n2313,
         DP_mult_204_n2312, DP_mult_204_n2311, DP_mult_204_n2310,
         DP_mult_204_n2309, DP_mult_204_n2308, DP_mult_204_n2307,
         DP_mult_204_n2306, DP_mult_204_n2305, DP_mult_204_n2304,
         DP_mult_204_n2303, DP_mult_204_n2302, DP_mult_204_n2301,
         DP_mult_204_n2300, DP_mult_204_n2299, DP_mult_204_n2298,
         DP_mult_204_n2297, DP_mult_204_n2296, DP_mult_204_n2295,
         DP_mult_204_n2294, DP_mult_204_n2293, DP_mult_204_n2292,
         DP_mult_204_n2291, DP_mult_204_n2290, DP_mult_204_n2289,
         DP_mult_204_n2288, DP_mult_204_n2287, DP_mult_204_n2286,
         DP_mult_204_n2285, DP_mult_204_n2284, DP_mult_204_n2283,
         DP_mult_204_n2282, DP_mult_204_n2281, DP_mult_204_n2280,
         DP_mult_204_n2279, DP_mult_204_n2278, DP_mult_204_n2277,
         DP_mult_204_n2276, DP_mult_204_n2275, DP_mult_204_n2274,
         DP_mult_204_n2273, DP_mult_204_n2272, DP_mult_204_n2271,
         DP_mult_204_n2270, DP_mult_204_n2269, DP_mult_204_n2268,
         DP_mult_204_n2267, DP_mult_204_n2266, DP_mult_204_n2265,
         DP_mult_204_n2264, DP_mult_204_n2263, DP_mult_204_n2262,
         DP_mult_204_n2261, DP_mult_204_n2260, DP_mult_204_n2259,
         DP_mult_204_n2258, DP_mult_204_n2257, DP_mult_204_n2256,
         DP_mult_204_n2255, DP_mult_204_n2254, DP_mult_204_n2253,
         DP_mult_204_n2252, DP_mult_204_n2251, DP_mult_204_n2250,
         DP_mult_204_n2249, DP_mult_204_n2248, DP_mult_204_n2247,
         DP_mult_204_n2246, DP_mult_204_n2245, DP_mult_204_n2244,
         DP_mult_204_n2243, DP_mult_204_n2242, DP_mult_204_n2241,
         DP_mult_204_n2240, DP_mult_204_n2239, DP_mult_204_n2238,
         DP_mult_204_n2237, DP_mult_204_n2236, DP_mult_204_n2235,
         DP_mult_204_n2234, DP_mult_204_n2233, DP_mult_204_n2232,
         DP_mult_204_n2231, DP_mult_204_n2230, DP_mult_204_n2229,
         DP_mult_204_n2228, DP_mult_204_n2227, DP_mult_204_n2226,
         DP_mult_204_n2225, DP_mult_204_n2224, DP_mult_204_n2223,
         DP_mult_204_n2222, DP_mult_204_n2221, DP_mult_204_n2220,
         DP_mult_204_n2219, DP_mult_204_n2218, DP_mult_204_n2217,
         DP_mult_204_n2216, DP_mult_204_n2215, DP_mult_204_n2214,
         DP_mult_204_n2213, DP_mult_204_n2212, DP_mult_204_n2211,
         DP_mult_204_n2210, DP_mult_204_n2209, DP_mult_204_n2208,
         DP_mult_204_n2207, DP_mult_204_n2206, DP_mult_204_n2205,
         DP_mult_204_n2204, DP_mult_204_n2203, DP_mult_204_n2202,
         DP_mult_204_n2201, DP_mult_204_n2200, DP_mult_204_n2199,
         DP_mult_204_n2198, DP_mult_204_n2197, DP_mult_204_n2196,
         DP_mult_204_n2195, DP_mult_204_n2194, DP_mult_204_n2193,
         DP_mult_204_n2192, DP_mult_204_n2191, DP_mult_204_n2190,
         DP_mult_204_n2189, DP_mult_204_n2188, DP_mult_204_n2187,
         DP_mult_204_n2186, DP_mult_204_n2185, DP_mult_204_n2184,
         DP_mult_204_n2183, DP_mult_204_n2182, DP_mult_204_n2181,
         DP_mult_204_n2180, DP_mult_204_n2179, DP_mult_204_n2178,
         DP_mult_204_n2177, DP_mult_204_n2176, DP_mult_204_n2175,
         DP_mult_204_n2174, DP_mult_204_n2173, DP_mult_204_n2172,
         DP_mult_204_n2171, DP_mult_204_n2170, DP_mult_204_n2169,
         DP_mult_204_n2168, DP_mult_204_n2167, DP_mult_204_n2166,
         DP_mult_204_n2165, DP_mult_204_n2164, DP_mult_204_n2163,
         DP_mult_204_n2162, DP_mult_204_n2161, DP_mult_204_n2160,
         DP_mult_204_n2159, DP_mult_204_n2158, DP_mult_204_n2157,
         DP_mult_204_n2156, DP_mult_204_n2155, DP_mult_204_n2154,
         DP_mult_204_n2153, DP_mult_204_n2152, DP_mult_204_n2151,
         DP_mult_204_n2150, DP_mult_204_n2149, DP_mult_204_n2148,
         DP_mult_204_n2147, DP_mult_204_n2146, DP_mult_204_n2145,
         DP_mult_204_n2144, DP_mult_204_n2143, DP_mult_204_n2142,
         DP_mult_204_n2141, DP_mult_204_n2140, DP_mult_204_n2139,
         DP_mult_204_n2138, DP_mult_204_n2137, DP_mult_204_n2136,
         DP_mult_204_n2135, DP_mult_204_n2134, DP_mult_204_n2133,
         DP_mult_204_n2132, DP_mult_204_n2131, DP_mult_204_n2130,
         DP_mult_204_n2129, DP_mult_204_n2128, DP_mult_204_n2127,
         DP_mult_204_n2126, DP_mult_204_n2125, DP_mult_204_n2124,
         DP_mult_204_n2123, DP_mult_204_n2122, DP_mult_204_n2121,
         DP_mult_204_n2120, DP_mult_204_n2119, DP_mult_204_n2118,
         DP_mult_204_n2117, DP_mult_204_n2116, DP_mult_204_n2115,
         DP_mult_204_n2114, DP_mult_204_n2113, DP_mult_204_n2112,
         DP_mult_204_n2111, DP_mult_204_n2110, DP_mult_204_n2109,
         DP_mult_204_n2108, DP_mult_204_n2107, DP_mult_204_n2106,
         DP_mult_204_n2105, DP_mult_204_n2104, DP_mult_204_n2103,
         DP_mult_204_n2102, DP_mult_204_n2101, DP_mult_204_n2100,
         DP_mult_204_n2099, DP_mult_204_n2098, DP_mult_204_n2097,
         DP_mult_204_n2096, DP_mult_204_n2095, DP_mult_204_n2094,
         DP_mult_204_n2093, DP_mult_204_n2092, DP_mult_204_n2091,
         DP_mult_204_n2090, DP_mult_204_n2089, DP_mult_204_n2088,
         DP_mult_204_n2087, DP_mult_204_n2086, DP_mult_204_n2085,
         DP_mult_204_n2084, DP_mult_204_n2083, DP_mult_204_n2082,
         DP_mult_204_n2081, DP_mult_204_n2080, DP_mult_204_n2079,
         DP_mult_204_n2078, DP_mult_204_n2077, DP_mult_204_n2076,
         DP_mult_204_n2075, DP_mult_204_n2074, DP_mult_204_n2073,
         DP_mult_204_n2072, DP_mult_204_n2071, DP_mult_204_n2070,
         DP_mult_204_n2069, DP_mult_204_n2068, DP_mult_204_n2067,
         DP_mult_204_n2066, DP_mult_204_n2065, DP_mult_204_n2064,
         DP_mult_204_n2063, DP_mult_204_n2062, DP_mult_204_n2061,
         DP_mult_204_n2060, DP_mult_204_n2059, DP_mult_204_n2058,
         DP_mult_204_n2057, DP_mult_204_n2056, DP_mult_204_n2055,
         DP_mult_204_n2054, DP_mult_204_n2053, DP_mult_204_n2052,
         DP_mult_204_n2051, DP_mult_204_n2050, DP_mult_204_n2049,
         DP_mult_204_n2048, DP_mult_204_n2047, DP_mult_204_n2046,
         DP_mult_204_n2045, DP_mult_204_n2044, DP_mult_204_n2043,
         DP_mult_204_n2042, DP_mult_204_n2041, DP_mult_204_n2040,
         DP_mult_204_n2039, DP_mult_204_n2038, DP_mult_204_n2037,
         DP_mult_204_n2036, DP_mult_204_n2035, DP_mult_204_n2034,
         DP_mult_204_n2033, DP_mult_204_n2032, DP_mult_204_n2031,
         DP_mult_204_n2030, DP_mult_204_n2029, DP_mult_204_n2028,
         DP_mult_204_n2027, DP_mult_204_n2026, DP_mult_204_n2025,
         DP_mult_204_n2024, DP_mult_204_n2023, DP_mult_204_n2022,
         DP_mult_204_n2021, DP_mult_204_n2020, DP_mult_204_n2019,
         DP_mult_204_n2018, DP_mult_204_n2017, DP_mult_204_n2016,
         DP_mult_204_n2015, DP_mult_204_n2014, DP_mult_204_n2013,
         DP_mult_204_n2012, DP_mult_204_n2011, DP_mult_204_n2010,
         DP_mult_204_n2009, DP_mult_204_n2008, DP_mult_204_n2007,
         DP_mult_204_n2006, DP_mult_204_n2005, DP_mult_204_n2004,
         DP_mult_204_n2003, DP_mult_204_n2002, DP_mult_204_n2001,
         DP_mult_204_n2000, DP_mult_204_n1999, DP_mult_204_n1998,
         DP_mult_204_n1997, DP_mult_204_n1996, DP_mult_204_n1995,
         DP_mult_204_n1994, DP_mult_204_n1993, DP_mult_204_n1992,
         DP_mult_204_n1991, DP_mult_204_n1990, DP_mult_204_n1989,
         DP_mult_204_n1988, DP_mult_204_n1987, DP_mult_204_n1986,
         DP_mult_204_n1985, DP_mult_204_n1984, DP_mult_204_n1983,
         DP_mult_204_n1982, DP_mult_204_n1981, DP_mult_204_n1980,
         DP_mult_204_n1979, DP_mult_204_n1978, DP_mult_204_n1977,
         DP_mult_204_n1976, DP_mult_204_n1975, DP_mult_204_n1974,
         DP_mult_204_n1973, DP_mult_204_n1972, DP_mult_204_n1971,
         DP_mult_204_n1970, DP_mult_204_n1969, DP_mult_204_n1968,
         DP_mult_204_n1967, DP_mult_204_n1966, DP_mult_204_n1965,
         DP_mult_204_n1964, DP_mult_204_n1963, DP_mult_204_n1962,
         DP_mult_204_n1961, DP_mult_204_n1960, DP_mult_204_n1959,
         DP_mult_204_n1958, DP_mult_204_n1957, DP_mult_204_n1956,
         DP_mult_204_n1955, DP_mult_204_n1954, DP_mult_204_n1953,
         DP_mult_204_n1952, DP_mult_204_n1951, DP_mult_204_n1950,
         DP_mult_204_n1949, DP_mult_204_n1948, DP_mult_204_n1947,
         DP_mult_204_n1946, DP_mult_204_n1945, DP_mult_204_n1944,
         DP_mult_204_n1943, DP_mult_204_n1942, DP_mult_204_n1941,
         DP_mult_204_n1940, DP_mult_204_n1939, DP_mult_204_n1938,
         DP_mult_204_n1937, DP_mult_204_n1936, DP_mult_204_n1935,
         DP_mult_204_n1934, DP_mult_204_n1933, DP_mult_204_n1932,
         DP_mult_204_n1931, DP_mult_204_n1930, DP_mult_204_n1929,
         DP_mult_204_n1817, DP_mult_204_n1816, DP_mult_204_n1815,
         DP_mult_204_n1814, DP_mult_204_n1813, DP_mult_204_n1812,
         DP_mult_204_n1811, DP_mult_204_n1810, DP_mult_204_n1809,
         DP_mult_204_n1808, DP_mult_204_n1807, DP_mult_204_n1806,
         DP_mult_204_n1781, DP_mult_204_n1780, DP_mult_204_n1779,
         DP_mult_204_n1778, DP_mult_204_n1777, DP_mult_204_n1776,
         DP_mult_204_n1775, DP_mult_204_n1774, DP_mult_204_n1773,
         DP_mult_204_n1772, DP_mult_204_n1771, DP_mult_204_n1770,
         DP_mult_204_n1769, DP_mult_204_n1768, DP_mult_204_n1767,
         DP_mult_204_n1766, DP_mult_204_n1765, DP_mult_204_n1764,
         DP_mult_204_n1763, DP_mult_204_n1762, DP_mult_204_n1761,
         DP_mult_204_n1760, DP_mult_204_n1759, DP_mult_204_n1758,
         DP_mult_204_n1757, DP_mult_204_n1756, DP_mult_204_n1755,
         DP_mult_204_n1754, DP_mult_204_n1753, DP_mult_204_n1752,
         DP_mult_204_n1751, DP_mult_204_n1750, DP_mult_204_n1749,
         DP_mult_204_n1748, DP_mult_204_n1747, DP_mult_204_n1746,
         DP_mult_204_n1745, DP_mult_204_n1744, DP_mult_204_n1743,
         DP_mult_204_n1742, DP_mult_204_n1741, DP_mult_204_n1740,
         DP_mult_204_n1739, DP_mult_204_n1738, DP_mult_204_n1737,
         DP_mult_204_n1736, DP_mult_204_n1735, DP_mult_204_n1734,
         DP_mult_204_n1733, DP_mult_204_n1732, DP_mult_204_n1731,
         DP_mult_204_n1730, DP_mult_204_n1729, DP_mult_204_n1728,
         DP_mult_204_n1727, DP_mult_204_n1726, DP_mult_204_n1725,
         DP_mult_204_n1724, DP_mult_204_n1723, DP_mult_204_n1722,
         DP_mult_204_n1721, DP_mult_204_n1720, DP_mult_204_n1719,
         DP_mult_204_n1718, DP_mult_204_n1717, DP_mult_204_n1716,
         DP_mult_204_n1715, DP_mult_204_n1714, DP_mult_204_n1713,
         DP_mult_204_n1712, DP_mult_204_n1711, DP_mult_204_n1710,
         DP_mult_204_n1709, DP_mult_204_n1708, DP_mult_204_n1707,
         DP_mult_204_n1706, DP_mult_204_n1705, DP_mult_204_n1704,
         DP_mult_204_n1703, DP_mult_204_n1702, DP_mult_204_n1701,
         DP_mult_204_n1700, DP_mult_204_n1699, DP_mult_204_n1698,
         DP_mult_204_n1697, DP_mult_204_n1696, DP_mult_204_n1695,
         DP_mult_204_n1694, DP_mult_204_n1693, DP_mult_204_n1692,
         DP_mult_204_n1691, DP_mult_204_n1690, DP_mult_204_n1689,
         DP_mult_204_n1688, DP_mult_204_n1687, DP_mult_204_n1686,
         DP_mult_204_n1685, DP_mult_204_n1684, DP_mult_204_n1683,
         DP_mult_204_n1682, DP_mult_204_n1681, DP_mult_204_n1680,
         DP_mult_204_n1679, DP_mult_204_n1678, DP_mult_204_n1677,
         DP_mult_204_n1676, DP_mult_204_n1675, DP_mult_204_n1674,
         DP_mult_204_n1673, DP_mult_204_n1672, DP_mult_204_n1671,
         DP_mult_204_n1670, DP_mult_204_n1669, DP_mult_204_n1668,
         DP_mult_204_n1667, DP_mult_204_n1666, DP_mult_204_n1665,
         DP_mult_204_n1664, DP_mult_204_n1663, DP_mult_204_n1662,
         DP_mult_204_n1661, DP_mult_204_n1660, DP_mult_204_n1659,
         DP_mult_204_n1658, DP_mult_204_n1657, DP_mult_204_n1656,
         DP_mult_204_n1655, DP_mult_204_n1654, DP_mult_204_n1653,
         DP_mult_204_n1652, DP_mult_204_n1651, DP_mult_204_n1650,
         DP_mult_204_n1649, DP_mult_204_n1648, DP_mult_204_n1647,
         DP_mult_204_n1646, DP_mult_204_n1645, DP_mult_204_n1644,
         DP_mult_204_n1643, DP_mult_204_n1642, DP_mult_204_n1641,
         DP_mult_204_n1640, DP_mult_204_n1639, DP_mult_204_n1638,
         DP_mult_204_n1637, DP_mult_204_n1636, DP_mult_204_n1635,
         DP_mult_204_n1634, DP_mult_204_n1633, DP_mult_204_n1632,
         DP_mult_204_n1631, DP_mult_204_n1630, DP_mult_204_n1629,
         DP_mult_204_n1628, DP_mult_204_n1627, DP_mult_204_n1626,
         DP_mult_204_n1625, DP_mult_204_n1624, DP_mult_204_n1623,
         DP_mult_204_n1622, DP_mult_204_n1621, DP_mult_204_n1620,
         DP_mult_204_n1619, DP_mult_204_n1618, DP_mult_204_n1617,
         DP_mult_204_n1616, DP_mult_204_n1615, DP_mult_204_n1614,
         DP_mult_204_n1613, DP_mult_204_n1612, DP_mult_204_n1611,
         DP_mult_204_n1610, DP_mult_204_n1609, DP_mult_204_n1608,
         DP_mult_204_n1607, DP_mult_204_n1606, DP_mult_204_n1605,
         DP_mult_204_n1604, DP_mult_204_n1603, DP_mult_204_n1602,
         DP_mult_204_n1601, DP_mult_204_n1600, DP_mult_204_n1599,
         DP_mult_204_n1598, DP_mult_204_n1597, DP_mult_204_n1596,
         DP_mult_204_n1595, DP_mult_204_n1594, DP_mult_204_n1593,
         DP_mult_204_n1592, DP_mult_204_n1591, DP_mult_204_n1590,
         DP_mult_204_n1589, DP_mult_204_n1588, DP_mult_204_n1587,
         DP_mult_204_n1586, DP_mult_204_n1585, DP_mult_204_n1584,
         DP_mult_204_n1583, DP_mult_204_n1582, DP_mult_204_n1581,
         DP_mult_204_n1580, DP_mult_204_n1579, DP_mult_204_n1578,
         DP_mult_204_n1577, DP_mult_204_n1576, DP_mult_204_n1575,
         DP_mult_204_n1574, DP_mult_204_n1573, DP_mult_204_n1572,
         DP_mult_204_n1571, DP_mult_204_n1570, DP_mult_204_n1569,
         DP_mult_204_n1568, DP_mult_204_n1567, DP_mult_204_n1566,
         DP_mult_204_n1565, DP_mult_204_n1564, DP_mult_204_n1563,
         DP_mult_204_n1562, DP_mult_204_n1561, DP_mult_204_n1560,
         DP_mult_204_n1559, DP_mult_204_n1558, DP_mult_204_n1557,
         DP_mult_204_n1556, DP_mult_204_n1555, DP_mult_204_n1554,
         DP_mult_204_n1553, DP_mult_204_n1552, DP_mult_204_n1551,
         DP_mult_204_n1550, DP_mult_204_n1549, DP_mult_204_n1548,
         DP_mult_204_n1547, DP_mult_204_n1546, DP_mult_204_n1545,
         DP_mult_204_n1544, DP_mult_204_n1543, DP_mult_204_n1542,
         DP_mult_204_n1541, DP_mult_204_n1540, DP_mult_204_n1539,
         DP_mult_204_n1538, DP_mult_204_n1537, DP_mult_204_n1536,
         DP_mult_204_n1535, DP_mult_204_n1534, DP_mult_204_n1533,
         DP_mult_204_n1532, DP_mult_204_n1531, DP_mult_204_n1530,
         DP_mult_204_n1529, DP_mult_204_n1528, DP_mult_204_n1527,
         DP_mult_204_n1526, DP_mult_204_n1525, DP_mult_204_n1524,
         DP_mult_204_n1523, DP_mult_204_n1522, DP_mult_204_n1521,
         DP_mult_204_n1520, DP_mult_204_n1519, DP_mult_204_n1518,
         DP_mult_204_n1517, DP_mult_204_n1516, DP_mult_204_n1515,
         DP_mult_204_n1514, DP_mult_204_n1513, DP_mult_204_n1512,
         DP_mult_204_n1511, DP_mult_204_n1510, DP_mult_204_n1509,
         DP_mult_204_n1508, DP_mult_204_n1507, DP_mult_204_n1506,
         DP_mult_204_n1505, DP_mult_204_n1504, DP_mult_204_n1503,
         DP_mult_204_n1502, DP_mult_204_n1501, DP_mult_204_n1500,
         DP_mult_204_n1499, DP_mult_204_n1498, DP_mult_204_n1497,
         DP_mult_204_n1496, DP_mult_204_n1495, DP_mult_204_n1494,
         DP_mult_204_n1493, DP_mult_204_n1492, DP_mult_204_n1491,
         DP_mult_204_n1490, DP_mult_204_n1489, DP_mult_204_n1488,
         DP_mult_204_n1487, DP_mult_204_n1486, DP_mult_204_n1485,
         DP_mult_204_n1484, DP_mult_204_n1483, DP_mult_204_n1482,
         DP_mult_204_n1481, DP_mult_204_n1480, DP_mult_204_n1479,
         DP_mult_204_n1478, DP_mult_204_n1477, DP_mult_204_n1476,
         DP_mult_204_n1475, DP_mult_204_n1474, DP_mult_204_n1473,
         DP_mult_204_n1472, DP_mult_204_n1471, DP_mult_204_n1470,
         DP_mult_204_n1469, DP_mult_204_n1468, DP_mult_204_n1467,
         DP_mult_204_n1466, DP_mult_204_n1465, DP_mult_204_n1464,
         DP_mult_204_n1463, DP_mult_204_n1462, DP_mult_204_n1461,
         DP_mult_204_n1460, DP_mult_204_n1459, DP_mult_204_n1458,
         DP_mult_204_n1457, DP_mult_204_n1456, DP_mult_204_n1455,
         DP_mult_204_n1454, DP_mult_204_n1453, DP_mult_204_n1452,
         DP_mult_204_n1451, DP_mult_204_n1450, DP_mult_204_n1449,
         DP_mult_204_n1448, DP_mult_204_n1447, DP_mult_204_n1446,
         DP_mult_204_n1445, DP_mult_204_n1444, DP_mult_204_n1443,
         DP_mult_204_n1442, DP_mult_204_n1441, DP_mult_204_n1440,
         DP_mult_204_n1439, DP_mult_204_n1438, DP_mult_204_n1437,
         DP_mult_204_n1436, DP_mult_204_n1435, DP_mult_204_n1434,
         DP_mult_204_n1433, DP_mult_204_n1432, DP_mult_204_n1431,
         DP_mult_204_n1430, DP_mult_204_n1429, DP_mult_204_n1428,
         DP_mult_204_n1427, DP_mult_204_n1426, DP_mult_204_n1425,
         DP_mult_204_n1424, DP_mult_204_n1423, DP_mult_204_n1422,
         DP_mult_204_n1421, DP_mult_204_n1420, DP_mult_204_n1419,
         DP_mult_204_n1418, DP_mult_204_n1417, DP_mult_204_n1416,
         DP_mult_204_n1415, DP_mult_204_n1414, DP_mult_204_n1413,
         DP_mult_204_n1412, DP_mult_204_n1411, DP_mult_204_n1410,
         DP_mult_204_n1409, DP_mult_204_n1408, DP_mult_204_n1407,
         DP_mult_204_n1406, DP_mult_204_n1405, DP_mult_204_n1404,
         DP_mult_204_n1403, DP_mult_204_n1402, DP_mult_204_n1401,
         DP_mult_204_n1400, DP_mult_204_n1399, DP_mult_204_n1398,
         DP_mult_204_n1397, DP_mult_204_n1396, DP_mult_204_n1395,
         DP_mult_204_n1394, DP_mult_204_n1393, DP_mult_204_n1392,
         DP_mult_204_n1391, DP_mult_204_n1390, DP_mult_204_n1389,
         DP_mult_204_n1388, DP_mult_204_n1387, DP_mult_204_n1386,
         DP_mult_204_n1385, DP_mult_204_n1384, DP_mult_204_n1383,
         DP_mult_204_n1382, DP_mult_204_n1381, DP_mult_204_n1380,
         DP_mult_204_n1379, DP_mult_204_n1378, DP_mult_204_n1377,
         DP_mult_204_n1376, DP_mult_204_n1375, DP_mult_204_n1374,
         DP_mult_204_n1373, DP_mult_204_n1372, DP_mult_204_n1371,
         DP_mult_204_n1370, DP_mult_204_n1369, DP_mult_204_n1368,
         DP_mult_204_n1367, DP_mult_204_n1366, DP_mult_204_n1365,
         DP_mult_204_n1364, DP_mult_204_n1363, DP_mult_204_n1362,
         DP_mult_204_n1361, DP_mult_204_n1360, DP_mult_204_n1359,
         DP_mult_204_n1358, DP_mult_204_n1357, DP_mult_204_n1356,
         DP_mult_204_n1355, DP_mult_204_n1354, DP_mult_204_n1353,
         DP_mult_204_n1352, DP_mult_204_n1351, DP_mult_204_n1350,
         DP_mult_204_n1349, DP_mult_204_n1348, DP_mult_204_n1347,
         DP_mult_204_n1346, DP_mult_204_n1345, DP_mult_204_n1344,
         DP_mult_204_n1343, DP_mult_204_n1342, DP_mult_204_n1341,
         DP_mult_204_n1340, DP_mult_204_n1339, DP_mult_204_n1338,
         DP_mult_204_n1337, DP_mult_204_n1336, DP_mult_204_n1335,
         DP_mult_204_n1334, DP_mult_204_n1333, DP_mult_204_n1332,
         DP_mult_204_n1331, DP_mult_204_n1330, DP_mult_204_n1329,
         DP_mult_204_n1328, DP_mult_204_n1327, DP_mult_204_n1326,
         DP_mult_204_n1325, DP_mult_204_n1324, DP_mult_204_n1323,
         DP_mult_204_n1322, DP_mult_204_n1321, DP_mult_204_n1320,
         DP_mult_204_n1319, DP_mult_204_n1318, DP_mult_204_n1317,
         DP_mult_204_n1316, DP_mult_204_n1315, DP_mult_204_n1314,
         DP_mult_204_n1313, DP_mult_204_n1312, DP_mult_204_n1311,
         DP_mult_204_n1310, DP_mult_204_n1309, DP_mult_204_n1308,
         DP_mult_204_n1307, DP_mult_204_n1306, DP_mult_204_n1305,
         DP_mult_204_n1304, DP_mult_204_n1303, DP_mult_204_n1302,
         DP_mult_204_n1301, DP_mult_204_n1300, DP_mult_204_n1299,
         DP_mult_204_n1298, DP_mult_204_n1297, DP_mult_204_n1296,
         DP_mult_204_n1295, DP_mult_204_n1294, DP_mult_204_n1293,
         DP_mult_204_n1292, DP_mult_204_n1291, DP_mult_204_n1290,
         DP_mult_204_n1289, DP_mult_204_n1288, DP_mult_204_n1287,
         DP_mult_204_n1286, DP_mult_204_n1285, DP_mult_204_n1284,
         DP_mult_204_n1283, DP_mult_204_n1282, DP_mult_204_n1281,
         DP_mult_204_n1280, DP_mult_204_n1279, DP_mult_204_n1278,
         DP_mult_204_n1277, DP_mult_204_n1276, DP_mult_204_n1275,
         DP_mult_204_n1274, DP_mult_204_n1273, DP_mult_204_n1272,
         DP_mult_204_n1271, DP_mult_204_n1270, DP_mult_204_n1269,
         DP_mult_204_n1268, DP_mult_204_n1267, DP_mult_204_n1266,
         DP_mult_204_n1265, DP_mult_204_n1264, DP_mult_204_n1263,
         DP_mult_204_n1261, DP_mult_204_n1260, DP_mult_204_n1259,
         DP_mult_204_n1258, DP_mult_204_n1257, DP_mult_204_n1256,
         DP_mult_204_n1255, DP_mult_204_n1254, DP_mult_204_n1253,
         DP_mult_204_n1252, DP_mult_204_n1251, DP_mult_204_n1250,
         DP_mult_204_n1249, DP_mult_204_n1248, DP_mult_204_n1247,
         DP_mult_204_n1246, DP_mult_204_n1245, DP_mult_204_n1244,
         DP_mult_204_n1243, DP_mult_204_n1242, DP_mult_204_n1241,
         DP_mult_204_n1240, DP_mult_204_n1239, DP_mult_204_n1238,
         DP_mult_204_n1237, DP_mult_204_n1236, DP_mult_204_n1235,
         DP_mult_204_n1234, DP_mult_204_n1233, DP_mult_204_n1232,
         DP_mult_204_n1231, DP_mult_204_n1230, DP_mult_204_n1229,
         DP_mult_204_n1228, DP_mult_204_n1227, DP_mult_204_n1226,
         DP_mult_204_n1225, DP_mult_204_n1224, DP_mult_204_n1223,
         DP_mult_204_n1222, DP_mult_204_n1221, DP_mult_204_n1220,
         DP_mult_204_n1219, DP_mult_204_n1218, DP_mult_204_n1217,
         DP_mult_204_n1216, DP_mult_204_n1215, DP_mult_204_n1214,
         DP_mult_204_n1213, DP_mult_204_n1212, DP_mult_204_n1211,
         DP_mult_204_n1210, DP_mult_204_n1209, DP_mult_204_n1208,
         DP_mult_204_n1207, DP_mult_204_n1206, DP_mult_204_n1205,
         DP_mult_204_n1204, DP_mult_204_n1203, DP_mult_204_n1202,
         DP_mult_204_n1201, DP_mult_204_n1200, DP_mult_204_n1199,
         DP_mult_204_n1198, DP_mult_204_n1197, DP_mult_204_n1196,
         DP_mult_204_n1195, DP_mult_204_n1194, DP_mult_204_n1193,
         DP_mult_204_n1192, DP_mult_204_n1191, DP_mult_204_n1190,
         DP_mult_204_n1189, DP_mult_204_n1188, DP_mult_204_n1187,
         DP_mult_204_n1186, DP_mult_204_n1185, DP_mult_204_n1184,
         DP_mult_204_n1183, DP_mult_204_n1182, DP_mult_204_n1181,
         DP_mult_204_n1180, DP_mult_204_n1179, DP_mult_204_n1178,
         DP_mult_204_n1177, DP_mult_204_n1176, DP_mult_204_n1175,
         DP_mult_204_n1174, DP_mult_204_n1173, DP_mult_204_n1172,
         DP_mult_204_n1171, DP_mult_204_n1170, DP_mult_204_n1169,
         DP_mult_204_n1168, DP_mult_204_n1167, DP_mult_204_n1166,
         DP_mult_204_n1165, DP_mult_204_n1164, DP_mult_204_n1163,
         DP_mult_204_n1162, DP_mult_204_n1161, DP_mult_204_n1160,
         DP_mult_204_n1159, DP_mult_204_n1158, DP_mult_204_n1157,
         DP_mult_204_n1156, DP_mult_204_n1155, DP_mult_204_n1154,
         DP_mult_204_n1153, DP_mult_204_n1152, DP_mult_204_n1151,
         DP_mult_204_n1150, DP_mult_204_n1149, DP_mult_204_n1148,
         DP_mult_204_n1147, DP_mult_204_n1146, DP_mult_204_n1145,
         DP_mult_204_n1144, DP_mult_204_n1143, DP_mult_204_n1142,
         DP_mult_204_n1141, DP_mult_204_n1140, DP_mult_204_n1139,
         DP_mult_204_n1138, DP_mult_204_n1137, DP_mult_204_n1136,
         DP_mult_204_n1135, DP_mult_204_n1134, DP_mult_204_n1133,
         DP_mult_204_n1132, DP_mult_204_n1131, DP_mult_204_n1130,
         DP_mult_204_n1129, DP_mult_204_n1128, DP_mult_204_n1127,
         DP_mult_204_n1126, DP_mult_204_n1125, DP_mult_204_n1124,
         DP_mult_204_n1123, DP_mult_204_n1122, DP_mult_204_n1121,
         DP_mult_204_n1120, DP_mult_204_n1119, DP_mult_204_n1118,
         DP_mult_204_n1117, DP_mult_204_n1116, DP_mult_204_n1115,
         DP_mult_204_n1114, DP_mult_204_n1113, DP_mult_204_n1112,
         DP_mult_204_n1111, DP_mult_204_n1110, DP_mult_204_n1109,
         DP_mult_204_n1108, DP_mult_204_n1107, DP_mult_204_n1106,
         DP_mult_204_n1105, DP_mult_204_n1104, DP_mult_204_n1103,
         DP_mult_204_n1102, DP_mult_204_n1101, DP_mult_204_n1100,
         DP_mult_204_n1099, DP_mult_204_n1098, DP_mult_204_n1097,
         DP_mult_204_n1096, DP_mult_204_n1095, DP_mult_204_n1094,
         DP_mult_204_n1093, DP_mult_204_n1092, DP_mult_204_n1091,
         DP_mult_204_n1090, DP_mult_204_n1089, DP_mult_204_n1088,
         DP_mult_204_n1087, DP_mult_204_n1086, DP_mult_204_n1085,
         DP_mult_204_n1084, DP_mult_204_n1083, DP_mult_204_n1082,
         DP_mult_204_n1081, DP_mult_204_n1080, DP_mult_204_n1079,
         DP_mult_204_n1078, DP_mult_204_n1077, DP_mult_204_n1076,
         DP_mult_204_n1075, DP_mult_204_n1074, DP_mult_204_n1073,
         DP_mult_204_n1072, DP_mult_204_n1071, DP_mult_204_n1070,
         DP_mult_204_n1069, DP_mult_204_n1068, DP_mult_204_n1067,
         DP_mult_204_n1066, DP_mult_204_n1065, DP_mult_204_n1064,
         DP_mult_204_n1063, DP_mult_204_n1062, DP_mult_204_n1061,
         DP_mult_204_n1060, DP_mult_204_n1059, DP_mult_204_n1058,
         DP_mult_204_n1057, DP_mult_204_n1056, DP_mult_204_n1055,
         DP_mult_204_n1054, DP_mult_204_n1053, DP_mult_204_n1052,
         DP_mult_204_n1051, DP_mult_204_n1050, DP_mult_204_n1049,
         DP_mult_204_n1048, DP_mult_204_n1047, DP_mult_204_n1046,
         DP_mult_204_n1045, DP_mult_204_n1044, DP_mult_204_n1043,
         DP_mult_204_n1042, DP_mult_204_n1041, DP_mult_204_n1040,
         DP_mult_204_n1039, DP_mult_204_n1038, DP_mult_204_n1037,
         DP_mult_204_n1036, DP_mult_204_n1035, DP_mult_204_n1034,
         DP_mult_204_n1033, DP_mult_204_n1032, DP_mult_204_n1031,
         DP_mult_204_n1030, DP_mult_204_n1029, DP_mult_204_n1028,
         DP_mult_204_n1027, DP_mult_204_n1026, DP_mult_204_n1025,
         DP_mult_204_n1024, DP_mult_204_n1023, DP_mult_204_n1022,
         DP_mult_204_n1021, DP_mult_204_n1020, DP_mult_204_n1019,
         DP_mult_204_n1018, DP_mult_204_n1017, DP_mult_204_n1016,
         DP_mult_204_n1015, DP_mult_204_n1014, DP_mult_204_n1013,
         DP_mult_204_n1012, DP_mult_204_n1011, DP_mult_204_n1010,
         DP_mult_204_n1009, DP_mult_204_n1008, DP_mult_204_n1007,
         DP_mult_204_n1006, DP_mult_204_n1005, DP_mult_204_n1004,
         DP_mult_204_n1003, DP_mult_204_n1002, DP_mult_204_n1001,
         DP_mult_204_n999, DP_mult_204_n998, DP_mult_204_n997,
         DP_mult_204_n996, DP_mult_204_n995, DP_mult_204_n994,
         DP_mult_204_n993, DP_mult_204_n992, DP_mult_204_n991,
         DP_mult_204_n990, DP_mult_204_n989, DP_mult_204_n988,
         DP_mult_204_n987, DP_mult_204_n986, DP_mult_204_n985,
         DP_mult_204_n984, DP_mult_204_n983, DP_mult_204_n982,
         DP_mult_204_n981, DP_mult_204_n980, DP_mult_204_n979,
         DP_mult_204_n978, DP_mult_204_n977, DP_mult_204_n976,
         DP_mult_204_n975, DP_mult_204_n974, DP_mult_204_n973,
         DP_mult_204_n972, DP_mult_204_n971, DP_mult_204_n970,
         DP_mult_204_n969, DP_mult_204_n968, DP_mult_204_n967,
         DP_mult_204_n966, DP_mult_204_n965, DP_mult_204_n964,
         DP_mult_204_n963, DP_mult_204_n962, DP_mult_204_n961,
         DP_mult_204_n959, DP_mult_204_n958, DP_mult_204_n957,
         DP_mult_204_n956, DP_mult_204_n955, DP_mult_204_n954,
         DP_mult_204_n953, DP_mult_204_n952, DP_mult_204_n951,
         DP_mult_204_n950, DP_mult_204_n949, DP_mult_204_n948,
         DP_mult_204_n947, DP_mult_204_n946, DP_mult_204_n945,
         DP_mult_204_n944, DP_mult_204_n943, DP_mult_204_n942,
         DP_mult_204_n941, DP_mult_204_n940, DP_mult_204_n939,
         DP_mult_204_n938, DP_mult_204_n937, DP_mult_204_n936,
         DP_mult_204_n935, DP_mult_204_n934, DP_mult_204_n933,
         DP_mult_204_n932, DP_mult_204_n931, DP_mult_204_n930,
         DP_mult_204_n929, DP_mult_204_n928, DP_mult_204_n927,
         DP_mult_204_n926, DP_mult_204_n925, DP_mult_204_n924,
         DP_mult_204_n923, DP_mult_204_n922, DP_mult_204_n921,
         DP_mult_204_n920, DP_mult_204_n919, DP_mult_204_n918,
         DP_mult_204_n917, DP_mult_204_n916, DP_mult_204_n915,
         DP_mult_204_n914, DP_mult_204_n913, DP_mult_204_n912,
         DP_mult_204_n911, DP_mult_204_n910, DP_mult_204_n909,
         DP_mult_204_n908, DP_mult_204_n907, DP_mult_204_n906,
         DP_mult_204_n905, DP_mult_204_n904, DP_mult_204_n903,
         DP_mult_204_n902, DP_mult_204_n901, DP_mult_204_n900,
         DP_mult_204_n899, DP_mult_204_n898, DP_mult_204_n897,
         DP_mult_204_n896, DP_mult_204_n895, DP_mult_204_n894,
         DP_mult_204_n893, DP_mult_204_n892, DP_mult_204_n891,
         DP_mult_204_n890, DP_mult_204_n889, DP_mult_204_n888,
         DP_mult_204_n887, DP_mult_204_n886, DP_mult_204_n885,
         DP_mult_204_n884, DP_mult_204_n883, DP_mult_204_n882,
         DP_mult_204_n881, DP_mult_204_n880, DP_mult_204_n879,
         DP_mult_204_n878, DP_mult_204_n877, DP_mult_204_n876,
         DP_mult_204_n875, DP_mult_204_n874, DP_mult_204_n873,
         DP_mult_204_n872, DP_mult_204_n871, DP_mult_204_n870,
         DP_mult_204_n869, DP_mult_204_n868, DP_mult_204_n867,
         DP_mult_204_n866, DP_mult_204_n865, DP_mult_204_n864,
         DP_mult_204_n863, DP_mult_204_n862, DP_mult_204_n861,
         DP_mult_204_n860, DP_mult_204_n859, DP_mult_204_n858,
         DP_mult_204_n857, DP_mult_204_n856, DP_mult_204_n855,
         DP_mult_204_n854, DP_mult_204_n853, DP_mult_204_n852,
         DP_mult_204_n851, DP_mult_204_n850, DP_mult_204_n849,
         DP_mult_204_n848, DP_mult_204_n847, DP_mult_204_n846,
         DP_mult_204_n845, DP_mult_204_n844, DP_mult_204_n843,
         DP_mult_204_n842, DP_mult_204_n841, DP_mult_204_n840,
         DP_mult_204_n839, DP_mult_204_n838, DP_mult_204_n837,
         DP_mult_204_n836, DP_mult_204_n835, DP_mult_204_n834,
         DP_mult_204_n833, DP_mult_204_n832, DP_mult_204_n831,
         DP_mult_204_n830, DP_mult_204_n829, DP_mult_204_n828,
         DP_mult_204_n827, DP_mult_204_n826, DP_mult_204_n825,
         DP_mult_204_n824, DP_mult_204_n823, DP_mult_204_n822,
         DP_mult_204_n821, DP_mult_204_n820, DP_mult_204_n819,
         DP_mult_204_n818, DP_mult_204_n817, DP_mult_204_n816,
         DP_mult_204_n815, DP_mult_204_n814, DP_mult_204_n813,
         DP_mult_204_n812, DP_mult_204_n811, DP_mult_204_n810,
         DP_mult_204_n809, DP_mult_204_n808, DP_mult_204_n807,
         DP_mult_204_n806, DP_mult_204_n805, DP_mult_204_n804,
         DP_mult_204_n803, DP_mult_204_n802, DP_mult_204_n801,
         DP_mult_204_n800, DP_mult_204_n799, DP_mult_204_n798,
         DP_mult_204_n797, DP_mult_204_n796, DP_mult_204_n795,
         DP_mult_204_n794, DP_mult_204_n793, DP_mult_204_n792,
         DP_mult_204_n791, DP_mult_204_n790, DP_mult_204_n789,
         DP_mult_204_n788, DP_mult_204_n787, DP_mult_204_n786,
         DP_mult_204_n785, DP_mult_204_n784, DP_mult_204_n783,
         DP_mult_204_n782, DP_mult_204_n781, DP_mult_204_n780,
         DP_mult_204_n779, DP_mult_204_n778, DP_mult_204_n777,
         DP_mult_204_n776, DP_mult_204_n775, DP_mult_204_n774,
         DP_mult_204_n773, DP_mult_204_n772, DP_mult_204_n771,
         DP_mult_204_n770, DP_mult_204_n769, DP_mult_204_n768,
         DP_mult_204_n767, DP_mult_204_n766, DP_mult_204_n765,
         DP_mult_204_n764, DP_mult_204_n763, DP_mult_204_n762,
         DP_mult_204_n761, DP_mult_204_n760, DP_mult_204_n759,
         DP_mult_204_n758, DP_mult_204_n757, DP_mult_204_n756,
         DP_mult_204_n755, DP_mult_204_n754, DP_mult_204_n753,
         DP_mult_204_n752, DP_mult_204_n751, DP_mult_204_n750,
         DP_mult_204_n749, DP_mult_204_n748, DP_mult_204_n747,
         DP_mult_204_n746, DP_mult_204_n745, DP_mult_204_n744,
         DP_mult_204_n743, DP_mult_204_n742, DP_mult_204_n741,
         DP_mult_204_n740, DP_mult_204_n739, DP_mult_204_n738,
         DP_mult_204_n737, DP_mult_204_n736, DP_mult_204_n735,
         DP_mult_204_n734, DP_mult_204_n733, DP_mult_204_n732,
         DP_mult_204_n731, DP_mult_204_n730, DP_mult_204_n729,
         DP_mult_204_n728, DP_mult_204_n727, DP_mult_204_n726,
         DP_mult_204_n725, DP_mult_204_n724, DP_mult_204_n723,
         DP_mult_204_n722, DP_mult_204_n721, DP_mult_204_n720,
         DP_mult_204_n719, DP_mult_204_n718, DP_mult_204_n717,
         DP_mult_204_n716, DP_mult_204_n715, DP_mult_204_n714,
         DP_mult_204_n713, DP_mult_204_n712, DP_mult_204_n711,
         DP_mult_204_n710, DP_mult_204_n709, DP_mult_204_n708,
         DP_mult_204_n707, DP_mult_204_n706, DP_mult_204_n705,
         DP_mult_204_n704, DP_mult_204_n703, DP_mult_204_n702,
         DP_mult_204_n701, DP_mult_204_n700, DP_mult_204_n699,
         DP_mult_204_n698, DP_mult_204_n697, DP_mult_204_n696,
         DP_mult_204_n695, DP_mult_204_n694, DP_mult_204_n693,
         DP_mult_204_n692, DP_mult_204_n691, DP_mult_204_n690,
         DP_mult_204_n689, DP_mult_204_n688, DP_mult_204_n687,
         DP_mult_204_n686, DP_mult_204_n685, DP_mult_204_n684,
         DP_mult_204_n683, DP_mult_204_n682, DP_mult_204_n681,
         DP_mult_204_n680, DP_mult_204_n679, DP_mult_204_n678,
         DP_mult_204_n677, DP_mult_204_n676, DP_mult_204_n672,
         DP_mult_204_n670, DP_mult_204_n668, DP_mult_204_n663,
         DP_mult_204_n662, DP_mult_204_n661, DP_mult_204_n657,
         DP_mult_204_n646, DP_mult_204_n645, DP_mult_204_n644,
         DP_mult_204_n643, DP_mult_204_n638, DP_mult_204_n637,
         DP_mult_204_n636, DP_mult_204_n635, DP_mult_204_n634,
         DP_mult_204_n633, DP_mult_204_n632, DP_mult_204_n631,
         DP_mult_204_n630, DP_mult_204_n629, DP_mult_204_n628,
         DP_mult_204_n627, DP_mult_204_n626, DP_mult_204_n625,
         DP_mult_204_n620, DP_mult_204_n611, DP_mult_204_n610,
         DP_mult_204_n609, DP_mult_204_n600, DP_mult_204_n599,
         DP_mult_204_n598, DP_mult_204_n597, DP_mult_204_n596,
         DP_mult_204_n595, DP_mult_204_n594, DP_mult_204_n593,
         DP_mult_204_n592, DP_mult_204_n591, DP_mult_204_n590,
         DP_mult_204_n589, DP_mult_204_n588, DP_mult_204_n583,
         DP_mult_204_n582, DP_mult_204_n581, DP_mult_204_n572,
         DP_mult_204_n570, DP_mult_204_n568, DP_mult_204_n567,
         DP_mult_204_n566, DP_mult_204_n565, DP_mult_204_n564,
         DP_mult_204_n563, DP_mult_204_n562, DP_mult_204_n561,
         DP_mult_204_n560, DP_mult_204_n559, DP_mult_204_n558,
         DP_mult_204_n555, DP_mult_204_n554, DP_mult_204_n553,
         DP_mult_204_n552, DP_mult_204_n551, DP_mult_204_n550,
         DP_mult_204_n547, DP_mult_204_n546, DP_mult_204_n545,
         DP_mult_204_n544, DP_mult_204_n543, DP_mult_204_n542,
         DP_mult_204_n541, DP_mult_204_n540, DP_mult_204_n539,
         DP_mult_204_n538, DP_mult_204_n536, DP_mult_204_n535,
         DP_mult_204_n534, DP_mult_204_n533, DP_mult_204_n532,
         DP_mult_204_n531, DP_mult_204_n526, DP_mult_204_n525,
         DP_mult_204_n524, DP_mult_204_n522, DP_mult_204_n521,
         DP_mult_204_n520, DP_mult_204_n519, DP_mult_204_n517,
         DP_mult_204_n516, DP_mult_204_n515, DP_mult_204_n514,
         DP_mult_204_n513, DP_mult_204_n512, DP_mult_204_n511,
         DP_mult_204_n508, DP_mult_204_n507, DP_mult_204_n506,
         DP_mult_204_n505, DP_mult_204_n504, DP_mult_204_n503,
         DP_mult_204_n502, DP_mult_204_n499, DP_mult_204_n498,
         DP_mult_204_n497, DP_mult_204_n496, DP_mult_204_n495,
         DP_mult_204_n492, DP_mult_204_n490, DP_mult_204_n489,
         DP_mult_204_n488, DP_mult_204_n487, DP_mult_204_n486,
         DP_mult_204_n483, DP_mult_204_n481, DP_mult_204_n480,
         DP_mult_204_n479, DP_mult_204_n478, DP_mult_204_n477,
         DP_mult_204_n476, DP_mult_204_n475, DP_mult_204_n474,
         DP_mult_204_n472, DP_mult_204_n468, DP_mult_204_n467,
         DP_mult_204_n466, DP_mult_204_n465, DP_mult_204_n464,
         DP_mult_204_n463, DP_mult_204_n462, DP_mult_204_n461,
         DP_mult_204_n459, DP_mult_204_n457, DP_mult_204_n456,
         DP_mult_204_n455, DP_mult_204_n454, DP_mult_204_n453,
         DP_mult_204_n452, DP_mult_204_n451, DP_mult_204_n450,
         DP_mult_204_n445, DP_mult_204_n439, DP_mult_204_n438,
         DP_mult_204_n437, DP_mult_204_n436, DP_mult_204_n435,
         DP_mult_204_n434, DP_mult_204_n432, DP_mult_204_n431,
         DP_mult_204_n430, DP_mult_204_n429, DP_mult_204_n428,
         DP_mult_204_n427, DP_mult_204_n426, DP_mult_204_n423,
         DP_mult_204_n422, DP_mult_204_n421, DP_mult_204_n420,
         DP_mult_204_n419, DP_mult_204_n418, DP_mult_204_n416,
         DP_mult_204_n412, DP_mult_204_n411, DP_mult_204_n410,
         DP_mult_204_n409, DP_mult_204_n407, DP_mult_204_n405,
         DP_mult_204_n402, DP_mult_204_n401, DP_mult_204_n400,
         DP_mult_204_n399, DP_mult_204_n398, DP_mult_204_n397,
         DP_mult_204_n396, DP_mult_204_n394, DP_mult_204_n390,
         DP_mult_204_n389, DP_mult_204_n388, DP_mult_204_n387,
         DP_mult_204_n384, DP_mult_204_n383, DP_mult_204_n382,
         DP_mult_204_n381, DP_mult_204_n380, DP_mult_204_n379,
         DP_mult_204_n378, DP_mult_204_n376, DP_mult_204_n372,
         DP_mult_204_n371, DP_mult_204_n370, DP_mult_204_n369,
         DP_mult_204_n367, DP_mult_204_n365, DP_mult_204_n364,
         DP_mult_204_n363, DP_mult_204_n362, DP_mult_204_n361,
         DP_mult_204_n360, DP_mult_204_n359, DP_mult_204_n356,
         DP_mult_204_n355, DP_mult_204_n354, DP_mult_204_n353,
         DP_mult_204_n352, DP_mult_204_n350, DP_mult_204_n348,
         DP_mult_204_n347, DP_mult_204_n346, DP_mult_204_n345,
         DP_mult_204_n344, DP_mult_204_n343, DP_mult_204_n342,
         DP_mult_204_n341, DP_mult_204_n339, DP_mult_204_n337,
         DP_mult_204_n336, DP_mult_204_n335, DP_mult_204_n334,
         DP_mult_204_n333, DP_mult_204_n332, DP_mult_204_n327,
         DP_mult_204_n326, DP_mult_204_n325, DP_mult_204_n322,
         DP_mult_204_n320, DP_mult_204_n319, DP_mult_204_n318,
         DP_mult_204_n317, DP_mult_204_n316, DP_mult_204_n315,
         DP_mult_204_n314, DP_mult_204_n313, DP_mult_204_n311,
         DP_mult_204_n310, DP_mult_204_n309, DP_mult_204_n308,
         DP_mult_204_n307, DP_mult_204_n306, DP_mult_204_n305,
         DP_mult_204_n304, DP_mult_204_n303, DP_mult_204_n302,
         DP_mult_204_n301, DP_mult_204_n297, DP_mult_204_n295,
         DP_mult_204_n293, DP_mult_204_n287, DP_mult_204_n285,
         DP_mult_204_n251, DP_mult_206_n2339, DP_mult_206_n2338,
         DP_mult_206_n2337, DP_mult_206_n2336, DP_mult_206_n2335,
         DP_mult_206_n2334, DP_mult_206_n2333, DP_mult_206_n2332,
         DP_mult_206_n2331, DP_mult_206_n2330, DP_mult_206_n2329,
         DP_mult_206_n2328, DP_mult_206_n2327, DP_mult_206_n2326,
         DP_mult_206_n2325, DP_mult_206_n2324, DP_mult_206_n2323,
         DP_mult_206_n2322, DP_mult_206_n2321, DP_mult_206_n2320,
         DP_mult_206_n2319, DP_mult_206_n2318, DP_mult_206_n2317,
         DP_mult_206_n2316, DP_mult_206_n2315, DP_mult_206_n2314,
         DP_mult_206_n2313, DP_mult_206_n2312, DP_mult_206_n2311,
         DP_mult_206_n2310, DP_mult_206_n2309, DP_mult_206_n2308,
         DP_mult_206_n2307, DP_mult_206_n2306, DP_mult_206_n2305,
         DP_mult_206_n2304, DP_mult_206_n2303, DP_mult_206_n2302,
         DP_mult_206_n2301, DP_mult_206_n2300, DP_mult_206_n2299,
         DP_mult_206_n2298, DP_mult_206_n2297, DP_mult_206_n2296,
         DP_mult_206_n2295, DP_mult_206_n2294, DP_mult_206_n2293,
         DP_mult_206_n2292, DP_mult_206_n2291, DP_mult_206_n2290,
         DP_mult_206_n2289, DP_mult_206_n2288, DP_mult_206_n2287,
         DP_mult_206_n2286, DP_mult_206_n2285, DP_mult_206_n2284,
         DP_mult_206_n2283, DP_mult_206_n2282, DP_mult_206_n2281,
         DP_mult_206_n2280, DP_mult_206_n2279, DP_mult_206_n2278,
         DP_mult_206_n2277, DP_mult_206_n2276, DP_mult_206_n2275,
         DP_mult_206_n2274, DP_mult_206_n2273, DP_mult_206_n2272,
         DP_mult_206_n2271, DP_mult_206_n2270, DP_mult_206_n2269,
         DP_mult_206_n2268, DP_mult_206_n2267, DP_mult_206_n2266,
         DP_mult_206_n2265, DP_mult_206_n2264, DP_mult_206_n2263,
         DP_mult_206_n2262, DP_mult_206_n2261, DP_mult_206_n2260,
         DP_mult_206_n2259, DP_mult_206_n2258, DP_mult_206_n2257,
         DP_mult_206_n2256, DP_mult_206_n2255, DP_mult_206_n2254,
         DP_mult_206_n2253, DP_mult_206_n2252, DP_mult_206_n2251,
         DP_mult_206_n2250, DP_mult_206_n2249, DP_mult_206_n2248,
         DP_mult_206_n2247, DP_mult_206_n2246, DP_mult_206_n2245,
         DP_mult_206_n2244, DP_mult_206_n2243, DP_mult_206_n2242,
         DP_mult_206_n2241, DP_mult_206_n2240, DP_mult_206_n2239,
         DP_mult_206_n2238, DP_mult_206_n2237, DP_mult_206_n2236,
         DP_mult_206_n2235, DP_mult_206_n2234, DP_mult_206_n2233,
         DP_mult_206_n2232, DP_mult_206_n2231, DP_mult_206_n2230,
         DP_mult_206_n2229, DP_mult_206_n2228, DP_mult_206_n2227,
         DP_mult_206_n2226, DP_mult_206_n2225, DP_mult_206_n2224,
         DP_mult_206_n2223, DP_mult_206_n2222, DP_mult_206_n2221,
         DP_mult_206_n2220, DP_mult_206_n2219, DP_mult_206_n2218,
         DP_mult_206_n2217, DP_mult_206_n2216, DP_mult_206_n2215,
         DP_mult_206_n2214, DP_mult_206_n2213, DP_mult_206_n2212,
         DP_mult_206_n2211, DP_mult_206_n2210, DP_mult_206_n2209,
         DP_mult_206_n2208, DP_mult_206_n2207, DP_mult_206_n2206,
         DP_mult_206_n2205, DP_mult_206_n2204, DP_mult_206_n2203,
         DP_mult_206_n2202, DP_mult_206_n2201, DP_mult_206_n2200,
         DP_mult_206_n2199, DP_mult_206_n2198, DP_mult_206_n2197,
         DP_mult_206_n2196, DP_mult_206_n2195, DP_mult_206_n2194,
         DP_mult_206_n2193, DP_mult_206_n2192, DP_mult_206_n2191,
         DP_mult_206_n2190, DP_mult_206_n2189, DP_mult_206_n2188,
         DP_mult_206_n2187, DP_mult_206_n2186, DP_mult_206_n2185,
         DP_mult_206_n2184, DP_mult_206_n2183, DP_mult_206_n2182,
         DP_mult_206_n2181, DP_mult_206_n2180, DP_mult_206_n2179,
         DP_mult_206_n2178, DP_mult_206_n2177, DP_mult_206_n2176,
         DP_mult_206_n2175, DP_mult_206_n2174, DP_mult_206_n2173,
         DP_mult_206_n2172, DP_mult_206_n2171, DP_mult_206_n2170,
         DP_mult_206_n2169, DP_mult_206_n2168, DP_mult_206_n2167,
         DP_mult_206_n2166, DP_mult_206_n2165, DP_mult_206_n2164,
         DP_mult_206_n2163, DP_mult_206_n2162, DP_mult_206_n2161,
         DP_mult_206_n2160, DP_mult_206_n2159, DP_mult_206_n2158,
         DP_mult_206_n2157, DP_mult_206_n2156, DP_mult_206_n2155,
         DP_mult_206_n2154, DP_mult_206_n2153, DP_mult_206_n2152,
         DP_mult_206_n2151, DP_mult_206_n2150, DP_mult_206_n2149,
         DP_mult_206_n2148, DP_mult_206_n2147, DP_mult_206_n2146,
         DP_mult_206_n2145, DP_mult_206_n2144, DP_mult_206_n2143,
         DP_mult_206_n2142, DP_mult_206_n2141, DP_mult_206_n2140,
         DP_mult_206_n2139, DP_mult_206_n2138, DP_mult_206_n2137,
         DP_mult_206_n2136, DP_mult_206_n2135, DP_mult_206_n2134,
         DP_mult_206_n2133, DP_mult_206_n2132, DP_mult_206_n2131,
         DP_mult_206_n2130, DP_mult_206_n2129, DP_mult_206_n2128,
         DP_mult_206_n2127, DP_mult_206_n2126, DP_mult_206_n2125,
         DP_mult_206_n2124, DP_mult_206_n2123, DP_mult_206_n2122,
         DP_mult_206_n2121, DP_mult_206_n2120, DP_mult_206_n2119,
         DP_mult_206_n2118, DP_mult_206_n2117, DP_mult_206_n2116,
         DP_mult_206_n2115, DP_mult_206_n2114, DP_mult_206_n2113,
         DP_mult_206_n2112, DP_mult_206_n2111, DP_mult_206_n2110,
         DP_mult_206_n2109, DP_mult_206_n2108, DP_mult_206_n2107,
         DP_mult_206_n2106, DP_mult_206_n2105, DP_mult_206_n2104,
         DP_mult_206_n2103, DP_mult_206_n2102, DP_mult_206_n2101,
         DP_mult_206_n2100, DP_mult_206_n2099, DP_mult_206_n2098,
         DP_mult_206_n2097, DP_mult_206_n2096, DP_mult_206_n2095,
         DP_mult_206_n2094, DP_mult_206_n2093, DP_mult_206_n2092,
         DP_mult_206_n2091, DP_mult_206_n2090, DP_mult_206_n2089,
         DP_mult_206_n2088, DP_mult_206_n2087, DP_mult_206_n2086,
         DP_mult_206_n2085, DP_mult_206_n2084, DP_mult_206_n2083,
         DP_mult_206_n2082, DP_mult_206_n2081, DP_mult_206_n2080,
         DP_mult_206_n2079, DP_mult_206_n2078, DP_mult_206_n2077,
         DP_mult_206_n2076, DP_mult_206_n2075, DP_mult_206_n2074,
         DP_mult_206_n2073, DP_mult_206_n2072, DP_mult_206_n2071,
         DP_mult_206_n2070, DP_mult_206_n2069, DP_mult_206_n2068,
         DP_mult_206_n2067, DP_mult_206_n2066, DP_mult_206_n2065,
         DP_mult_206_n2064, DP_mult_206_n2063, DP_mult_206_n2062,
         DP_mult_206_n2061, DP_mult_206_n2060, DP_mult_206_n2059,
         DP_mult_206_n2058, DP_mult_206_n2057, DP_mult_206_n2056,
         DP_mult_206_n2055, DP_mult_206_n2054, DP_mult_206_n2053,
         DP_mult_206_n2052, DP_mult_206_n2051, DP_mult_206_n2050,
         DP_mult_206_n2049, DP_mult_206_n2048, DP_mult_206_n2047,
         DP_mult_206_n2046, DP_mult_206_n2045, DP_mult_206_n2044,
         DP_mult_206_n2043, DP_mult_206_n2042, DP_mult_206_n2041,
         DP_mult_206_n2040, DP_mult_206_n2039, DP_mult_206_n2038,
         DP_mult_206_n2037, DP_mult_206_n2036, DP_mult_206_n2035,
         DP_mult_206_n2034, DP_mult_206_n2033, DP_mult_206_n2032,
         DP_mult_206_n2031, DP_mult_206_n2030, DP_mult_206_n2029,
         DP_mult_206_n2028, DP_mult_206_n2027, DP_mult_206_n2026,
         DP_mult_206_n2025, DP_mult_206_n2024, DP_mult_206_n2023,
         DP_mult_206_n2022, DP_mult_206_n2021, DP_mult_206_n2020,
         DP_mult_206_n2019, DP_mult_206_n2018, DP_mult_206_n2017,
         DP_mult_206_n2016, DP_mult_206_n2015, DP_mult_206_n2014,
         DP_mult_206_n2013, DP_mult_206_n2012, DP_mult_206_n2011,
         DP_mult_206_n2010, DP_mult_206_n2009, DP_mult_206_n2008,
         DP_mult_206_n2007, DP_mult_206_n2006, DP_mult_206_n2005,
         DP_mult_206_n2004, DP_mult_206_n2003, DP_mult_206_n2002,
         DP_mult_206_n2001, DP_mult_206_n2000, DP_mult_206_n1999,
         DP_mult_206_n1998, DP_mult_206_n1997, DP_mult_206_n1996,
         DP_mult_206_n1995, DP_mult_206_n1994, DP_mult_206_n1993,
         DP_mult_206_n1992, DP_mult_206_n1991, DP_mult_206_n1990,
         DP_mult_206_n1989, DP_mult_206_n1988, DP_mult_206_n1987,
         DP_mult_206_n1986, DP_mult_206_n1985, DP_mult_206_n1984,
         DP_mult_206_n1983, DP_mult_206_n1982, DP_mult_206_n1981,
         DP_mult_206_n1980, DP_mult_206_n1979, DP_mult_206_n1978,
         DP_mult_206_n1977, DP_mult_206_n1976, DP_mult_206_n1975,
         DP_mult_206_n1974, DP_mult_206_n1973, DP_mult_206_n1972,
         DP_mult_206_n1971, DP_mult_206_n1970, DP_mult_206_n1969,
         DP_mult_206_n1968, DP_mult_206_n1967, DP_mult_206_n1966,
         DP_mult_206_n1965, DP_mult_206_n1964, DP_mult_206_n1963,
         DP_mult_206_n1962, DP_mult_206_n1961, DP_mult_206_n1960,
         DP_mult_206_n1959, DP_mult_206_n1958, DP_mult_206_n1957,
         DP_mult_206_n1956, DP_mult_206_n1955, DP_mult_206_n1954,
         DP_mult_206_n1953, DP_mult_206_n1952, DP_mult_206_n1951,
         DP_mult_206_n1950, DP_mult_206_n1949, DP_mult_206_n1948,
         DP_mult_206_n1947, DP_mult_206_n1946, DP_mult_206_n1945,
         DP_mult_206_n1944, DP_mult_206_n1943, DP_mult_206_n1942,
         DP_mult_206_n1941, DP_mult_206_n1940, DP_mult_206_n1939,
         DP_mult_206_n1938, DP_mult_206_n1937, DP_mult_206_n1936,
         DP_mult_206_n1935, DP_mult_206_n1934, DP_mult_206_n1933,
         DP_mult_206_n1932, DP_mult_206_n1931, DP_mult_206_n1930,
         DP_mult_206_n1929, DP_mult_206_n1817, DP_mult_206_n1816,
         DP_mult_206_n1815, DP_mult_206_n1814, DP_mult_206_n1812,
         DP_mult_206_n1811, DP_mult_206_n1810, DP_mult_206_n1809,
         DP_mult_206_n1808, DP_mult_206_n1807, DP_mult_206_n1806,
         DP_mult_206_n1781, DP_mult_206_n1780, DP_mult_206_n1779,
         DP_mult_206_n1778, DP_mult_206_n1777, DP_mult_206_n1776,
         DP_mult_206_n1775, DP_mult_206_n1774, DP_mult_206_n1773,
         DP_mult_206_n1772, DP_mult_206_n1771, DP_mult_206_n1770,
         DP_mult_206_n1769, DP_mult_206_n1768, DP_mult_206_n1767,
         DP_mult_206_n1766, DP_mult_206_n1765, DP_mult_206_n1764,
         DP_mult_206_n1763, DP_mult_206_n1762, DP_mult_206_n1761,
         DP_mult_206_n1760, DP_mult_206_n1759, DP_mult_206_n1758,
         DP_mult_206_n1757, DP_mult_206_n1756, DP_mult_206_n1755,
         DP_mult_206_n1754, DP_mult_206_n1753, DP_mult_206_n1752,
         DP_mult_206_n1751, DP_mult_206_n1750, DP_mult_206_n1749,
         DP_mult_206_n1748, DP_mult_206_n1747, DP_mult_206_n1746,
         DP_mult_206_n1745, DP_mult_206_n1744, DP_mult_206_n1743,
         DP_mult_206_n1742, DP_mult_206_n1741, DP_mult_206_n1740,
         DP_mult_206_n1739, DP_mult_206_n1738, DP_mult_206_n1737,
         DP_mult_206_n1736, DP_mult_206_n1735, DP_mult_206_n1734,
         DP_mult_206_n1733, DP_mult_206_n1732, DP_mult_206_n1731,
         DP_mult_206_n1730, DP_mult_206_n1729, DP_mult_206_n1728,
         DP_mult_206_n1727, DP_mult_206_n1726, DP_mult_206_n1725,
         DP_mult_206_n1724, DP_mult_206_n1723, DP_mult_206_n1722,
         DP_mult_206_n1721, DP_mult_206_n1720, DP_mult_206_n1719,
         DP_mult_206_n1718, DP_mult_206_n1717, DP_mult_206_n1716,
         DP_mult_206_n1715, DP_mult_206_n1714, DP_mult_206_n1713,
         DP_mult_206_n1712, DP_mult_206_n1711, DP_mult_206_n1710,
         DP_mult_206_n1709, DP_mult_206_n1708, DP_mult_206_n1707,
         DP_mult_206_n1706, DP_mult_206_n1705, DP_mult_206_n1704,
         DP_mult_206_n1703, DP_mult_206_n1702, DP_mult_206_n1701,
         DP_mult_206_n1700, DP_mult_206_n1699, DP_mult_206_n1698,
         DP_mult_206_n1697, DP_mult_206_n1696, DP_mult_206_n1695,
         DP_mult_206_n1694, DP_mult_206_n1693, DP_mult_206_n1692,
         DP_mult_206_n1691, DP_mult_206_n1690, DP_mult_206_n1689,
         DP_mult_206_n1688, DP_mult_206_n1687, DP_mult_206_n1686,
         DP_mult_206_n1685, DP_mult_206_n1684, DP_mult_206_n1683,
         DP_mult_206_n1682, DP_mult_206_n1681, DP_mult_206_n1680,
         DP_mult_206_n1679, DP_mult_206_n1678, DP_mult_206_n1677,
         DP_mult_206_n1676, DP_mult_206_n1675, DP_mult_206_n1674,
         DP_mult_206_n1673, DP_mult_206_n1672, DP_mult_206_n1671,
         DP_mult_206_n1670, DP_mult_206_n1669, DP_mult_206_n1668,
         DP_mult_206_n1667, DP_mult_206_n1666, DP_mult_206_n1665,
         DP_mult_206_n1664, DP_mult_206_n1663, DP_mult_206_n1662,
         DP_mult_206_n1661, DP_mult_206_n1660, DP_mult_206_n1659,
         DP_mult_206_n1658, DP_mult_206_n1657, DP_mult_206_n1656,
         DP_mult_206_n1655, DP_mult_206_n1654, DP_mult_206_n1653,
         DP_mult_206_n1652, DP_mult_206_n1651, DP_mult_206_n1650,
         DP_mult_206_n1649, DP_mult_206_n1648, DP_mult_206_n1647,
         DP_mult_206_n1646, DP_mult_206_n1645, DP_mult_206_n1644,
         DP_mult_206_n1643, DP_mult_206_n1642, DP_mult_206_n1641,
         DP_mult_206_n1640, DP_mult_206_n1639, DP_mult_206_n1638,
         DP_mult_206_n1637, DP_mult_206_n1636, DP_mult_206_n1635,
         DP_mult_206_n1634, DP_mult_206_n1633, DP_mult_206_n1632,
         DP_mult_206_n1631, DP_mult_206_n1630, DP_mult_206_n1629,
         DP_mult_206_n1628, DP_mult_206_n1627, DP_mult_206_n1626,
         DP_mult_206_n1625, DP_mult_206_n1624, DP_mult_206_n1623,
         DP_mult_206_n1622, DP_mult_206_n1621, DP_mult_206_n1620,
         DP_mult_206_n1619, DP_mult_206_n1618, DP_mult_206_n1617,
         DP_mult_206_n1616, DP_mult_206_n1615, DP_mult_206_n1614,
         DP_mult_206_n1613, DP_mult_206_n1612, DP_mult_206_n1611,
         DP_mult_206_n1610, DP_mult_206_n1609, DP_mult_206_n1608,
         DP_mult_206_n1607, DP_mult_206_n1606, DP_mult_206_n1605,
         DP_mult_206_n1604, DP_mult_206_n1603, DP_mult_206_n1602,
         DP_mult_206_n1601, DP_mult_206_n1600, DP_mult_206_n1599,
         DP_mult_206_n1598, DP_mult_206_n1597, DP_mult_206_n1596,
         DP_mult_206_n1595, DP_mult_206_n1594, DP_mult_206_n1593,
         DP_mult_206_n1592, DP_mult_206_n1591, DP_mult_206_n1590,
         DP_mult_206_n1589, DP_mult_206_n1588, DP_mult_206_n1587,
         DP_mult_206_n1586, DP_mult_206_n1585, DP_mult_206_n1584,
         DP_mult_206_n1583, DP_mult_206_n1582, DP_mult_206_n1581,
         DP_mult_206_n1580, DP_mult_206_n1579, DP_mult_206_n1578,
         DP_mult_206_n1577, DP_mult_206_n1576, DP_mult_206_n1575,
         DP_mult_206_n1574, DP_mult_206_n1573, DP_mult_206_n1572,
         DP_mult_206_n1571, DP_mult_206_n1570, DP_mult_206_n1569,
         DP_mult_206_n1568, DP_mult_206_n1567, DP_mult_206_n1566,
         DP_mult_206_n1565, DP_mult_206_n1564, DP_mult_206_n1563,
         DP_mult_206_n1562, DP_mult_206_n1561, DP_mult_206_n1560,
         DP_mult_206_n1559, DP_mult_206_n1558, DP_mult_206_n1557,
         DP_mult_206_n1556, DP_mult_206_n1555, DP_mult_206_n1554,
         DP_mult_206_n1553, DP_mult_206_n1552, DP_mult_206_n1551,
         DP_mult_206_n1550, DP_mult_206_n1549, DP_mult_206_n1548,
         DP_mult_206_n1547, DP_mult_206_n1546, DP_mult_206_n1545,
         DP_mult_206_n1544, DP_mult_206_n1543, DP_mult_206_n1542,
         DP_mult_206_n1541, DP_mult_206_n1540, DP_mult_206_n1539,
         DP_mult_206_n1538, DP_mult_206_n1537, DP_mult_206_n1536,
         DP_mult_206_n1535, DP_mult_206_n1534, DP_mult_206_n1533,
         DP_mult_206_n1532, DP_mult_206_n1531, DP_mult_206_n1530,
         DP_mult_206_n1529, DP_mult_206_n1528, DP_mult_206_n1527,
         DP_mult_206_n1526, DP_mult_206_n1525, DP_mult_206_n1524,
         DP_mult_206_n1523, DP_mult_206_n1522, DP_mult_206_n1521,
         DP_mult_206_n1520, DP_mult_206_n1519, DP_mult_206_n1518,
         DP_mult_206_n1517, DP_mult_206_n1516, DP_mult_206_n1515,
         DP_mult_206_n1514, DP_mult_206_n1513, DP_mult_206_n1512,
         DP_mult_206_n1511, DP_mult_206_n1510, DP_mult_206_n1509,
         DP_mult_206_n1508, DP_mult_206_n1507, DP_mult_206_n1506,
         DP_mult_206_n1505, DP_mult_206_n1504, DP_mult_206_n1503,
         DP_mult_206_n1502, DP_mult_206_n1501, DP_mult_206_n1500,
         DP_mult_206_n1499, DP_mult_206_n1498, DP_mult_206_n1497,
         DP_mult_206_n1496, DP_mult_206_n1495, DP_mult_206_n1494,
         DP_mult_206_n1493, DP_mult_206_n1492, DP_mult_206_n1491,
         DP_mult_206_n1490, DP_mult_206_n1489, DP_mult_206_n1488,
         DP_mult_206_n1487, DP_mult_206_n1486, DP_mult_206_n1485,
         DP_mult_206_n1484, DP_mult_206_n1483, DP_mult_206_n1482,
         DP_mult_206_n1481, DP_mult_206_n1480, DP_mult_206_n1479,
         DP_mult_206_n1478, DP_mult_206_n1477, DP_mult_206_n1476,
         DP_mult_206_n1475, DP_mult_206_n1474, DP_mult_206_n1473,
         DP_mult_206_n1472, DP_mult_206_n1471, DP_mult_206_n1470,
         DP_mult_206_n1469, DP_mult_206_n1468, DP_mult_206_n1467,
         DP_mult_206_n1466, DP_mult_206_n1465, DP_mult_206_n1464,
         DP_mult_206_n1463, DP_mult_206_n1462, DP_mult_206_n1461,
         DP_mult_206_n1460, DP_mult_206_n1459, DP_mult_206_n1458,
         DP_mult_206_n1457, DP_mult_206_n1456, DP_mult_206_n1455,
         DP_mult_206_n1454, DP_mult_206_n1453, DP_mult_206_n1452,
         DP_mult_206_n1451, DP_mult_206_n1450, DP_mult_206_n1449,
         DP_mult_206_n1448, DP_mult_206_n1447, DP_mult_206_n1446,
         DP_mult_206_n1445, DP_mult_206_n1444, DP_mult_206_n1443,
         DP_mult_206_n1442, DP_mult_206_n1441, DP_mult_206_n1440,
         DP_mult_206_n1439, DP_mult_206_n1438, DP_mult_206_n1437,
         DP_mult_206_n1436, DP_mult_206_n1435, DP_mult_206_n1434,
         DP_mult_206_n1433, DP_mult_206_n1432, DP_mult_206_n1431,
         DP_mult_206_n1430, DP_mult_206_n1429, DP_mult_206_n1428,
         DP_mult_206_n1427, DP_mult_206_n1426, DP_mult_206_n1425,
         DP_mult_206_n1424, DP_mult_206_n1423, DP_mult_206_n1422,
         DP_mult_206_n1421, DP_mult_206_n1420, DP_mult_206_n1419,
         DP_mult_206_n1418, DP_mult_206_n1417, DP_mult_206_n1416,
         DP_mult_206_n1415, DP_mult_206_n1414, DP_mult_206_n1413,
         DP_mult_206_n1412, DP_mult_206_n1411, DP_mult_206_n1410,
         DP_mult_206_n1409, DP_mult_206_n1408, DP_mult_206_n1407,
         DP_mult_206_n1406, DP_mult_206_n1405, DP_mult_206_n1404,
         DP_mult_206_n1403, DP_mult_206_n1402, DP_mult_206_n1401,
         DP_mult_206_n1400, DP_mult_206_n1399, DP_mult_206_n1398,
         DP_mult_206_n1397, DP_mult_206_n1396, DP_mult_206_n1395,
         DP_mult_206_n1394, DP_mult_206_n1393, DP_mult_206_n1392,
         DP_mult_206_n1391, DP_mult_206_n1390, DP_mult_206_n1389,
         DP_mult_206_n1388, DP_mult_206_n1387, DP_mult_206_n1386,
         DP_mult_206_n1385, DP_mult_206_n1384, DP_mult_206_n1383,
         DP_mult_206_n1382, DP_mult_206_n1381, DP_mult_206_n1380,
         DP_mult_206_n1379, DP_mult_206_n1378, DP_mult_206_n1377,
         DP_mult_206_n1376, DP_mult_206_n1375, DP_mult_206_n1374,
         DP_mult_206_n1373, DP_mult_206_n1372, DP_mult_206_n1371,
         DP_mult_206_n1370, DP_mult_206_n1369, DP_mult_206_n1368,
         DP_mult_206_n1367, DP_mult_206_n1366, DP_mult_206_n1365,
         DP_mult_206_n1364, DP_mult_206_n1363, DP_mult_206_n1362,
         DP_mult_206_n1361, DP_mult_206_n1360, DP_mult_206_n1359,
         DP_mult_206_n1358, DP_mult_206_n1357, DP_mult_206_n1356,
         DP_mult_206_n1355, DP_mult_206_n1354, DP_mult_206_n1353,
         DP_mult_206_n1352, DP_mult_206_n1351, DP_mult_206_n1350,
         DP_mult_206_n1349, DP_mult_206_n1348, DP_mult_206_n1347,
         DP_mult_206_n1346, DP_mult_206_n1345, DP_mult_206_n1344,
         DP_mult_206_n1343, DP_mult_206_n1342, DP_mult_206_n1341,
         DP_mult_206_n1340, DP_mult_206_n1339, DP_mult_206_n1338,
         DP_mult_206_n1337, DP_mult_206_n1336, DP_mult_206_n1335,
         DP_mult_206_n1334, DP_mult_206_n1333, DP_mult_206_n1332,
         DP_mult_206_n1331, DP_mult_206_n1330, DP_mult_206_n1329,
         DP_mult_206_n1328, DP_mult_206_n1327, DP_mult_206_n1326,
         DP_mult_206_n1325, DP_mult_206_n1324, DP_mult_206_n1323,
         DP_mult_206_n1322, DP_mult_206_n1321, DP_mult_206_n1320,
         DP_mult_206_n1319, DP_mult_206_n1318, DP_mult_206_n1317,
         DP_mult_206_n1316, DP_mult_206_n1315, DP_mult_206_n1314,
         DP_mult_206_n1313, DP_mult_206_n1312, DP_mult_206_n1311,
         DP_mult_206_n1310, DP_mult_206_n1309, DP_mult_206_n1308,
         DP_mult_206_n1307, DP_mult_206_n1306, DP_mult_206_n1305,
         DP_mult_206_n1304, DP_mult_206_n1303, DP_mult_206_n1302,
         DP_mult_206_n1301, DP_mult_206_n1300, DP_mult_206_n1299,
         DP_mult_206_n1298, DP_mult_206_n1297, DP_mult_206_n1296,
         DP_mult_206_n1295, DP_mult_206_n1294, DP_mult_206_n1293,
         DP_mult_206_n1292, DP_mult_206_n1291, DP_mult_206_n1290,
         DP_mult_206_n1289, DP_mult_206_n1288, DP_mult_206_n1287,
         DP_mult_206_n1286, DP_mult_206_n1285, DP_mult_206_n1284,
         DP_mult_206_n1283, DP_mult_206_n1282, DP_mult_206_n1281,
         DP_mult_206_n1280, DP_mult_206_n1279, DP_mult_206_n1278,
         DP_mult_206_n1277, DP_mult_206_n1276, DP_mult_206_n1275,
         DP_mult_206_n1274, DP_mult_206_n1273, DP_mult_206_n1272,
         DP_mult_206_n1271, DP_mult_206_n1270, DP_mult_206_n1269,
         DP_mult_206_n1268, DP_mult_206_n1267, DP_mult_206_n1266,
         DP_mult_206_n1265, DP_mult_206_n1264, DP_mult_206_n1263,
         DP_mult_206_n1262, DP_mult_206_n1261, DP_mult_206_n1260,
         DP_mult_206_n1259, DP_mult_206_n1258, DP_mult_206_n1257,
         DP_mult_206_n1256, DP_mult_206_n1255, DP_mult_206_n1254,
         DP_mult_206_n1253, DP_mult_206_n1252, DP_mult_206_n1251,
         DP_mult_206_n1250, DP_mult_206_n1249, DP_mult_206_n1248,
         DP_mult_206_n1247, DP_mult_206_n1246, DP_mult_206_n1245,
         DP_mult_206_n1244, DP_mult_206_n1243, DP_mult_206_n1242,
         DP_mult_206_n1241, DP_mult_206_n1240, DP_mult_206_n1239,
         DP_mult_206_n1238, DP_mult_206_n1237, DP_mult_206_n1236,
         DP_mult_206_n1235, DP_mult_206_n1234, DP_mult_206_n1233,
         DP_mult_206_n1232, DP_mult_206_n1231, DP_mult_206_n1230,
         DP_mult_206_n1229, DP_mult_206_n1228, DP_mult_206_n1227,
         DP_mult_206_n1226, DP_mult_206_n1225, DP_mult_206_n1224,
         DP_mult_206_n1223, DP_mult_206_n1222, DP_mult_206_n1221,
         DP_mult_206_n1220, DP_mult_206_n1219, DP_mult_206_n1218,
         DP_mult_206_n1217, DP_mult_206_n1216, DP_mult_206_n1215,
         DP_mult_206_n1214, DP_mult_206_n1213, DP_mult_206_n1212,
         DP_mult_206_n1211, DP_mult_206_n1210, DP_mult_206_n1209,
         DP_mult_206_n1208, DP_mult_206_n1207, DP_mult_206_n1206,
         DP_mult_206_n1205, DP_mult_206_n1204, DP_mult_206_n1203,
         DP_mult_206_n1202, DP_mult_206_n1201, DP_mult_206_n1200,
         DP_mult_206_n1199, DP_mult_206_n1198, DP_mult_206_n1197,
         DP_mult_206_n1196, DP_mult_206_n1195, DP_mult_206_n1194,
         DP_mult_206_n1193, DP_mult_206_n1192, DP_mult_206_n1191,
         DP_mult_206_n1190, DP_mult_206_n1189, DP_mult_206_n1188,
         DP_mult_206_n1187, DP_mult_206_n1186, DP_mult_206_n1185,
         DP_mult_206_n1184, DP_mult_206_n1183, DP_mult_206_n1182,
         DP_mult_206_n1181, DP_mult_206_n1180, DP_mult_206_n1179,
         DP_mult_206_n1178, DP_mult_206_n1177, DP_mult_206_n1176,
         DP_mult_206_n1175, DP_mult_206_n1174, DP_mult_206_n1173,
         DP_mult_206_n1172, DP_mult_206_n1171, DP_mult_206_n1170,
         DP_mult_206_n1169, DP_mult_206_n1168, DP_mult_206_n1167,
         DP_mult_206_n1166, DP_mult_206_n1165, DP_mult_206_n1164,
         DP_mult_206_n1163, DP_mult_206_n1162, DP_mult_206_n1161,
         DP_mult_206_n1160, DP_mult_206_n1159, DP_mult_206_n1158,
         DP_mult_206_n1157, DP_mult_206_n1156, DP_mult_206_n1155,
         DP_mult_206_n1154, DP_mult_206_n1153, DP_mult_206_n1152,
         DP_mult_206_n1151, DP_mult_206_n1150, DP_mult_206_n1149,
         DP_mult_206_n1148, DP_mult_206_n1147, DP_mult_206_n1146,
         DP_mult_206_n1145, DP_mult_206_n1144, DP_mult_206_n1143,
         DP_mult_206_n1142, DP_mult_206_n1141, DP_mult_206_n1140,
         DP_mult_206_n1139, DP_mult_206_n1138, DP_mult_206_n1137,
         DP_mult_206_n1136, DP_mult_206_n1135, DP_mult_206_n1134,
         DP_mult_206_n1133, DP_mult_206_n1132, DP_mult_206_n1131,
         DP_mult_206_n1130, DP_mult_206_n1129, DP_mult_206_n1128,
         DP_mult_206_n1127, DP_mult_206_n1126, DP_mult_206_n1125,
         DP_mult_206_n1124, DP_mult_206_n1123, DP_mult_206_n1122,
         DP_mult_206_n1121, DP_mult_206_n1120, DP_mult_206_n1119,
         DP_mult_206_n1118, DP_mult_206_n1117, DP_mult_206_n1116,
         DP_mult_206_n1115, DP_mult_206_n1114, DP_mult_206_n1113,
         DP_mult_206_n1112, DP_mult_206_n1111, DP_mult_206_n1110,
         DP_mult_206_n1109, DP_mult_206_n1108, DP_mult_206_n1107,
         DP_mult_206_n1106, DP_mult_206_n1105, DP_mult_206_n1104,
         DP_mult_206_n1103, DP_mult_206_n1102, DP_mult_206_n1101,
         DP_mult_206_n1100, DP_mult_206_n1099, DP_mult_206_n1098,
         DP_mult_206_n1097, DP_mult_206_n1096, DP_mult_206_n1095,
         DP_mult_206_n1094, DP_mult_206_n1093, DP_mult_206_n1092,
         DP_mult_206_n1091, DP_mult_206_n1090, DP_mult_206_n1089,
         DP_mult_206_n1088, DP_mult_206_n1087, DP_mult_206_n1086,
         DP_mult_206_n1085, DP_mult_206_n1084, DP_mult_206_n1083,
         DP_mult_206_n1082, DP_mult_206_n1081, DP_mult_206_n1080,
         DP_mult_206_n1079, DP_mult_206_n1078, DP_mult_206_n1077,
         DP_mult_206_n1076, DP_mult_206_n1075, DP_mult_206_n1074,
         DP_mult_206_n1073, DP_mult_206_n1072, DP_mult_206_n1071,
         DP_mult_206_n1070, DP_mult_206_n1069, DP_mult_206_n1068,
         DP_mult_206_n1067, DP_mult_206_n1066, DP_mult_206_n1065,
         DP_mult_206_n1064, DP_mult_206_n1063, DP_mult_206_n1062,
         DP_mult_206_n1061, DP_mult_206_n1060, DP_mult_206_n1059,
         DP_mult_206_n1058, DP_mult_206_n1057, DP_mult_206_n1056,
         DP_mult_206_n1055, DP_mult_206_n1054, DP_mult_206_n1053,
         DP_mult_206_n1052, DP_mult_206_n1051, DP_mult_206_n1050,
         DP_mult_206_n1049, DP_mult_206_n1048, DP_mult_206_n1047,
         DP_mult_206_n1046, DP_mult_206_n1045, DP_mult_206_n1044,
         DP_mult_206_n1043, DP_mult_206_n1042, DP_mult_206_n1041,
         DP_mult_206_n1040, DP_mult_206_n1039, DP_mult_206_n1038,
         DP_mult_206_n1037, DP_mult_206_n1036, DP_mult_206_n1035,
         DP_mult_206_n1034, DP_mult_206_n1033, DP_mult_206_n1032,
         DP_mult_206_n1031, DP_mult_206_n1030, DP_mult_206_n1029,
         DP_mult_206_n1028, DP_mult_206_n1027, DP_mult_206_n1026,
         DP_mult_206_n1025, DP_mult_206_n1024, DP_mult_206_n1023,
         DP_mult_206_n1022, DP_mult_206_n1021, DP_mult_206_n1020,
         DP_mult_206_n1019, DP_mult_206_n1018, DP_mult_206_n1017,
         DP_mult_206_n1016, DP_mult_206_n1015, DP_mult_206_n1014,
         DP_mult_206_n1013, DP_mult_206_n1012, DP_mult_206_n1011,
         DP_mult_206_n1010, DP_mult_206_n1009, DP_mult_206_n1008,
         DP_mult_206_n1007, DP_mult_206_n1006, DP_mult_206_n1005,
         DP_mult_206_n1004, DP_mult_206_n1003, DP_mult_206_n1002,
         DP_mult_206_n1001, DP_mult_206_n1000, DP_mult_206_n999,
         DP_mult_206_n998, DP_mult_206_n997, DP_mult_206_n996,
         DP_mult_206_n995, DP_mult_206_n994, DP_mult_206_n993,
         DP_mult_206_n992, DP_mult_206_n991, DP_mult_206_n990,
         DP_mult_206_n989, DP_mult_206_n988, DP_mult_206_n987,
         DP_mult_206_n986, DP_mult_206_n985, DP_mult_206_n984,
         DP_mult_206_n983, DP_mult_206_n982, DP_mult_206_n981,
         DP_mult_206_n980, DP_mult_206_n979, DP_mult_206_n978,
         DP_mult_206_n977, DP_mult_206_n976, DP_mult_206_n975,
         DP_mult_206_n974, DP_mult_206_n973, DP_mult_206_n972,
         DP_mult_206_n971, DP_mult_206_n970, DP_mult_206_n969,
         DP_mult_206_n968, DP_mult_206_n967, DP_mult_206_n966,
         DP_mult_206_n965, DP_mult_206_n964, DP_mult_206_n963,
         DP_mult_206_n962, DP_mult_206_n961, DP_mult_206_n960,
         DP_mult_206_n959, DP_mult_206_n957, DP_mult_206_n956,
         DP_mult_206_n955, DP_mult_206_n954, DP_mult_206_n953,
         DP_mult_206_n952, DP_mult_206_n951, DP_mult_206_n950,
         DP_mult_206_n949, DP_mult_206_n948, DP_mult_206_n947,
         DP_mult_206_n946, DP_mult_206_n945, DP_mult_206_n944,
         DP_mult_206_n943, DP_mult_206_n942, DP_mult_206_n941,
         DP_mult_206_n940, DP_mult_206_n939, DP_mult_206_n938,
         DP_mult_206_n937, DP_mult_206_n936, DP_mult_206_n935,
         DP_mult_206_n934, DP_mult_206_n933, DP_mult_206_n932,
         DP_mult_206_n931, DP_mult_206_n930, DP_mult_206_n929,
         DP_mult_206_n928, DP_mult_206_n927, DP_mult_206_n926,
         DP_mult_206_n925, DP_mult_206_n924, DP_mult_206_n923,
         DP_mult_206_n922, DP_mult_206_n921, DP_mult_206_n920,
         DP_mult_206_n919, DP_mult_206_n918, DP_mult_206_n917,
         DP_mult_206_n915, DP_mult_206_n914, DP_mult_206_n913,
         DP_mult_206_n912, DP_mult_206_n911, DP_mult_206_n910,
         DP_mult_206_n909, DP_mult_206_n908, DP_mult_206_n907,
         DP_mult_206_n906, DP_mult_206_n905, DP_mult_206_n904,
         DP_mult_206_n903, DP_mult_206_n902, DP_mult_206_n901,
         DP_mult_206_n900, DP_mult_206_n899, DP_mult_206_n898,
         DP_mult_206_n897, DP_mult_206_n896, DP_mult_206_n895,
         DP_mult_206_n894, DP_mult_206_n893, DP_mult_206_n892,
         DP_mult_206_n891, DP_mult_206_n890, DP_mult_206_n889,
         DP_mult_206_n888, DP_mult_206_n887, DP_mult_206_n886,
         DP_mult_206_n885, DP_mult_206_n884, DP_mult_206_n883,
         DP_mult_206_n882, DP_mult_206_n881, DP_mult_206_n880,
         DP_mult_206_n879, DP_mult_206_n878, DP_mult_206_n877,
         DP_mult_206_n876, DP_mult_206_n875, DP_mult_206_n874,
         DP_mult_206_n873, DP_mult_206_n872, DP_mult_206_n871,
         DP_mult_206_n870, DP_mult_206_n869, DP_mult_206_n868,
         DP_mult_206_n867, DP_mult_206_n866, DP_mult_206_n865,
         DP_mult_206_n864, DP_mult_206_n863, DP_mult_206_n861,
         DP_mult_206_n860, DP_mult_206_n859, DP_mult_206_n858,
         DP_mult_206_n857, DP_mult_206_n856, DP_mult_206_n855,
         DP_mult_206_n854, DP_mult_206_n853, DP_mult_206_n852,
         DP_mult_206_n851, DP_mult_206_n850, DP_mult_206_n849,
         DP_mult_206_n848, DP_mult_206_n847, DP_mult_206_n846,
         DP_mult_206_n845, DP_mult_206_n844, DP_mult_206_n843,
         DP_mult_206_n842, DP_mult_206_n841, DP_mult_206_n840,
         DP_mult_206_n839, DP_mult_206_n838, DP_mult_206_n836,
         DP_mult_206_n835, DP_mult_206_n834, DP_mult_206_n833,
         DP_mult_206_n832, DP_mult_206_n831, DP_mult_206_n830,
         DP_mult_206_n829, DP_mult_206_n828, DP_mult_206_n827,
         DP_mult_206_n826, DP_mult_206_n825, DP_mult_206_n824,
         DP_mult_206_n823, DP_mult_206_n822, DP_mult_206_n821,
         DP_mult_206_n820, DP_mult_206_n819, DP_mult_206_n818,
         DP_mult_206_n817, DP_mult_206_n816, DP_mult_206_n815,
         DP_mult_206_n814, DP_mult_206_n813, DP_mult_206_n812,
         DP_mult_206_n811, DP_mult_206_n810, DP_mult_206_n809,
         DP_mult_206_n808, DP_mult_206_n807, DP_mult_206_n806,
         DP_mult_206_n805, DP_mult_206_n804, DP_mult_206_n803,
         DP_mult_206_n802, DP_mult_206_n801, DP_mult_206_n800,
         DP_mult_206_n799, DP_mult_206_n798, DP_mult_206_n797,
         DP_mult_206_n796, DP_mult_206_n795, DP_mult_206_n794,
         DP_mult_206_n793, DP_mult_206_n792, DP_mult_206_n791,
         DP_mult_206_n790, DP_mult_206_n789, DP_mult_206_n788,
         DP_mult_206_n787, DP_mult_206_n786, DP_mult_206_n785,
         DP_mult_206_n784, DP_mult_206_n783, DP_mult_206_n782,
         DP_mult_206_n781, DP_mult_206_n780, DP_mult_206_n779,
         DP_mult_206_n778, DP_mult_206_n777, DP_mult_206_n776,
         DP_mult_206_n775, DP_mult_206_n774, DP_mult_206_n773,
         DP_mult_206_n772, DP_mult_206_n771, DP_mult_206_n770,
         DP_mult_206_n769, DP_mult_206_n768, DP_mult_206_n767,
         DP_mult_206_n766, DP_mult_206_n765, DP_mult_206_n764,
         DP_mult_206_n763, DP_mult_206_n762, DP_mult_206_n761,
         DP_mult_206_n760, DP_mult_206_n759, DP_mult_206_n758,
         DP_mult_206_n757, DP_mult_206_n756, DP_mult_206_n755,
         DP_mult_206_n754, DP_mult_206_n753, DP_mult_206_n752,
         DP_mult_206_n751, DP_mult_206_n750, DP_mult_206_n749,
         DP_mult_206_n748, DP_mult_206_n747, DP_mult_206_n746,
         DP_mult_206_n745, DP_mult_206_n744, DP_mult_206_n743,
         DP_mult_206_n742, DP_mult_206_n741, DP_mult_206_n740,
         DP_mult_206_n739, DP_mult_206_n738, DP_mult_206_n737,
         DP_mult_206_n736, DP_mult_206_n735, DP_mult_206_n734,
         DP_mult_206_n733, DP_mult_206_n732, DP_mult_206_n731,
         DP_mult_206_n730, DP_mult_206_n729, DP_mult_206_n728,
         DP_mult_206_n727, DP_mult_206_n726, DP_mult_206_n725,
         DP_mult_206_n724, DP_mult_206_n723, DP_mult_206_n722,
         DP_mult_206_n721, DP_mult_206_n720, DP_mult_206_n719,
         DP_mult_206_n718, DP_mult_206_n717, DP_mult_206_n716,
         DP_mult_206_n715, DP_mult_206_n714, DP_mult_206_n713,
         DP_mult_206_n712, DP_mult_206_n711, DP_mult_206_n710,
         DP_mult_206_n709, DP_mult_206_n708, DP_mult_206_n707,
         DP_mult_206_n706, DP_mult_206_n705, DP_mult_206_n704,
         DP_mult_206_n703, DP_mult_206_n702, DP_mult_206_n701,
         DP_mult_206_n700, DP_mult_206_n699, DP_mult_206_n698,
         DP_mult_206_n697, DP_mult_206_n696, DP_mult_206_n695,
         DP_mult_206_n694, DP_mult_206_n693, DP_mult_206_n692,
         DP_mult_206_n691, DP_mult_206_n690, DP_mult_206_n689,
         DP_mult_206_n688, DP_mult_206_n687, DP_mult_206_n686,
         DP_mult_206_n685, DP_mult_206_n684, DP_mult_206_n683,
         DP_mult_206_n682, DP_mult_206_n681, DP_mult_206_n680,
         DP_mult_206_n679, DP_mult_206_n678, DP_mult_206_n677,
         DP_mult_206_n676, DP_mult_206_n674, DP_mult_206_n673,
         DP_mult_206_n671, DP_mult_206_n670, DP_mult_206_n668,
         DP_mult_206_n667, DP_mult_206_n666, DP_mult_206_n663,
         DP_mult_206_n662, DP_mult_206_n661, DP_mult_206_n657,
         DP_mult_206_n646, DP_mult_206_n645, DP_mult_206_n644,
         DP_mult_206_n643, DP_mult_206_n638, DP_mult_206_n637,
         DP_mult_206_n636, DP_mult_206_n635, DP_mult_206_n634,
         DP_mult_206_n633, DP_mult_206_n632, DP_mult_206_n631,
         DP_mult_206_n630, DP_mult_206_n629, DP_mult_206_n628,
         DP_mult_206_n627, DP_mult_206_n626, DP_mult_206_n625,
         DP_mult_206_n620, DP_mult_206_n611, DP_mult_206_n610,
         DP_mult_206_n609, DP_mult_206_n600, DP_mult_206_n599,
         DP_mult_206_n598, DP_mult_206_n597, DP_mult_206_n596,
         DP_mult_206_n595, DP_mult_206_n594, DP_mult_206_n593,
         DP_mult_206_n592, DP_mult_206_n591, DP_mult_206_n590,
         DP_mult_206_n589, DP_mult_206_n588, DP_mult_206_n583,
         DP_mult_206_n582, DP_mult_206_n581, DP_mult_206_n572,
         DP_mult_206_n571, DP_mult_206_n570, DP_mult_206_n569,
         DP_mult_206_n568, DP_mult_206_n567, DP_mult_206_n566,
         DP_mult_206_n565, DP_mult_206_n564, DP_mult_206_n563,
         DP_mult_206_n562, DP_mult_206_n561, DP_mult_206_n560,
         DP_mult_206_n559, DP_mult_206_n558, DP_mult_206_n555,
         DP_mult_206_n553, DP_mult_206_n552, DP_mult_206_n551,
         DP_mult_206_n550, DP_mult_206_n547, DP_mult_206_n546,
         DP_mult_206_n545, DP_mult_206_n544, DP_mult_206_n543,
         DP_mult_206_n542, DP_mult_206_n541, DP_mult_206_n540,
         DP_mult_206_n539, DP_mult_206_n538, DP_mult_206_n537,
         DP_mult_206_n536, DP_mult_206_n535, DP_mult_206_n534,
         DP_mult_206_n533, DP_mult_206_n532, DP_mult_206_n531,
         DP_mult_206_n526, DP_mult_206_n525, DP_mult_206_n524,
         DP_mult_206_n523, DP_mult_206_n522, DP_mult_206_n521,
         DP_mult_206_n520, DP_mult_206_n519, DP_mult_206_n517,
         DP_mult_206_n516, DP_mult_206_n515, DP_mult_206_n514,
         DP_mult_206_n513, DP_mult_206_n512, DP_mult_206_n511,
         DP_mult_206_n508, DP_mult_206_n507, DP_mult_206_n506,
         DP_mult_206_n505, DP_mult_206_n504, DP_mult_206_n503,
         DP_mult_206_n502, DP_mult_206_n501, DP_mult_206_n499,
         DP_mult_206_n498, DP_mult_206_n497, DP_mult_206_n496,
         DP_mult_206_n495, DP_mult_206_n492, DP_mult_206_n491,
         DP_mult_206_n490, DP_mult_206_n489, DP_mult_206_n488,
         DP_mult_206_n487, DP_mult_206_n486, DP_mult_206_n483,
         DP_mult_206_n481, DP_mult_206_n480, DP_mult_206_n479,
         DP_mult_206_n478, DP_mult_206_n477, DP_mult_206_n476,
         DP_mult_206_n475, DP_mult_206_n474, DP_mult_206_n472,
         DP_mult_206_n468, DP_mult_206_n467, DP_mult_206_n466,
         DP_mult_206_n465, DP_mult_206_n464, DP_mult_206_n463,
         DP_mult_206_n462, DP_mult_206_n461, DP_mult_206_n459,
         DP_mult_206_n457, DP_mult_206_n456, DP_mult_206_n455,
         DP_mult_206_n454, DP_mult_206_n453, DP_mult_206_n452,
         DP_mult_206_n451, DP_mult_206_n450, DP_mult_206_n448,
         DP_mult_206_n445, DP_mult_206_n439, DP_mult_206_n438,
         DP_mult_206_n437, DP_mult_206_n436, DP_mult_206_n435,
         DP_mult_206_n434, DP_mult_206_n432, DP_mult_206_n431,
         DP_mult_206_n430, DP_mult_206_n429, DP_mult_206_n428,
         DP_mult_206_n427, DP_mult_206_n426, DP_mult_206_n423,
         DP_mult_206_n422, DP_mult_206_n421, DP_mult_206_n420,
         DP_mult_206_n419, DP_mult_206_n418, DP_mult_206_n416,
         DP_mult_206_n412, DP_mult_206_n411, DP_mult_206_n410,
         DP_mult_206_n409, DP_mult_206_n407, DP_mult_206_n405,
         DP_mult_206_n402, DP_mult_206_n401, DP_mult_206_n400,
         DP_mult_206_n399, DP_mult_206_n398, DP_mult_206_n397,
         DP_mult_206_n396, DP_mult_206_n394, DP_mult_206_n390,
         DP_mult_206_n389, DP_mult_206_n388, DP_mult_206_n387,
         DP_mult_206_n384, DP_mult_206_n383, DP_mult_206_n382,
         DP_mult_206_n381, DP_mult_206_n380, DP_mult_206_n379,
         DP_mult_206_n378, DP_mult_206_n376, DP_mult_206_n372,
         DP_mult_206_n371, DP_mult_206_n370, DP_mult_206_n369,
         DP_mult_206_n367, DP_mult_206_n365, DP_mult_206_n364,
         DP_mult_206_n363, DP_mult_206_n362, DP_mult_206_n361,
         DP_mult_206_n360, DP_mult_206_n359, DP_mult_206_n356,
         DP_mult_206_n355, DP_mult_206_n354, DP_mult_206_n353,
         DP_mult_206_n352, DP_mult_206_n350, DP_mult_206_n348,
         DP_mult_206_n347, DP_mult_206_n346, DP_mult_206_n345,
         DP_mult_206_n344, DP_mult_206_n343, DP_mult_206_n342,
         DP_mult_206_n341, DP_mult_206_n339, DP_mult_206_n337,
         DP_mult_206_n336, DP_mult_206_n335, DP_mult_206_n334,
         DP_mult_206_n333, DP_mult_206_n332, DP_mult_206_n327,
         DP_mult_206_n326, DP_mult_206_n325, DP_mult_206_n320,
         DP_mult_206_n319, DP_mult_206_n318, DP_mult_206_n317,
         DP_mult_206_n316, DP_mult_206_n315, DP_mult_206_n314,
         DP_mult_206_n313, DP_mult_206_n312, DP_mult_206_n311,
         DP_mult_206_n310, DP_mult_206_n309, DP_mult_206_n308,
         DP_mult_206_n307, DP_mult_206_n306, DP_mult_206_n305,
         DP_mult_206_n304, DP_mult_206_n303, DP_mult_206_n302,
         DP_mult_206_n301, DP_mult_206_n285, DP_mult_206_n253,
         DP_mult_206_n251, DP_mult_207_n2331, DP_mult_207_n2330,
         DP_mult_207_n2329, DP_mult_207_n2328, DP_mult_207_n2327,
         DP_mult_207_n2326, DP_mult_207_n2325, DP_mult_207_n2324,
         DP_mult_207_n2323, DP_mult_207_n2322, DP_mult_207_n2321,
         DP_mult_207_n2320, DP_mult_207_n2319, DP_mult_207_n2318,
         DP_mult_207_n2317, DP_mult_207_n2316, DP_mult_207_n2315,
         DP_mult_207_n2314, DP_mult_207_n2313, DP_mult_207_n2312,
         DP_mult_207_n2311, DP_mult_207_n2310, DP_mult_207_n2309,
         DP_mult_207_n2308, DP_mult_207_n2307, DP_mult_207_n2306,
         DP_mult_207_n2305, DP_mult_207_n2304, DP_mult_207_n2303,
         DP_mult_207_n2302, DP_mult_207_n2301, DP_mult_207_n2300,
         DP_mult_207_n2299, DP_mult_207_n2298, DP_mult_207_n2297,
         DP_mult_207_n2296, DP_mult_207_n2295, DP_mult_207_n2294,
         DP_mult_207_n2293, DP_mult_207_n2292, DP_mult_207_n2291,
         DP_mult_207_n2290, DP_mult_207_n2289, DP_mult_207_n2288,
         DP_mult_207_n2287, DP_mult_207_n2286, DP_mult_207_n2285,
         DP_mult_207_n2284, DP_mult_207_n2283, DP_mult_207_n2282,
         DP_mult_207_n2281, DP_mult_207_n2280, DP_mult_207_n2279,
         DP_mult_207_n2278, DP_mult_207_n2277, DP_mult_207_n2276,
         DP_mult_207_n2275, DP_mult_207_n2274, DP_mult_207_n2273,
         DP_mult_207_n2272, DP_mult_207_n2271, DP_mult_207_n2270,
         DP_mult_207_n2269, DP_mult_207_n2268, DP_mult_207_n2267,
         DP_mult_207_n2266, DP_mult_207_n2265, DP_mult_207_n2264,
         DP_mult_207_n2263, DP_mult_207_n2262, DP_mult_207_n2261,
         DP_mult_207_n2260, DP_mult_207_n2259, DP_mult_207_n2258,
         DP_mult_207_n2257, DP_mult_207_n2256, DP_mult_207_n2255,
         DP_mult_207_n2254, DP_mult_207_n2253, DP_mult_207_n2252,
         DP_mult_207_n2251, DP_mult_207_n2250, DP_mult_207_n2249,
         DP_mult_207_n2248, DP_mult_207_n2247, DP_mult_207_n2246,
         DP_mult_207_n2245, DP_mult_207_n2244, DP_mult_207_n2243,
         DP_mult_207_n2242, DP_mult_207_n2241, DP_mult_207_n2240,
         DP_mult_207_n2239, DP_mult_207_n2238, DP_mult_207_n2237,
         DP_mult_207_n2236, DP_mult_207_n2235, DP_mult_207_n2234,
         DP_mult_207_n2233, DP_mult_207_n2232, DP_mult_207_n2231,
         DP_mult_207_n2230, DP_mult_207_n2229, DP_mult_207_n2228,
         DP_mult_207_n2227, DP_mult_207_n2226, DP_mult_207_n2225,
         DP_mult_207_n2224, DP_mult_207_n2223, DP_mult_207_n2222,
         DP_mult_207_n2221, DP_mult_207_n2220, DP_mult_207_n2219,
         DP_mult_207_n2218, DP_mult_207_n2217, DP_mult_207_n2216,
         DP_mult_207_n2215, DP_mult_207_n2214, DP_mult_207_n2213,
         DP_mult_207_n2212, DP_mult_207_n2211, DP_mult_207_n2210,
         DP_mult_207_n2209, DP_mult_207_n2208, DP_mult_207_n2207,
         DP_mult_207_n2206, DP_mult_207_n2205, DP_mult_207_n2204,
         DP_mult_207_n2203, DP_mult_207_n2202, DP_mult_207_n2201,
         DP_mult_207_n2200, DP_mult_207_n2199, DP_mult_207_n2198,
         DP_mult_207_n2197, DP_mult_207_n2196, DP_mult_207_n2195,
         DP_mult_207_n2194, DP_mult_207_n2193, DP_mult_207_n2192,
         DP_mult_207_n2191, DP_mult_207_n2190, DP_mult_207_n2189,
         DP_mult_207_n2188, DP_mult_207_n2187, DP_mult_207_n2186,
         DP_mult_207_n2185, DP_mult_207_n2184, DP_mult_207_n2183,
         DP_mult_207_n2182, DP_mult_207_n2181, DP_mult_207_n2180,
         DP_mult_207_n2179, DP_mult_207_n2178, DP_mult_207_n2177,
         DP_mult_207_n2176, DP_mult_207_n2175, DP_mult_207_n2174,
         DP_mult_207_n2173, DP_mult_207_n2172, DP_mult_207_n2171,
         DP_mult_207_n2170, DP_mult_207_n2169, DP_mult_207_n2168,
         DP_mult_207_n2167, DP_mult_207_n2166, DP_mult_207_n2165,
         DP_mult_207_n2164, DP_mult_207_n2163, DP_mult_207_n2162,
         DP_mult_207_n2161, DP_mult_207_n2160, DP_mult_207_n2159,
         DP_mult_207_n2158, DP_mult_207_n2157, DP_mult_207_n2156,
         DP_mult_207_n2155, DP_mult_207_n2154, DP_mult_207_n2153,
         DP_mult_207_n2152, DP_mult_207_n2151, DP_mult_207_n2150,
         DP_mult_207_n2149, DP_mult_207_n2148, DP_mult_207_n2147,
         DP_mult_207_n2146, DP_mult_207_n2145, DP_mult_207_n2144,
         DP_mult_207_n2143, DP_mult_207_n2142, DP_mult_207_n2141,
         DP_mult_207_n2140, DP_mult_207_n2139, DP_mult_207_n2138,
         DP_mult_207_n2137, DP_mult_207_n2136, DP_mult_207_n2135,
         DP_mult_207_n2134, DP_mult_207_n2133, DP_mult_207_n2132,
         DP_mult_207_n2131, DP_mult_207_n2130, DP_mult_207_n2129,
         DP_mult_207_n2128, DP_mult_207_n2127, DP_mult_207_n2126,
         DP_mult_207_n2125, DP_mult_207_n2124, DP_mult_207_n2123,
         DP_mult_207_n2122, DP_mult_207_n2121, DP_mult_207_n2120,
         DP_mult_207_n2119, DP_mult_207_n2118, DP_mult_207_n2117,
         DP_mult_207_n2116, DP_mult_207_n2115, DP_mult_207_n2114,
         DP_mult_207_n2113, DP_mult_207_n2112, DP_mult_207_n2111,
         DP_mult_207_n2110, DP_mult_207_n2109, DP_mult_207_n2108,
         DP_mult_207_n2107, DP_mult_207_n2106, DP_mult_207_n2105,
         DP_mult_207_n2104, DP_mult_207_n2103, DP_mult_207_n2102,
         DP_mult_207_n2101, DP_mult_207_n2100, DP_mult_207_n2099,
         DP_mult_207_n2098, DP_mult_207_n2097, DP_mult_207_n2096,
         DP_mult_207_n2095, DP_mult_207_n2094, DP_mult_207_n2093,
         DP_mult_207_n2092, DP_mult_207_n2091, DP_mult_207_n2090,
         DP_mult_207_n2089, DP_mult_207_n2088, DP_mult_207_n2087,
         DP_mult_207_n2086, DP_mult_207_n2085, DP_mult_207_n2084,
         DP_mult_207_n2083, DP_mult_207_n2082, DP_mult_207_n2081,
         DP_mult_207_n2080, DP_mult_207_n2079, DP_mult_207_n2078,
         DP_mult_207_n2077, DP_mult_207_n2076, DP_mult_207_n2075,
         DP_mult_207_n2074, DP_mult_207_n2073, DP_mult_207_n2072,
         DP_mult_207_n2071, DP_mult_207_n2070, DP_mult_207_n2069,
         DP_mult_207_n2068, DP_mult_207_n2067, DP_mult_207_n2066,
         DP_mult_207_n2065, DP_mult_207_n2064, DP_mult_207_n2063,
         DP_mult_207_n2062, DP_mult_207_n2061, DP_mult_207_n2060,
         DP_mult_207_n2059, DP_mult_207_n2058, DP_mult_207_n2057,
         DP_mult_207_n2056, DP_mult_207_n2055, DP_mult_207_n2054,
         DP_mult_207_n2053, DP_mult_207_n2052, DP_mult_207_n2051,
         DP_mult_207_n2050, DP_mult_207_n2049, DP_mult_207_n2048,
         DP_mult_207_n2047, DP_mult_207_n2046, DP_mult_207_n2045,
         DP_mult_207_n2044, DP_mult_207_n2043, DP_mult_207_n2042,
         DP_mult_207_n2041, DP_mult_207_n2040, DP_mult_207_n2039,
         DP_mult_207_n2038, DP_mult_207_n2037, DP_mult_207_n2036,
         DP_mult_207_n2035, DP_mult_207_n2034, DP_mult_207_n2033,
         DP_mult_207_n2032, DP_mult_207_n2031, DP_mult_207_n2030,
         DP_mult_207_n2029, DP_mult_207_n2028, DP_mult_207_n2027,
         DP_mult_207_n2026, DP_mult_207_n2025, DP_mult_207_n2024,
         DP_mult_207_n2023, DP_mult_207_n2022, DP_mult_207_n2021,
         DP_mult_207_n2020, DP_mult_207_n2019, DP_mult_207_n2018,
         DP_mult_207_n2017, DP_mult_207_n2016, DP_mult_207_n2015,
         DP_mult_207_n2014, DP_mult_207_n2013, DP_mult_207_n2012,
         DP_mult_207_n2011, DP_mult_207_n2010, DP_mult_207_n2009,
         DP_mult_207_n2008, DP_mult_207_n2007, DP_mult_207_n2006,
         DP_mult_207_n2005, DP_mult_207_n2004, DP_mult_207_n2003,
         DP_mult_207_n2002, DP_mult_207_n2001, DP_mult_207_n2000,
         DP_mult_207_n1999, DP_mult_207_n1998, DP_mult_207_n1997,
         DP_mult_207_n1996, DP_mult_207_n1995, DP_mult_207_n1994,
         DP_mult_207_n1993, DP_mult_207_n1992, DP_mult_207_n1991,
         DP_mult_207_n1990, DP_mult_207_n1989, DP_mult_207_n1988,
         DP_mult_207_n1987, DP_mult_207_n1986, DP_mult_207_n1985,
         DP_mult_207_n1984, DP_mult_207_n1983, DP_mult_207_n1982,
         DP_mult_207_n1981, DP_mult_207_n1980, DP_mult_207_n1979,
         DP_mult_207_n1978, DP_mult_207_n1977, DP_mult_207_n1976,
         DP_mult_207_n1975, DP_mult_207_n1974, DP_mult_207_n1973,
         DP_mult_207_n1972, DP_mult_207_n1971, DP_mult_207_n1970,
         DP_mult_207_n1969, DP_mult_207_n1968, DP_mult_207_n1967,
         DP_mult_207_n1966, DP_mult_207_n1965, DP_mult_207_n1964,
         DP_mult_207_n1963, DP_mult_207_n1962, DP_mult_207_n1961,
         DP_mult_207_n1960, DP_mult_207_n1959, DP_mult_207_n1958,
         DP_mult_207_n1957, DP_mult_207_n1956, DP_mult_207_n1955,
         DP_mult_207_n1954, DP_mult_207_n1953, DP_mult_207_n1952,
         DP_mult_207_n1951, DP_mult_207_n1950, DP_mult_207_n1949,
         DP_mult_207_n1948, DP_mult_207_n1947, DP_mult_207_n1946,
         DP_mult_207_n1945, DP_mult_207_n1944, DP_mult_207_n1943,
         DP_mult_207_n1942, DP_mult_207_n1941, DP_mult_207_n1940,
         DP_mult_207_n1939, DP_mult_207_n1938, DP_mult_207_n1937,
         DP_mult_207_n1936, DP_mult_207_n1935, DP_mult_207_n1934,
         DP_mult_207_n1933, DP_mult_207_n1932, DP_mult_207_n1931,
         DP_mult_207_n1930, DP_mult_207_n1929, DP_mult_207_n1817,
         DP_mult_207_n1816, DP_mult_207_n1815, DP_mult_207_n1814,
         DP_mult_207_n1813, DP_mult_207_n1812, DP_mult_207_n1811,
         DP_mult_207_n1810, DP_mult_207_n1809, DP_mult_207_n1808,
         DP_mult_207_n1806, DP_mult_207_n1781, DP_mult_207_n1780,
         DP_mult_207_n1779, DP_mult_207_n1778, DP_mult_207_n1777,
         DP_mult_207_n1776, DP_mult_207_n1775, DP_mult_207_n1774,
         DP_mult_207_n1773, DP_mult_207_n1772, DP_mult_207_n1771,
         DP_mult_207_n1770, DP_mult_207_n1769, DP_mult_207_n1768,
         DP_mult_207_n1767, DP_mult_207_n1766, DP_mult_207_n1765,
         DP_mult_207_n1764, DP_mult_207_n1763, DP_mult_207_n1762,
         DP_mult_207_n1761, DP_mult_207_n1760, DP_mult_207_n1759,
         DP_mult_207_n1758, DP_mult_207_n1757, DP_mult_207_n1756,
         DP_mult_207_n1755, DP_mult_207_n1754, DP_mult_207_n1753,
         DP_mult_207_n1752, DP_mult_207_n1751, DP_mult_207_n1750,
         DP_mult_207_n1749, DP_mult_207_n1748, DP_mult_207_n1747,
         DP_mult_207_n1746, DP_mult_207_n1745, DP_mult_207_n1744,
         DP_mult_207_n1743, DP_mult_207_n1742, DP_mult_207_n1741,
         DP_mult_207_n1740, DP_mult_207_n1739, DP_mult_207_n1738,
         DP_mult_207_n1737, DP_mult_207_n1736, DP_mult_207_n1735,
         DP_mult_207_n1734, DP_mult_207_n1733, DP_mult_207_n1732,
         DP_mult_207_n1731, DP_mult_207_n1730, DP_mult_207_n1729,
         DP_mult_207_n1728, DP_mult_207_n1727, DP_mult_207_n1726,
         DP_mult_207_n1725, DP_mult_207_n1724, DP_mult_207_n1723,
         DP_mult_207_n1722, DP_mult_207_n1721, DP_mult_207_n1720,
         DP_mult_207_n1719, DP_mult_207_n1718, DP_mult_207_n1717,
         DP_mult_207_n1716, DP_mult_207_n1715, DP_mult_207_n1714,
         DP_mult_207_n1713, DP_mult_207_n1712, DP_mult_207_n1711,
         DP_mult_207_n1710, DP_mult_207_n1709, DP_mult_207_n1708,
         DP_mult_207_n1707, DP_mult_207_n1706, DP_mult_207_n1705,
         DP_mult_207_n1704, DP_mult_207_n1703, DP_mult_207_n1702,
         DP_mult_207_n1701, DP_mult_207_n1700, DP_mult_207_n1699,
         DP_mult_207_n1698, DP_mult_207_n1697, DP_mult_207_n1696,
         DP_mult_207_n1695, DP_mult_207_n1694, DP_mult_207_n1693,
         DP_mult_207_n1692, DP_mult_207_n1691, DP_mult_207_n1690,
         DP_mult_207_n1689, DP_mult_207_n1688, DP_mult_207_n1687,
         DP_mult_207_n1686, DP_mult_207_n1685, DP_mult_207_n1684,
         DP_mult_207_n1683, DP_mult_207_n1682, DP_mult_207_n1681,
         DP_mult_207_n1680, DP_mult_207_n1679, DP_mult_207_n1678,
         DP_mult_207_n1677, DP_mult_207_n1676, DP_mult_207_n1675,
         DP_mult_207_n1674, DP_mult_207_n1673, DP_mult_207_n1672,
         DP_mult_207_n1671, DP_mult_207_n1670, DP_mult_207_n1669,
         DP_mult_207_n1668, DP_mult_207_n1667, DP_mult_207_n1666,
         DP_mult_207_n1665, DP_mult_207_n1664, DP_mult_207_n1663,
         DP_mult_207_n1662, DP_mult_207_n1661, DP_mult_207_n1660,
         DP_mult_207_n1659, DP_mult_207_n1658, DP_mult_207_n1657,
         DP_mult_207_n1656, DP_mult_207_n1655, DP_mult_207_n1654,
         DP_mult_207_n1653, DP_mult_207_n1652, DP_mult_207_n1651,
         DP_mult_207_n1650, DP_mult_207_n1649, DP_mult_207_n1648,
         DP_mult_207_n1647, DP_mult_207_n1646, DP_mult_207_n1645,
         DP_mult_207_n1644, DP_mult_207_n1643, DP_mult_207_n1642,
         DP_mult_207_n1641, DP_mult_207_n1640, DP_mult_207_n1639,
         DP_mult_207_n1638, DP_mult_207_n1637, DP_mult_207_n1636,
         DP_mult_207_n1635, DP_mult_207_n1634, DP_mult_207_n1633,
         DP_mult_207_n1632, DP_mult_207_n1631, DP_mult_207_n1630,
         DP_mult_207_n1629, DP_mult_207_n1628, DP_mult_207_n1627,
         DP_mult_207_n1626, DP_mult_207_n1625, DP_mult_207_n1624,
         DP_mult_207_n1623, DP_mult_207_n1622, DP_mult_207_n1621,
         DP_mult_207_n1620, DP_mult_207_n1619, DP_mult_207_n1618,
         DP_mult_207_n1617, DP_mult_207_n1616, DP_mult_207_n1615,
         DP_mult_207_n1614, DP_mult_207_n1613, DP_mult_207_n1612,
         DP_mult_207_n1611, DP_mult_207_n1610, DP_mult_207_n1609,
         DP_mult_207_n1608, DP_mult_207_n1607, DP_mult_207_n1606,
         DP_mult_207_n1605, DP_mult_207_n1604, DP_mult_207_n1603,
         DP_mult_207_n1602, DP_mult_207_n1601, DP_mult_207_n1600,
         DP_mult_207_n1599, DP_mult_207_n1598, DP_mult_207_n1597,
         DP_mult_207_n1596, DP_mult_207_n1595, DP_mult_207_n1594,
         DP_mult_207_n1593, DP_mult_207_n1592, DP_mult_207_n1591,
         DP_mult_207_n1590, DP_mult_207_n1589, DP_mult_207_n1588,
         DP_mult_207_n1587, DP_mult_207_n1586, DP_mult_207_n1585,
         DP_mult_207_n1584, DP_mult_207_n1583, DP_mult_207_n1582,
         DP_mult_207_n1581, DP_mult_207_n1580, DP_mult_207_n1579,
         DP_mult_207_n1578, DP_mult_207_n1577, DP_mult_207_n1576,
         DP_mult_207_n1575, DP_mult_207_n1574, DP_mult_207_n1573,
         DP_mult_207_n1572, DP_mult_207_n1571, DP_mult_207_n1570,
         DP_mult_207_n1569, DP_mult_207_n1568, DP_mult_207_n1567,
         DP_mult_207_n1566, DP_mult_207_n1565, DP_mult_207_n1564,
         DP_mult_207_n1563, DP_mult_207_n1562, DP_mult_207_n1561,
         DP_mult_207_n1560, DP_mult_207_n1559, DP_mult_207_n1558,
         DP_mult_207_n1557, DP_mult_207_n1556, DP_mult_207_n1555,
         DP_mult_207_n1554, DP_mult_207_n1553, DP_mult_207_n1552,
         DP_mult_207_n1551, DP_mult_207_n1550, DP_mult_207_n1549,
         DP_mult_207_n1548, DP_mult_207_n1547, DP_mult_207_n1546,
         DP_mult_207_n1545, DP_mult_207_n1544, DP_mult_207_n1543,
         DP_mult_207_n1542, DP_mult_207_n1541, DP_mult_207_n1540,
         DP_mult_207_n1539, DP_mult_207_n1538, DP_mult_207_n1537,
         DP_mult_207_n1536, DP_mult_207_n1535, DP_mult_207_n1534,
         DP_mult_207_n1533, DP_mult_207_n1532, DP_mult_207_n1531,
         DP_mult_207_n1530, DP_mult_207_n1529, DP_mult_207_n1528,
         DP_mult_207_n1527, DP_mult_207_n1526, DP_mult_207_n1525,
         DP_mult_207_n1524, DP_mult_207_n1523, DP_mult_207_n1522,
         DP_mult_207_n1521, DP_mult_207_n1520, DP_mult_207_n1519,
         DP_mult_207_n1518, DP_mult_207_n1517, DP_mult_207_n1516,
         DP_mult_207_n1515, DP_mult_207_n1514, DP_mult_207_n1513,
         DP_mult_207_n1512, DP_mult_207_n1511, DP_mult_207_n1510,
         DP_mult_207_n1509, DP_mult_207_n1508, DP_mult_207_n1507,
         DP_mult_207_n1506, DP_mult_207_n1505, DP_mult_207_n1504,
         DP_mult_207_n1503, DP_mult_207_n1502, DP_mult_207_n1501,
         DP_mult_207_n1500, DP_mult_207_n1499, DP_mult_207_n1498,
         DP_mult_207_n1497, DP_mult_207_n1496, DP_mult_207_n1495,
         DP_mult_207_n1494, DP_mult_207_n1493, DP_mult_207_n1492,
         DP_mult_207_n1491, DP_mult_207_n1490, DP_mult_207_n1489,
         DP_mult_207_n1488, DP_mult_207_n1487, DP_mult_207_n1486,
         DP_mult_207_n1485, DP_mult_207_n1484, DP_mult_207_n1483,
         DP_mult_207_n1482, DP_mult_207_n1481, DP_mult_207_n1480,
         DP_mult_207_n1479, DP_mult_207_n1478, DP_mult_207_n1477,
         DP_mult_207_n1476, DP_mult_207_n1475, DP_mult_207_n1474,
         DP_mult_207_n1473, DP_mult_207_n1472, DP_mult_207_n1471,
         DP_mult_207_n1470, DP_mult_207_n1469, DP_mult_207_n1468,
         DP_mult_207_n1467, DP_mult_207_n1466, DP_mult_207_n1465,
         DP_mult_207_n1464, DP_mult_207_n1463, DP_mult_207_n1462,
         DP_mult_207_n1461, DP_mult_207_n1460, DP_mult_207_n1459,
         DP_mult_207_n1458, DP_mult_207_n1457, DP_mult_207_n1456,
         DP_mult_207_n1455, DP_mult_207_n1454, DP_mult_207_n1453,
         DP_mult_207_n1452, DP_mult_207_n1451, DP_mult_207_n1450,
         DP_mult_207_n1449, DP_mult_207_n1448, DP_mult_207_n1447,
         DP_mult_207_n1446, DP_mult_207_n1445, DP_mult_207_n1444,
         DP_mult_207_n1443, DP_mult_207_n1442, DP_mult_207_n1441,
         DP_mult_207_n1440, DP_mult_207_n1439, DP_mult_207_n1438,
         DP_mult_207_n1437, DP_mult_207_n1436, DP_mult_207_n1435,
         DP_mult_207_n1434, DP_mult_207_n1433, DP_mult_207_n1432,
         DP_mult_207_n1431, DP_mult_207_n1430, DP_mult_207_n1429,
         DP_mult_207_n1428, DP_mult_207_n1427, DP_mult_207_n1426,
         DP_mult_207_n1425, DP_mult_207_n1424, DP_mult_207_n1423,
         DP_mult_207_n1422, DP_mult_207_n1421, DP_mult_207_n1420,
         DP_mult_207_n1419, DP_mult_207_n1418, DP_mult_207_n1417,
         DP_mult_207_n1416, DP_mult_207_n1415, DP_mult_207_n1414,
         DP_mult_207_n1413, DP_mult_207_n1412, DP_mult_207_n1411,
         DP_mult_207_n1410, DP_mult_207_n1409, DP_mult_207_n1408,
         DP_mult_207_n1407, DP_mult_207_n1406, DP_mult_207_n1405,
         DP_mult_207_n1404, DP_mult_207_n1403, DP_mult_207_n1402,
         DP_mult_207_n1401, DP_mult_207_n1400, DP_mult_207_n1399,
         DP_mult_207_n1398, DP_mult_207_n1397, DP_mult_207_n1396,
         DP_mult_207_n1395, DP_mult_207_n1394, DP_mult_207_n1393,
         DP_mult_207_n1392, DP_mult_207_n1391, DP_mult_207_n1390,
         DP_mult_207_n1389, DP_mult_207_n1388, DP_mult_207_n1387,
         DP_mult_207_n1386, DP_mult_207_n1385, DP_mult_207_n1384,
         DP_mult_207_n1383, DP_mult_207_n1382, DP_mult_207_n1381,
         DP_mult_207_n1380, DP_mult_207_n1379, DP_mult_207_n1378,
         DP_mult_207_n1377, DP_mult_207_n1376, DP_mult_207_n1375,
         DP_mult_207_n1374, DP_mult_207_n1373, DP_mult_207_n1372,
         DP_mult_207_n1371, DP_mult_207_n1370, DP_mult_207_n1369,
         DP_mult_207_n1368, DP_mult_207_n1367, DP_mult_207_n1366,
         DP_mult_207_n1365, DP_mult_207_n1364, DP_mult_207_n1363,
         DP_mult_207_n1362, DP_mult_207_n1361, DP_mult_207_n1360,
         DP_mult_207_n1359, DP_mult_207_n1358, DP_mult_207_n1357,
         DP_mult_207_n1356, DP_mult_207_n1355, DP_mult_207_n1354,
         DP_mult_207_n1353, DP_mult_207_n1352, DP_mult_207_n1351,
         DP_mult_207_n1350, DP_mult_207_n1349, DP_mult_207_n1348,
         DP_mult_207_n1347, DP_mult_207_n1346, DP_mult_207_n1345,
         DP_mult_207_n1344, DP_mult_207_n1343, DP_mult_207_n1342,
         DP_mult_207_n1341, DP_mult_207_n1340, DP_mult_207_n1339,
         DP_mult_207_n1338, DP_mult_207_n1337, DP_mult_207_n1336,
         DP_mult_207_n1335, DP_mult_207_n1334, DP_mult_207_n1333,
         DP_mult_207_n1332, DP_mult_207_n1331, DP_mult_207_n1330,
         DP_mult_207_n1329, DP_mult_207_n1328, DP_mult_207_n1327,
         DP_mult_207_n1326, DP_mult_207_n1325, DP_mult_207_n1324,
         DP_mult_207_n1323, DP_mult_207_n1322, DP_mult_207_n1321,
         DP_mult_207_n1320, DP_mult_207_n1319, DP_mult_207_n1318,
         DP_mult_207_n1317, DP_mult_207_n1316, DP_mult_207_n1315,
         DP_mult_207_n1314, DP_mult_207_n1313, DP_mult_207_n1312,
         DP_mult_207_n1311, DP_mult_207_n1310, DP_mult_207_n1309,
         DP_mult_207_n1308, DP_mult_207_n1307, DP_mult_207_n1306,
         DP_mult_207_n1305, DP_mult_207_n1304, DP_mult_207_n1303,
         DP_mult_207_n1302, DP_mult_207_n1301, DP_mult_207_n1300,
         DP_mult_207_n1299, DP_mult_207_n1298, DP_mult_207_n1297,
         DP_mult_207_n1296, DP_mult_207_n1295, DP_mult_207_n1294,
         DP_mult_207_n1293, DP_mult_207_n1292, DP_mult_207_n1291,
         DP_mult_207_n1290, DP_mult_207_n1289, DP_mult_207_n1288,
         DP_mult_207_n1287, DP_mult_207_n1286, DP_mult_207_n1285,
         DP_mult_207_n1284, DP_mult_207_n1283, DP_mult_207_n1282,
         DP_mult_207_n1281, DP_mult_207_n1280, DP_mult_207_n1279,
         DP_mult_207_n1278, DP_mult_207_n1277, DP_mult_207_n1276,
         DP_mult_207_n1275, DP_mult_207_n1274, DP_mult_207_n1273,
         DP_mult_207_n1272, DP_mult_207_n1271, DP_mult_207_n1270,
         DP_mult_207_n1269, DP_mult_207_n1268, DP_mult_207_n1267,
         DP_mult_207_n1266, DP_mult_207_n1265, DP_mult_207_n1264,
         DP_mult_207_n1263, DP_mult_207_n1262, DP_mult_207_n1261,
         DP_mult_207_n1260, DP_mult_207_n1259, DP_mult_207_n1258,
         DP_mult_207_n1257, DP_mult_207_n1256, DP_mult_207_n1255,
         DP_mult_207_n1254, DP_mult_207_n1253, DP_mult_207_n1252,
         DP_mult_207_n1251, DP_mult_207_n1250, DP_mult_207_n1249,
         DP_mult_207_n1248, DP_mult_207_n1247, DP_mult_207_n1246,
         DP_mult_207_n1245, DP_mult_207_n1244, DP_mult_207_n1243,
         DP_mult_207_n1242, DP_mult_207_n1241, DP_mult_207_n1240,
         DP_mult_207_n1239, DP_mult_207_n1238, DP_mult_207_n1237,
         DP_mult_207_n1236, DP_mult_207_n1235, DP_mult_207_n1234,
         DP_mult_207_n1233, DP_mult_207_n1232, DP_mult_207_n1231,
         DP_mult_207_n1230, DP_mult_207_n1229, DP_mult_207_n1228,
         DP_mult_207_n1227, DP_mult_207_n1226, DP_mult_207_n1225,
         DP_mult_207_n1224, DP_mult_207_n1223, DP_mult_207_n1222,
         DP_mult_207_n1221, DP_mult_207_n1220, DP_mult_207_n1219,
         DP_mult_207_n1218, DP_mult_207_n1217, DP_mult_207_n1216,
         DP_mult_207_n1215, DP_mult_207_n1214, DP_mult_207_n1213,
         DP_mult_207_n1212, DP_mult_207_n1211, DP_mult_207_n1210,
         DP_mult_207_n1209, DP_mult_207_n1208, DP_mult_207_n1207,
         DP_mult_207_n1206, DP_mult_207_n1205, DP_mult_207_n1204,
         DP_mult_207_n1203, DP_mult_207_n1202, DP_mult_207_n1201,
         DP_mult_207_n1200, DP_mult_207_n1199, DP_mult_207_n1198,
         DP_mult_207_n1197, DP_mult_207_n1196, DP_mult_207_n1195,
         DP_mult_207_n1194, DP_mult_207_n1193, DP_mult_207_n1192,
         DP_mult_207_n1191, DP_mult_207_n1190, DP_mult_207_n1189,
         DP_mult_207_n1188, DP_mult_207_n1187, DP_mult_207_n1186,
         DP_mult_207_n1185, DP_mult_207_n1184, DP_mult_207_n1183,
         DP_mult_207_n1182, DP_mult_207_n1181, DP_mult_207_n1180,
         DP_mult_207_n1179, DP_mult_207_n1178, DP_mult_207_n1177,
         DP_mult_207_n1176, DP_mult_207_n1175, DP_mult_207_n1174,
         DP_mult_207_n1173, DP_mult_207_n1172, DP_mult_207_n1171,
         DP_mult_207_n1170, DP_mult_207_n1169, DP_mult_207_n1168,
         DP_mult_207_n1167, DP_mult_207_n1166, DP_mult_207_n1165,
         DP_mult_207_n1164, DP_mult_207_n1163, DP_mult_207_n1162,
         DP_mult_207_n1161, DP_mult_207_n1160, DP_mult_207_n1159,
         DP_mult_207_n1158, DP_mult_207_n1157, DP_mult_207_n1156,
         DP_mult_207_n1155, DP_mult_207_n1154, DP_mult_207_n1153,
         DP_mult_207_n1152, DP_mult_207_n1151, DP_mult_207_n1150,
         DP_mult_207_n1149, DP_mult_207_n1148, DP_mult_207_n1147,
         DP_mult_207_n1146, DP_mult_207_n1145, DP_mult_207_n1144,
         DP_mult_207_n1143, DP_mult_207_n1142, DP_mult_207_n1141,
         DP_mult_207_n1140, DP_mult_207_n1139, DP_mult_207_n1138,
         DP_mult_207_n1137, DP_mult_207_n1136, DP_mult_207_n1135,
         DP_mult_207_n1134, DP_mult_207_n1133, DP_mult_207_n1132,
         DP_mult_207_n1131, DP_mult_207_n1130, DP_mult_207_n1129,
         DP_mult_207_n1128, DP_mult_207_n1127, DP_mult_207_n1126,
         DP_mult_207_n1125, DP_mult_207_n1124, DP_mult_207_n1123,
         DP_mult_207_n1122, DP_mult_207_n1121, DP_mult_207_n1120,
         DP_mult_207_n1119, DP_mult_207_n1118, DP_mult_207_n1117,
         DP_mult_207_n1116, DP_mult_207_n1115, DP_mult_207_n1114,
         DP_mult_207_n1113, DP_mult_207_n1112, DP_mult_207_n1111,
         DP_mult_207_n1110, DP_mult_207_n1109, DP_mult_207_n1108,
         DP_mult_207_n1107, DP_mult_207_n1106, DP_mult_207_n1105,
         DP_mult_207_n1104, DP_mult_207_n1103, DP_mult_207_n1102,
         DP_mult_207_n1101, DP_mult_207_n1100, DP_mult_207_n1099,
         DP_mult_207_n1098, DP_mult_207_n1097, DP_mult_207_n1096,
         DP_mult_207_n1095, DP_mult_207_n1094, DP_mult_207_n1093,
         DP_mult_207_n1092, DP_mult_207_n1091, DP_mult_207_n1090,
         DP_mult_207_n1089, DP_mult_207_n1088, DP_mult_207_n1087,
         DP_mult_207_n1086, DP_mult_207_n1085, DP_mult_207_n1084,
         DP_mult_207_n1083, DP_mult_207_n1082, DP_mult_207_n1081,
         DP_mult_207_n1080, DP_mult_207_n1079, DP_mult_207_n1078,
         DP_mult_207_n1077, DP_mult_207_n1076, DP_mult_207_n1075,
         DP_mult_207_n1074, DP_mult_207_n1073, DP_mult_207_n1072,
         DP_mult_207_n1071, DP_mult_207_n1070, DP_mult_207_n1069,
         DP_mult_207_n1068, DP_mult_207_n1067, DP_mult_207_n1066,
         DP_mult_207_n1065, DP_mult_207_n1064, DP_mult_207_n1063,
         DP_mult_207_n1062, DP_mult_207_n1061, DP_mult_207_n1060,
         DP_mult_207_n1059, DP_mult_207_n1058, DP_mult_207_n1057,
         DP_mult_207_n1056, DP_mult_207_n1055, DP_mult_207_n1054,
         DP_mult_207_n1053, DP_mult_207_n1052, DP_mult_207_n1051,
         DP_mult_207_n1050, DP_mult_207_n1049, DP_mult_207_n1048,
         DP_mult_207_n1047, DP_mult_207_n1046, DP_mult_207_n1045,
         DP_mult_207_n1044, DP_mult_207_n1043, DP_mult_207_n1042,
         DP_mult_207_n1041, DP_mult_207_n1040, DP_mult_207_n1039,
         DP_mult_207_n1038, DP_mult_207_n1037, DP_mult_207_n1036,
         DP_mult_207_n1035, DP_mult_207_n1034, DP_mult_207_n1033,
         DP_mult_207_n1032, DP_mult_207_n1031, DP_mult_207_n1030,
         DP_mult_207_n1029, DP_mult_207_n1028, DP_mult_207_n1027,
         DP_mult_207_n1026, DP_mult_207_n1025, DP_mult_207_n1024,
         DP_mult_207_n1023, DP_mult_207_n1022, DP_mult_207_n1021,
         DP_mult_207_n1020, DP_mult_207_n1019, DP_mult_207_n1018,
         DP_mult_207_n1017, DP_mult_207_n1016, DP_mult_207_n1015,
         DP_mult_207_n1014, DP_mult_207_n1013, DP_mult_207_n1012,
         DP_mult_207_n1011, DP_mult_207_n1010, DP_mult_207_n1009,
         DP_mult_207_n1008, DP_mult_207_n1007, DP_mult_207_n1006,
         DP_mult_207_n1005, DP_mult_207_n1004, DP_mult_207_n1003,
         DP_mult_207_n1002, DP_mult_207_n1001, DP_mult_207_n1000,
         DP_mult_207_n999, DP_mult_207_n998, DP_mult_207_n997,
         DP_mult_207_n996, DP_mult_207_n995, DP_mult_207_n994,
         DP_mult_207_n993, DP_mult_207_n992, DP_mult_207_n991,
         DP_mult_207_n990, DP_mult_207_n989, DP_mult_207_n988,
         DP_mult_207_n987, DP_mult_207_n986, DP_mult_207_n985,
         DP_mult_207_n984, DP_mult_207_n983, DP_mult_207_n982,
         DP_mult_207_n981, DP_mult_207_n980, DP_mult_207_n979,
         DP_mult_207_n978, DP_mult_207_n977, DP_mult_207_n976,
         DP_mult_207_n975, DP_mult_207_n974, DP_mult_207_n973,
         DP_mult_207_n972, DP_mult_207_n971, DP_mult_207_n970,
         DP_mult_207_n969, DP_mult_207_n968, DP_mult_207_n967,
         DP_mult_207_n966, DP_mult_207_n965, DP_mult_207_n964,
         DP_mult_207_n963, DP_mult_207_n962, DP_mult_207_n961,
         DP_mult_207_n960, DP_mult_207_n959, DP_mult_207_n958,
         DP_mult_207_n957, DP_mult_207_n956, DP_mult_207_n955,
         DP_mult_207_n954, DP_mult_207_n953, DP_mult_207_n952,
         DP_mult_207_n951, DP_mult_207_n950, DP_mult_207_n949,
         DP_mult_207_n948, DP_mult_207_n947, DP_mult_207_n946,
         DP_mult_207_n945, DP_mult_207_n944, DP_mult_207_n943,
         DP_mult_207_n942, DP_mult_207_n941, DP_mult_207_n940,
         DP_mult_207_n939, DP_mult_207_n938, DP_mult_207_n937,
         DP_mult_207_n936, DP_mult_207_n935, DP_mult_207_n934,
         DP_mult_207_n933, DP_mult_207_n932, DP_mult_207_n931,
         DP_mult_207_n930, DP_mult_207_n929, DP_mult_207_n928,
         DP_mult_207_n927, DP_mult_207_n926, DP_mult_207_n925,
         DP_mult_207_n924, DP_mult_207_n923, DP_mult_207_n922,
         DP_mult_207_n921, DP_mult_207_n920, DP_mult_207_n918,
         DP_mult_207_n917, DP_mult_207_n916, DP_mult_207_n915,
         DP_mult_207_n914, DP_mult_207_n913, DP_mult_207_n912,
         DP_mult_207_n911, DP_mult_207_n910, DP_mult_207_n909,
         DP_mult_207_n908, DP_mult_207_n907, DP_mult_207_n906,
         DP_mult_207_n905, DP_mult_207_n904, DP_mult_207_n903,
         DP_mult_207_n902, DP_mult_207_n901, DP_mult_207_n900,
         DP_mult_207_n899, DP_mult_207_n898, DP_mult_207_n897,
         DP_mult_207_n896, DP_mult_207_n895, DP_mult_207_n894,
         DP_mult_207_n893, DP_mult_207_n892, DP_mult_207_n891,
         DP_mult_207_n890, DP_mult_207_n889, DP_mult_207_n888,
         DP_mult_207_n887, DP_mult_207_n886, DP_mult_207_n885,
         DP_mult_207_n884, DP_mult_207_n883, DP_mult_207_n882,
         DP_mult_207_n881, DP_mult_207_n880, DP_mult_207_n879,
         DP_mult_207_n878, DP_mult_207_n877, DP_mult_207_n876,
         DP_mult_207_n875, DP_mult_207_n874, DP_mult_207_n873,
         DP_mult_207_n872, DP_mult_207_n871, DP_mult_207_n870,
         DP_mult_207_n869, DP_mult_207_n868, DP_mult_207_n867,
         DP_mult_207_n866, DP_mult_207_n865, DP_mult_207_n864,
         DP_mult_207_n863, DP_mult_207_n862, DP_mult_207_n861,
         DP_mult_207_n860, DP_mult_207_n859, DP_mult_207_n858,
         DP_mult_207_n857, DP_mult_207_n856, DP_mult_207_n855,
         DP_mult_207_n854, DP_mult_207_n853, DP_mult_207_n852,
         DP_mult_207_n851, DP_mult_207_n850, DP_mult_207_n849,
         DP_mult_207_n848, DP_mult_207_n847, DP_mult_207_n846,
         DP_mult_207_n845, DP_mult_207_n844, DP_mult_207_n843,
         DP_mult_207_n842, DP_mult_207_n841, DP_mult_207_n840,
         DP_mult_207_n839, DP_mult_207_n838, DP_mult_207_n837,
         DP_mult_207_n836, DP_mult_207_n835, DP_mult_207_n834,
         DP_mult_207_n833, DP_mult_207_n832, DP_mult_207_n831,
         DP_mult_207_n830, DP_mult_207_n829, DP_mult_207_n828,
         DP_mult_207_n827, DP_mult_207_n826, DP_mult_207_n825,
         DP_mult_207_n824, DP_mult_207_n823, DP_mult_207_n822,
         DP_mult_207_n821, DP_mult_207_n820, DP_mult_207_n819,
         DP_mult_207_n818, DP_mult_207_n817, DP_mult_207_n816,
         DP_mult_207_n815, DP_mult_207_n814, DP_mult_207_n813,
         DP_mult_207_n812, DP_mult_207_n811, DP_mult_207_n810,
         DP_mult_207_n809, DP_mult_207_n808, DP_mult_207_n807,
         DP_mult_207_n806, DP_mult_207_n805, DP_mult_207_n804,
         DP_mult_207_n803, DP_mult_207_n802, DP_mult_207_n801,
         DP_mult_207_n800, DP_mult_207_n799, DP_mult_207_n798,
         DP_mult_207_n797, DP_mult_207_n796, DP_mult_207_n795,
         DP_mult_207_n794, DP_mult_207_n793, DP_mult_207_n792,
         DP_mult_207_n791, DP_mult_207_n790, DP_mult_207_n789,
         DP_mult_207_n788, DP_mult_207_n787, DP_mult_207_n786,
         DP_mult_207_n785, DP_mult_207_n784, DP_mult_207_n783,
         DP_mult_207_n782, DP_mult_207_n781, DP_mult_207_n780,
         DP_mult_207_n779, DP_mult_207_n778, DP_mult_207_n777,
         DP_mult_207_n776, DP_mult_207_n775, DP_mult_207_n774,
         DP_mult_207_n773, DP_mult_207_n772, DP_mult_207_n771,
         DP_mult_207_n770, DP_mult_207_n769, DP_mult_207_n768,
         DP_mult_207_n767, DP_mult_207_n766, DP_mult_207_n765,
         DP_mult_207_n764, DP_mult_207_n763, DP_mult_207_n762,
         DP_mult_207_n761, DP_mult_207_n760, DP_mult_207_n759,
         DP_mult_207_n758, DP_mult_207_n757, DP_mult_207_n756,
         DP_mult_207_n755, DP_mult_207_n754, DP_mult_207_n753,
         DP_mult_207_n752, DP_mult_207_n751, DP_mult_207_n750,
         DP_mult_207_n749, DP_mult_207_n748, DP_mult_207_n747,
         DP_mult_207_n746, DP_mult_207_n745, DP_mult_207_n744,
         DP_mult_207_n743, DP_mult_207_n742, DP_mult_207_n741,
         DP_mult_207_n740, DP_mult_207_n739, DP_mult_207_n738,
         DP_mult_207_n737, DP_mult_207_n736, DP_mult_207_n735,
         DP_mult_207_n734, DP_mult_207_n733, DP_mult_207_n732,
         DP_mult_207_n731, DP_mult_207_n730, DP_mult_207_n729,
         DP_mult_207_n728, DP_mult_207_n727, DP_mult_207_n726,
         DP_mult_207_n725, DP_mult_207_n724, DP_mult_207_n723,
         DP_mult_207_n722, DP_mult_207_n721, DP_mult_207_n720,
         DP_mult_207_n719, DP_mult_207_n718, DP_mult_207_n717,
         DP_mult_207_n716, DP_mult_207_n715, DP_mult_207_n714,
         DP_mult_207_n713, DP_mult_207_n712, DP_mult_207_n711,
         DP_mult_207_n710, DP_mult_207_n709, DP_mult_207_n708,
         DP_mult_207_n707, DP_mult_207_n706, DP_mult_207_n705,
         DP_mult_207_n704, DP_mult_207_n703, DP_mult_207_n702,
         DP_mult_207_n701, DP_mult_207_n700, DP_mult_207_n699,
         DP_mult_207_n698, DP_mult_207_n697, DP_mult_207_n696,
         DP_mult_207_n695, DP_mult_207_n694, DP_mult_207_n693,
         DP_mult_207_n692, DP_mult_207_n691, DP_mult_207_n690,
         DP_mult_207_n689, DP_mult_207_n688, DP_mult_207_n687,
         DP_mult_207_n686, DP_mult_207_n685, DP_mult_207_n684,
         DP_mult_207_n683, DP_mult_207_n682, DP_mult_207_n681,
         DP_mult_207_n680, DP_mult_207_n679, DP_mult_207_n678,
         DP_mult_207_n677, DP_mult_207_n676, DP_mult_207_n672,
         DP_mult_207_n670, DP_mult_207_n668, DP_mult_207_n666,
         DP_mult_207_n663, DP_mult_207_n662, DP_mult_207_n661,
         DP_mult_207_n657, DP_mult_207_n646, DP_mult_207_n645,
         DP_mult_207_n644, DP_mult_207_n643, DP_mult_207_n638,
         DP_mult_207_n637, DP_mult_207_n636, DP_mult_207_n635,
         DP_mult_207_n634, DP_mult_207_n633, DP_mult_207_n632,
         DP_mult_207_n631, DP_mult_207_n630, DP_mult_207_n629,
         DP_mult_207_n628, DP_mult_207_n627, DP_mult_207_n626,
         DP_mult_207_n625, DP_mult_207_n620, DP_mult_207_n611,
         DP_mult_207_n610, DP_mult_207_n609, DP_mult_207_n600,
         DP_mult_207_n599, DP_mult_207_n598, DP_mult_207_n597,
         DP_mult_207_n596, DP_mult_207_n595, DP_mult_207_n594,
         DP_mult_207_n593, DP_mult_207_n592, DP_mult_207_n591,
         DP_mult_207_n590, DP_mult_207_n589, DP_mult_207_n588,
         DP_mult_207_n583, DP_mult_207_n582, DP_mult_207_n581,
         DP_mult_207_n572, DP_mult_207_n571, DP_mult_207_n570,
         DP_mult_207_n569, DP_mult_207_n568, DP_mult_207_n567,
         DP_mult_207_n566, DP_mult_207_n565, DP_mult_207_n564,
         DP_mult_207_n563, DP_mult_207_n562, DP_mult_207_n561,
         DP_mult_207_n560, DP_mult_207_n559, DP_mult_207_n558,
         DP_mult_207_n555, DP_mult_207_n553, DP_mult_207_n552,
         DP_mult_207_n551, DP_mult_207_n550, DP_mult_207_n547,
         DP_mult_207_n546, DP_mult_207_n545, DP_mult_207_n544,
         DP_mult_207_n543, DP_mult_207_n542, DP_mult_207_n541,
         DP_mult_207_n540, DP_mult_207_n539, DP_mult_207_n538,
         DP_mult_207_n537, DP_mult_207_n536, DP_mult_207_n535,
         DP_mult_207_n534, DP_mult_207_n533, DP_mult_207_n532,
         DP_mult_207_n531, DP_mult_207_n526, DP_mult_207_n525,
         DP_mult_207_n524, DP_mult_207_n523, DP_mult_207_n522,
         DP_mult_207_n521, DP_mult_207_n520, DP_mult_207_n519,
         DP_mult_207_n517, DP_mult_207_n516, DP_mult_207_n515,
         DP_mult_207_n514, DP_mult_207_n513, DP_mult_207_n512,
         DP_mult_207_n511, DP_mult_207_n508, DP_mult_207_n505,
         DP_mult_207_n504, DP_mult_207_n503, DP_mult_207_n502,
         DP_mult_207_n501, DP_mult_207_n499, DP_mult_207_n498,
         DP_mult_207_n497, DP_mult_207_n496, DP_mult_207_n495,
         DP_mult_207_n492, DP_mult_207_n491, DP_mult_207_n490,
         DP_mult_207_n488, DP_mult_207_n487, DP_mult_207_n486,
         DP_mult_207_n483, DP_mult_207_n481, DP_mult_207_n480,
         DP_mult_207_n479, DP_mult_207_n478, DP_mult_207_n477,
         DP_mult_207_n476, DP_mult_207_n475, DP_mult_207_n474,
         DP_mult_207_n472, DP_mult_207_n468, DP_mult_207_n467,
         DP_mult_207_n466, DP_mult_207_n465, DP_mult_207_n464,
         DP_mult_207_n463, DP_mult_207_n462, DP_mult_207_n461,
         DP_mult_207_n459, DP_mult_207_n457, DP_mult_207_n456,
         DP_mult_207_n455, DP_mult_207_n454, DP_mult_207_n453,
         DP_mult_207_n452, DP_mult_207_n451, DP_mult_207_n450,
         DP_mult_207_n445, DP_mult_207_n439, DP_mult_207_n438,
         DP_mult_207_n437, DP_mult_207_n436, DP_mult_207_n435,
         DP_mult_207_n434, DP_mult_207_n432, DP_mult_207_n431,
         DP_mult_207_n430, DP_mult_207_n429, DP_mult_207_n428,
         DP_mult_207_n427, DP_mult_207_n426, DP_mult_207_n423,
         DP_mult_207_n422, DP_mult_207_n421, DP_mult_207_n420,
         DP_mult_207_n419, DP_mult_207_n418, DP_mult_207_n416,
         DP_mult_207_n412, DP_mult_207_n411, DP_mult_207_n410,
         DP_mult_207_n409, DP_mult_207_n407, DP_mult_207_n405,
         DP_mult_207_n402, DP_mult_207_n401, DP_mult_207_n400,
         DP_mult_207_n399, DP_mult_207_n398, DP_mult_207_n397,
         DP_mult_207_n396, DP_mult_207_n394, DP_mult_207_n390,
         DP_mult_207_n389, DP_mult_207_n388, DP_mult_207_n387,
         DP_mult_207_n384, DP_mult_207_n383, DP_mult_207_n382,
         DP_mult_207_n381, DP_mult_207_n380, DP_mult_207_n379,
         DP_mult_207_n378, DP_mult_207_n376, DP_mult_207_n372,
         DP_mult_207_n371, DP_mult_207_n370, DP_mult_207_n369,
         DP_mult_207_n367, DP_mult_207_n365, DP_mult_207_n364,
         DP_mult_207_n363, DP_mult_207_n362, DP_mult_207_n361,
         DP_mult_207_n360, DP_mult_207_n359, DP_mult_207_n356,
         DP_mult_207_n355, DP_mult_207_n354, DP_mult_207_n353,
         DP_mult_207_n352, DP_mult_207_n350, DP_mult_207_n348,
         DP_mult_207_n347, DP_mult_207_n346, DP_mult_207_n345,
         DP_mult_207_n344, DP_mult_207_n343, DP_mult_207_n342,
         DP_mult_207_n341, DP_mult_207_n339, DP_mult_207_n337,
         DP_mult_207_n336, DP_mult_207_n335, DP_mult_207_n334,
         DP_mult_207_n333, DP_mult_207_n332, DP_mult_207_n327,
         DP_mult_207_n326, DP_mult_207_n325, DP_mult_207_n320,
         DP_mult_207_n319, DP_mult_207_n318, DP_mult_207_n317,
         DP_mult_207_n316, DP_mult_207_n315, DP_mult_207_n314,
         DP_mult_207_n313, DP_mult_207_n311, DP_mult_207_n310,
         DP_mult_207_n309, DP_mult_207_n308, DP_mult_207_n307,
         DP_mult_207_n306, DP_mult_207_n305, DP_mult_207_n304,
         DP_mult_207_n303, DP_mult_207_n302, DP_mult_207_n301,
         DP_mult_207_n265, DP_mult_207_n259, DP_mult_207_n251,
         DP_mult_208_n2282, DP_mult_208_n2281, DP_mult_208_n2280,
         DP_mult_208_n2279, DP_mult_208_n2278, DP_mult_208_n2277,
         DP_mult_208_n2276, DP_mult_208_n2275, DP_mult_208_n2274,
         DP_mult_208_n2273, DP_mult_208_n2272, DP_mult_208_n2271,
         DP_mult_208_n2270, DP_mult_208_n2269, DP_mult_208_n2268,
         DP_mult_208_n2267, DP_mult_208_n2266, DP_mult_208_n2265,
         DP_mult_208_n2264, DP_mult_208_n2263, DP_mult_208_n2262,
         DP_mult_208_n2261, DP_mult_208_n2260, DP_mult_208_n2259,
         DP_mult_208_n2258, DP_mult_208_n2257, DP_mult_208_n2256,
         DP_mult_208_n2255, DP_mult_208_n2254, DP_mult_208_n2253,
         DP_mult_208_n2252, DP_mult_208_n2251, DP_mult_208_n2250,
         DP_mult_208_n2249, DP_mult_208_n2248, DP_mult_208_n2247,
         DP_mult_208_n2246, DP_mult_208_n2245, DP_mult_208_n2244,
         DP_mult_208_n2243, DP_mult_208_n2242, DP_mult_208_n2241,
         DP_mult_208_n2240, DP_mult_208_n2239, DP_mult_208_n2238,
         DP_mult_208_n2237, DP_mult_208_n2236, DP_mult_208_n2235,
         DP_mult_208_n2234, DP_mult_208_n2233, DP_mult_208_n2232,
         DP_mult_208_n2231, DP_mult_208_n2230, DP_mult_208_n2229,
         DP_mult_208_n2228, DP_mult_208_n2227, DP_mult_208_n2226,
         DP_mult_208_n2225, DP_mult_208_n2224, DP_mult_208_n2223,
         DP_mult_208_n2222, DP_mult_208_n2221, DP_mult_208_n2220,
         DP_mult_208_n2219, DP_mult_208_n2218, DP_mult_208_n2217,
         DP_mult_208_n2216, DP_mult_208_n2215, DP_mult_208_n2214,
         DP_mult_208_n2213, DP_mult_208_n2212, DP_mult_208_n2211,
         DP_mult_208_n2210, DP_mult_208_n2209, DP_mult_208_n2208,
         DP_mult_208_n2207, DP_mult_208_n2206, DP_mult_208_n2205,
         DP_mult_208_n2204, DP_mult_208_n2203, DP_mult_208_n2202,
         DP_mult_208_n2201, DP_mult_208_n2200, DP_mult_208_n2199,
         DP_mult_208_n2198, DP_mult_208_n2197, DP_mult_208_n2196,
         DP_mult_208_n2195, DP_mult_208_n2194, DP_mult_208_n2193,
         DP_mult_208_n2192, DP_mult_208_n2191, DP_mult_208_n2190,
         DP_mult_208_n2189, DP_mult_208_n2188, DP_mult_208_n2187,
         DP_mult_208_n2186, DP_mult_208_n2185, DP_mult_208_n2184,
         DP_mult_208_n2183, DP_mult_208_n2182, DP_mult_208_n2181,
         DP_mult_208_n2180, DP_mult_208_n2179, DP_mult_208_n2178,
         DP_mult_208_n2177, DP_mult_208_n2176, DP_mult_208_n2175,
         DP_mult_208_n2174, DP_mult_208_n2173, DP_mult_208_n2172,
         DP_mult_208_n2171, DP_mult_208_n2170, DP_mult_208_n2169,
         DP_mult_208_n2168, DP_mult_208_n2167, DP_mult_208_n2166,
         DP_mult_208_n2165, DP_mult_208_n2164, DP_mult_208_n2163,
         DP_mult_208_n2162, DP_mult_208_n2161, DP_mult_208_n2160,
         DP_mult_208_n2159, DP_mult_208_n2158, DP_mult_208_n2157,
         DP_mult_208_n2156, DP_mult_208_n2155, DP_mult_208_n2154,
         DP_mult_208_n2153, DP_mult_208_n2152, DP_mult_208_n2151,
         DP_mult_208_n2150, DP_mult_208_n2149, DP_mult_208_n2148,
         DP_mult_208_n2147, DP_mult_208_n2146, DP_mult_208_n2145,
         DP_mult_208_n2144, DP_mult_208_n2143, DP_mult_208_n2142,
         DP_mult_208_n2141, DP_mult_208_n2140, DP_mult_208_n2139,
         DP_mult_208_n2138, DP_mult_208_n2137, DP_mult_208_n2136,
         DP_mult_208_n2135, DP_mult_208_n2134, DP_mult_208_n2133,
         DP_mult_208_n2132, DP_mult_208_n2131, DP_mult_208_n2130,
         DP_mult_208_n2129, DP_mult_208_n2128, DP_mult_208_n2127,
         DP_mult_208_n2126, DP_mult_208_n2125, DP_mult_208_n2124,
         DP_mult_208_n2123, DP_mult_208_n2122, DP_mult_208_n2121,
         DP_mult_208_n2120, DP_mult_208_n2119, DP_mult_208_n2118,
         DP_mult_208_n2117, DP_mult_208_n2116, DP_mult_208_n2115,
         DP_mult_208_n2114, DP_mult_208_n2113, DP_mult_208_n2112,
         DP_mult_208_n2111, DP_mult_208_n2110, DP_mult_208_n2109,
         DP_mult_208_n2108, DP_mult_208_n2107, DP_mult_208_n2106,
         DP_mult_208_n2105, DP_mult_208_n2104, DP_mult_208_n2103,
         DP_mult_208_n2102, DP_mult_208_n2101, DP_mult_208_n2100,
         DP_mult_208_n2099, DP_mult_208_n2098, DP_mult_208_n2097,
         DP_mult_208_n2096, DP_mult_208_n2095, DP_mult_208_n2094,
         DP_mult_208_n2093, DP_mult_208_n2092, DP_mult_208_n2091,
         DP_mult_208_n2090, DP_mult_208_n2089, DP_mult_208_n2088,
         DP_mult_208_n2087, DP_mult_208_n2086, DP_mult_208_n2085,
         DP_mult_208_n2084, DP_mult_208_n2083, DP_mult_208_n2082,
         DP_mult_208_n2081, DP_mult_208_n2080, DP_mult_208_n2079,
         DP_mult_208_n2078, DP_mult_208_n2077, DP_mult_208_n2076,
         DP_mult_208_n2075, DP_mult_208_n2074, DP_mult_208_n2073,
         DP_mult_208_n2072, DP_mult_208_n2071, DP_mult_208_n2070,
         DP_mult_208_n2069, DP_mult_208_n2068, DP_mult_208_n2067,
         DP_mult_208_n2066, DP_mult_208_n2065, DP_mult_208_n2064,
         DP_mult_208_n2063, DP_mult_208_n2062, DP_mult_208_n2061,
         DP_mult_208_n2060, DP_mult_208_n2059, DP_mult_208_n2058,
         DP_mult_208_n2057, DP_mult_208_n2056, DP_mult_208_n2055,
         DP_mult_208_n2054, DP_mult_208_n2053, DP_mult_208_n2052,
         DP_mult_208_n2051, DP_mult_208_n2050, DP_mult_208_n2049,
         DP_mult_208_n2048, DP_mult_208_n2047, DP_mult_208_n2046,
         DP_mult_208_n2045, DP_mult_208_n2044, DP_mult_208_n2043,
         DP_mult_208_n2042, DP_mult_208_n2041, DP_mult_208_n2040,
         DP_mult_208_n2039, DP_mult_208_n2038, DP_mult_208_n2037,
         DP_mult_208_n2036, DP_mult_208_n2035, DP_mult_208_n2034,
         DP_mult_208_n2033, DP_mult_208_n2032, DP_mult_208_n2031,
         DP_mult_208_n2030, DP_mult_208_n2029, DP_mult_208_n2028,
         DP_mult_208_n2027, DP_mult_208_n2026, DP_mult_208_n2025,
         DP_mult_208_n2024, DP_mult_208_n2023, DP_mult_208_n2022,
         DP_mult_208_n2021, DP_mult_208_n2020, DP_mult_208_n2019,
         DP_mult_208_n2018, DP_mult_208_n2017, DP_mult_208_n2016,
         DP_mult_208_n2015, DP_mult_208_n2014, DP_mult_208_n2013,
         DP_mult_208_n2012, DP_mult_208_n2011, DP_mult_208_n2010,
         DP_mult_208_n2009, DP_mult_208_n2008, DP_mult_208_n2007,
         DP_mult_208_n2006, DP_mult_208_n2005, DP_mult_208_n2004,
         DP_mult_208_n2003, DP_mult_208_n2002, DP_mult_208_n2001,
         DP_mult_208_n2000, DP_mult_208_n1999, DP_mult_208_n1998,
         DP_mult_208_n1997, DP_mult_208_n1996, DP_mult_208_n1995,
         DP_mult_208_n1994, DP_mult_208_n1993, DP_mult_208_n1992,
         DP_mult_208_n1991, DP_mult_208_n1990, DP_mult_208_n1989,
         DP_mult_208_n1988, DP_mult_208_n1987, DP_mult_208_n1986,
         DP_mult_208_n1985, DP_mult_208_n1984, DP_mult_208_n1983,
         DP_mult_208_n1982, DP_mult_208_n1981, DP_mult_208_n1980,
         DP_mult_208_n1979, DP_mult_208_n1978, DP_mult_208_n1977,
         DP_mult_208_n1976, DP_mult_208_n1975, DP_mult_208_n1974,
         DP_mult_208_n1973, DP_mult_208_n1972, DP_mult_208_n1971,
         DP_mult_208_n1970, DP_mult_208_n1969, DP_mult_208_n1968,
         DP_mult_208_n1967, DP_mult_208_n1966, DP_mult_208_n1965,
         DP_mult_208_n1964, DP_mult_208_n1963, DP_mult_208_n1962,
         DP_mult_208_n1961, DP_mult_208_n1960, DP_mult_208_n1959,
         DP_mult_208_n1958, DP_mult_208_n1957, DP_mult_208_n1956,
         DP_mult_208_n1955, DP_mult_208_n1954, DP_mult_208_n1953,
         DP_mult_208_n1952, DP_mult_208_n1951, DP_mult_208_n1950,
         DP_mult_208_n1949, DP_mult_208_n1948, DP_mult_208_n1947,
         DP_mult_208_n1946, DP_mult_208_n1945, DP_mult_208_n1944,
         DP_mult_208_n1943, DP_mult_208_n1942, DP_mult_208_n1941,
         DP_mult_208_n1940, DP_mult_208_n1939, DP_mult_208_n1938,
         DP_mult_208_n1937, DP_mult_208_n1936, DP_mult_208_n1935,
         DP_mult_208_n1934, DP_mult_208_n1933, DP_mult_208_n1932,
         DP_mult_208_n1931, DP_mult_208_n1930, DP_mult_208_n1929,
         DP_mult_208_n1817, DP_mult_208_n1816, DP_mult_208_n1815,
         DP_mult_208_n1814, DP_mult_208_n1813, DP_mult_208_n1811,
         DP_mult_208_n1810, DP_mult_208_n1809, DP_mult_208_n1808,
         DP_mult_208_n1807, DP_mult_208_n1806, DP_mult_208_n1781,
         DP_mult_208_n1780, DP_mult_208_n1779, DP_mult_208_n1778,
         DP_mult_208_n1777, DP_mult_208_n1776, DP_mult_208_n1775,
         DP_mult_208_n1774, DP_mult_208_n1773, DP_mult_208_n1772,
         DP_mult_208_n1771, DP_mult_208_n1770, DP_mult_208_n1769,
         DP_mult_208_n1768, DP_mult_208_n1767, DP_mult_208_n1766,
         DP_mult_208_n1765, DP_mult_208_n1764, DP_mult_208_n1763,
         DP_mult_208_n1762, DP_mult_208_n1761, DP_mult_208_n1760,
         DP_mult_208_n1759, DP_mult_208_n1758, DP_mult_208_n1757,
         DP_mult_208_n1756, DP_mult_208_n1755, DP_mult_208_n1754,
         DP_mult_208_n1753, DP_mult_208_n1752, DP_mult_208_n1751,
         DP_mult_208_n1750, DP_mult_208_n1749, DP_mult_208_n1748,
         DP_mult_208_n1747, DP_mult_208_n1746, DP_mult_208_n1745,
         DP_mult_208_n1744, DP_mult_208_n1743, DP_mult_208_n1742,
         DP_mult_208_n1741, DP_mult_208_n1740, DP_mult_208_n1739,
         DP_mult_208_n1738, DP_mult_208_n1737, DP_mult_208_n1736,
         DP_mult_208_n1735, DP_mult_208_n1734, DP_mult_208_n1733,
         DP_mult_208_n1732, DP_mult_208_n1731, DP_mult_208_n1730,
         DP_mult_208_n1729, DP_mult_208_n1728, DP_mult_208_n1727,
         DP_mult_208_n1726, DP_mult_208_n1725, DP_mult_208_n1724,
         DP_mult_208_n1723, DP_mult_208_n1722, DP_mult_208_n1721,
         DP_mult_208_n1720, DP_mult_208_n1719, DP_mult_208_n1718,
         DP_mult_208_n1717, DP_mult_208_n1716, DP_mult_208_n1715,
         DP_mult_208_n1714, DP_mult_208_n1713, DP_mult_208_n1712,
         DP_mult_208_n1711, DP_mult_208_n1710, DP_mult_208_n1709,
         DP_mult_208_n1708, DP_mult_208_n1707, DP_mult_208_n1706,
         DP_mult_208_n1705, DP_mult_208_n1704, DP_mult_208_n1703,
         DP_mult_208_n1702, DP_mult_208_n1701, DP_mult_208_n1700,
         DP_mult_208_n1699, DP_mult_208_n1698, DP_mult_208_n1697,
         DP_mult_208_n1696, DP_mult_208_n1695, DP_mult_208_n1694,
         DP_mult_208_n1693, DP_mult_208_n1692, DP_mult_208_n1691,
         DP_mult_208_n1690, DP_mult_208_n1689, DP_mult_208_n1688,
         DP_mult_208_n1687, DP_mult_208_n1686, DP_mult_208_n1685,
         DP_mult_208_n1684, DP_mult_208_n1683, DP_mult_208_n1682,
         DP_mult_208_n1681, DP_mult_208_n1680, DP_mult_208_n1679,
         DP_mult_208_n1678, DP_mult_208_n1677, DP_mult_208_n1676,
         DP_mult_208_n1675, DP_mult_208_n1674, DP_mult_208_n1673,
         DP_mult_208_n1672, DP_mult_208_n1671, DP_mult_208_n1670,
         DP_mult_208_n1669, DP_mult_208_n1668, DP_mult_208_n1667,
         DP_mult_208_n1666, DP_mult_208_n1665, DP_mult_208_n1664,
         DP_mult_208_n1663, DP_mult_208_n1662, DP_mult_208_n1661,
         DP_mult_208_n1660, DP_mult_208_n1659, DP_mult_208_n1658,
         DP_mult_208_n1657, DP_mult_208_n1656, DP_mult_208_n1655,
         DP_mult_208_n1654, DP_mult_208_n1653, DP_mult_208_n1652,
         DP_mult_208_n1651, DP_mult_208_n1650, DP_mult_208_n1649,
         DP_mult_208_n1648, DP_mult_208_n1647, DP_mult_208_n1646,
         DP_mult_208_n1645, DP_mult_208_n1644, DP_mult_208_n1643,
         DP_mult_208_n1642, DP_mult_208_n1641, DP_mult_208_n1640,
         DP_mult_208_n1639, DP_mult_208_n1638, DP_mult_208_n1637,
         DP_mult_208_n1636, DP_mult_208_n1635, DP_mult_208_n1634,
         DP_mult_208_n1633, DP_mult_208_n1632, DP_mult_208_n1631,
         DP_mult_208_n1630, DP_mult_208_n1629, DP_mult_208_n1628,
         DP_mult_208_n1627, DP_mult_208_n1626, DP_mult_208_n1625,
         DP_mult_208_n1624, DP_mult_208_n1623, DP_mult_208_n1622,
         DP_mult_208_n1621, DP_mult_208_n1620, DP_mult_208_n1619,
         DP_mult_208_n1618, DP_mult_208_n1617, DP_mult_208_n1616,
         DP_mult_208_n1615, DP_mult_208_n1614, DP_mult_208_n1613,
         DP_mult_208_n1612, DP_mult_208_n1611, DP_mult_208_n1610,
         DP_mult_208_n1609, DP_mult_208_n1608, DP_mult_208_n1607,
         DP_mult_208_n1606, DP_mult_208_n1605, DP_mult_208_n1604,
         DP_mult_208_n1603, DP_mult_208_n1602, DP_mult_208_n1601,
         DP_mult_208_n1600, DP_mult_208_n1599, DP_mult_208_n1598,
         DP_mult_208_n1597, DP_mult_208_n1596, DP_mult_208_n1595,
         DP_mult_208_n1594, DP_mult_208_n1593, DP_mult_208_n1592,
         DP_mult_208_n1591, DP_mult_208_n1590, DP_mult_208_n1589,
         DP_mult_208_n1588, DP_mult_208_n1587, DP_mult_208_n1586,
         DP_mult_208_n1585, DP_mult_208_n1584, DP_mult_208_n1583,
         DP_mult_208_n1582, DP_mult_208_n1581, DP_mult_208_n1580,
         DP_mult_208_n1579, DP_mult_208_n1578, DP_mult_208_n1577,
         DP_mult_208_n1576, DP_mult_208_n1575, DP_mult_208_n1574,
         DP_mult_208_n1573, DP_mult_208_n1572, DP_mult_208_n1571,
         DP_mult_208_n1570, DP_mult_208_n1569, DP_mult_208_n1568,
         DP_mult_208_n1567, DP_mult_208_n1566, DP_mult_208_n1565,
         DP_mult_208_n1564, DP_mult_208_n1563, DP_mult_208_n1562,
         DP_mult_208_n1561, DP_mult_208_n1560, DP_mult_208_n1559,
         DP_mult_208_n1558, DP_mult_208_n1557, DP_mult_208_n1556,
         DP_mult_208_n1555, DP_mult_208_n1554, DP_mult_208_n1553,
         DP_mult_208_n1552, DP_mult_208_n1551, DP_mult_208_n1550,
         DP_mult_208_n1549, DP_mult_208_n1548, DP_mult_208_n1547,
         DP_mult_208_n1546, DP_mult_208_n1545, DP_mult_208_n1544,
         DP_mult_208_n1543, DP_mult_208_n1542, DP_mult_208_n1541,
         DP_mult_208_n1540, DP_mult_208_n1539, DP_mult_208_n1538,
         DP_mult_208_n1537, DP_mult_208_n1536, DP_mult_208_n1535,
         DP_mult_208_n1534, DP_mult_208_n1533, DP_mult_208_n1532,
         DP_mult_208_n1531, DP_mult_208_n1530, DP_mult_208_n1529,
         DP_mult_208_n1528, DP_mult_208_n1527, DP_mult_208_n1526,
         DP_mult_208_n1525, DP_mult_208_n1524, DP_mult_208_n1523,
         DP_mult_208_n1522, DP_mult_208_n1521, DP_mult_208_n1520,
         DP_mult_208_n1519, DP_mult_208_n1518, DP_mult_208_n1517,
         DP_mult_208_n1516, DP_mult_208_n1515, DP_mult_208_n1514,
         DP_mult_208_n1513, DP_mult_208_n1512, DP_mult_208_n1511,
         DP_mult_208_n1510, DP_mult_208_n1509, DP_mult_208_n1508,
         DP_mult_208_n1507, DP_mult_208_n1506, DP_mult_208_n1505,
         DP_mult_208_n1504, DP_mult_208_n1503, DP_mult_208_n1502,
         DP_mult_208_n1501, DP_mult_208_n1500, DP_mult_208_n1499,
         DP_mult_208_n1498, DP_mult_208_n1497, DP_mult_208_n1496,
         DP_mult_208_n1495, DP_mult_208_n1494, DP_mult_208_n1493,
         DP_mult_208_n1492, DP_mult_208_n1491, DP_mult_208_n1490,
         DP_mult_208_n1489, DP_mult_208_n1488, DP_mult_208_n1487,
         DP_mult_208_n1486, DP_mult_208_n1485, DP_mult_208_n1484,
         DP_mult_208_n1483, DP_mult_208_n1482, DP_mult_208_n1481,
         DP_mult_208_n1480, DP_mult_208_n1479, DP_mult_208_n1478,
         DP_mult_208_n1477, DP_mult_208_n1476, DP_mult_208_n1475,
         DP_mult_208_n1474, DP_mult_208_n1473, DP_mult_208_n1472,
         DP_mult_208_n1471, DP_mult_208_n1470, DP_mult_208_n1469,
         DP_mult_208_n1468, DP_mult_208_n1467, DP_mult_208_n1466,
         DP_mult_208_n1465, DP_mult_208_n1464, DP_mult_208_n1463,
         DP_mult_208_n1462, DP_mult_208_n1461, DP_mult_208_n1460,
         DP_mult_208_n1459, DP_mult_208_n1458, DP_mult_208_n1457,
         DP_mult_208_n1456, DP_mult_208_n1455, DP_mult_208_n1454,
         DP_mult_208_n1453, DP_mult_208_n1452, DP_mult_208_n1451,
         DP_mult_208_n1450, DP_mult_208_n1449, DP_mult_208_n1448,
         DP_mult_208_n1447, DP_mult_208_n1446, DP_mult_208_n1445,
         DP_mult_208_n1444, DP_mult_208_n1443, DP_mult_208_n1442,
         DP_mult_208_n1441, DP_mult_208_n1440, DP_mult_208_n1439,
         DP_mult_208_n1438, DP_mult_208_n1437, DP_mult_208_n1436,
         DP_mult_208_n1435, DP_mult_208_n1434, DP_mult_208_n1433,
         DP_mult_208_n1432, DP_mult_208_n1431, DP_mult_208_n1430,
         DP_mult_208_n1429, DP_mult_208_n1428, DP_mult_208_n1427,
         DP_mult_208_n1426, DP_mult_208_n1425, DP_mult_208_n1424,
         DP_mult_208_n1423, DP_mult_208_n1422, DP_mult_208_n1421,
         DP_mult_208_n1420, DP_mult_208_n1419, DP_mult_208_n1418,
         DP_mult_208_n1417, DP_mult_208_n1416, DP_mult_208_n1415,
         DP_mult_208_n1414, DP_mult_208_n1413, DP_mult_208_n1412,
         DP_mult_208_n1411, DP_mult_208_n1410, DP_mult_208_n1409,
         DP_mult_208_n1408, DP_mult_208_n1407, DP_mult_208_n1406,
         DP_mult_208_n1405, DP_mult_208_n1404, DP_mult_208_n1403,
         DP_mult_208_n1402, DP_mult_208_n1401, DP_mult_208_n1400,
         DP_mult_208_n1399, DP_mult_208_n1398, DP_mult_208_n1397,
         DP_mult_208_n1396, DP_mult_208_n1395, DP_mult_208_n1394,
         DP_mult_208_n1393, DP_mult_208_n1392, DP_mult_208_n1391,
         DP_mult_208_n1390, DP_mult_208_n1389, DP_mult_208_n1388,
         DP_mult_208_n1387, DP_mult_208_n1386, DP_mult_208_n1385,
         DP_mult_208_n1384, DP_mult_208_n1383, DP_mult_208_n1382,
         DP_mult_208_n1381, DP_mult_208_n1380, DP_mult_208_n1379,
         DP_mult_208_n1378, DP_mult_208_n1377, DP_mult_208_n1376,
         DP_mult_208_n1375, DP_mult_208_n1374, DP_mult_208_n1373,
         DP_mult_208_n1372, DP_mult_208_n1371, DP_mult_208_n1370,
         DP_mult_208_n1369, DP_mult_208_n1368, DP_mult_208_n1367,
         DP_mult_208_n1366, DP_mult_208_n1365, DP_mult_208_n1364,
         DP_mult_208_n1363, DP_mult_208_n1362, DP_mult_208_n1361,
         DP_mult_208_n1360, DP_mult_208_n1359, DP_mult_208_n1358,
         DP_mult_208_n1357, DP_mult_208_n1356, DP_mult_208_n1355,
         DP_mult_208_n1354, DP_mult_208_n1353, DP_mult_208_n1352,
         DP_mult_208_n1351, DP_mult_208_n1350, DP_mult_208_n1349,
         DP_mult_208_n1348, DP_mult_208_n1347, DP_mult_208_n1346,
         DP_mult_208_n1345, DP_mult_208_n1344, DP_mult_208_n1343,
         DP_mult_208_n1342, DP_mult_208_n1341, DP_mult_208_n1340,
         DP_mult_208_n1339, DP_mult_208_n1338, DP_mult_208_n1337,
         DP_mult_208_n1336, DP_mult_208_n1335, DP_mult_208_n1334,
         DP_mult_208_n1333, DP_mult_208_n1332, DP_mult_208_n1331,
         DP_mult_208_n1330, DP_mult_208_n1329, DP_mult_208_n1328,
         DP_mult_208_n1327, DP_mult_208_n1326, DP_mult_208_n1325,
         DP_mult_208_n1324, DP_mult_208_n1323, DP_mult_208_n1322,
         DP_mult_208_n1321, DP_mult_208_n1320, DP_mult_208_n1319,
         DP_mult_208_n1318, DP_mult_208_n1317, DP_mult_208_n1316,
         DP_mult_208_n1315, DP_mult_208_n1314, DP_mult_208_n1313,
         DP_mult_208_n1312, DP_mult_208_n1311, DP_mult_208_n1310,
         DP_mult_208_n1309, DP_mult_208_n1308, DP_mult_208_n1307,
         DP_mult_208_n1306, DP_mult_208_n1305, DP_mult_208_n1304,
         DP_mult_208_n1303, DP_mult_208_n1302, DP_mult_208_n1301,
         DP_mult_208_n1300, DP_mult_208_n1299, DP_mult_208_n1298,
         DP_mult_208_n1297, DP_mult_208_n1296, DP_mult_208_n1295,
         DP_mult_208_n1294, DP_mult_208_n1293, DP_mult_208_n1292,
         DP_mult_208_n1291, DP_mult_208_n1290, DP_mult_208_n1289,
         DP_mult_208_n1288, DP_mult_208_n1287, DP_mult_208_n1286,
         DP_mult_208_n1285, DP_mult_208_n1284, DP_mult_208_n1283,
         DP_mult_208_n1282, DP_mult_208_n1281, DP_mult_208_n1280,
         DP_mult_208_n1279, DP_mult_208_n1278, DP_mult_208_n1277,
         DP_mult_208_n1276, DP_mult_208_n1275, DP_mult_208_n1274,
         DP_mult_208_n1273, DP_mult_208_n1272, DP_mult_208_n1271,
         DP_mult_208_n1270, DP_mult_208_n1269, DP_mult_208_n1268,
         DP_mult_208_n1267, DP_mult_208_n1266, DP_mult_208_n1265,
         DP_mult_208_n1264, DP_mult_208_n1263, DP_mult_208_n1262,
         DP_mult_208_n1261, DP_mult_208_n1260, DP_mult_208_n1259,
         DP_mult_208_n1258, DP_mult_208_n1257, DP_mult_208_n1256,
         DP_mult_208_n1255, DP_mult_208_n1254, DP_mult_208_n1253,
         DP_mult_208_n1252, DP_mult_208_n1251, DP_mult_208_n1250,
         DP_mult_208_n1249, DP_mult_208_n1248, DP_mult_208_n1247,
         DP_mult_208_n1246, DP_mult_208_n1245, DP_mult_208_n1244,
         DP_mult_208_n1243, DP_mult_208_n1242, DP_mult_208_n1241,
         DP_mult_208_n1240, DP_mult_208_n1239, DP_mult_208_n1238,
         DP_mult_208_n1237, DP_mult_208_n1236, DP_mult_208_n1235,
         DP_mult_208_n1234, DP_mult_208_n1233, DP_mult_208_n1232,
         DP_mult_208_n1231, DP_mult_208_n1230, DP_mult_208_n1229,
         DP_mult_208_n1228, DP_mult_208_n1227, DP_mult_208_n1226,
         DP_mult_208_n1225, DP_mult_208_n1224, DP_mult_208_n1223,
         DP_mult_208_n1222, DP_mult_208_n1221, DP_mult_208_n1220,
         DP_mult_208_n1219, DP_mult_208_n1218, DP_mult_208_n1217,
         DP_mult_208_n1216, DP_mult_208_n1215, DP_mult_208_n1214,
         DP_mult_208_n1213, DP_mult_208_n1212, DP_mult_208_n1211,
         DP_mult_208_n1210, DP_mult_208_n1209, DP_mult_208_n1208,
         DP_mult_208_n1207, DP_mult_208_n1206, DP_mult_208_n1205,
         DP_mult_208_n1204, DP_mult_208_n1203, DP_mult_208_n1202,
         DP_mult_208_n1201, DP_mult_208_n1200, DP_mult_208_n1199,
         DP_mult_208_n1198, DP_mult_208_n1197, DP_mult_208_n1196,
         DP_mult_208_n1195, DP_mult_208_n1194, DP_mult_208_n1193,
         DP_mult_208_n1192, DP_mult_208_n1191, DP_mult_208_n1190,
         DP_mult_208_n1189, DP_mult_208_n1188, DP_mult_208_n1187,
         DP_mult_208_n1186, DP_mult_208_n1185, DP_mult_208_n1184,
         DP_mult_208_n1183, DP_mult_208_n1182, DP_mult_208_n1181,
         DP_mult_208_n1180, DP_mult_208_n1179, DP_mult_208_n1178,
         DP_mult_208_n1177, DP_mult_208_n1176, DP_mult_208_n1175,
         DP_mult_208_n1174, DP_mult_208_n1173, DP_mult_208_n1172,
         DP_mult_208_n1171, DP_mult_208_n1170, DP_mult_208_n1169,
         DP_mult_208_n1168, DP_mult_208_n1167, DP_mult_208_n1166,
         DP_mult_208_n1165, DP_mult_208_n1164, DP_mult_208_n1163,
         DP_mult_208_n1162, DP_mult_208_n1161, DP_mult_208_n1160,
         DP_mult_208_n1159, DP_mult_208_n1158, DP_mult_208_n1157,
         DP_mult_208_n1156, DP_mult_208_n1155, DP_mult_208_n1154,
         DP_mult_208_n1153, DP_mult_208_n1152, DP_mult_208_n1151,
         DP_mult_208_n1150, DP_mult_208_n1149, DP_mult_208_n1148,
         DP_mult_208_n1147, DP_mult_208_n1146, DP_mult_208_n1145,
         DP_mult_208_n1144, DP_mult_208_n1143, DP_mult_208_n1142,
         DP_mult_208_n1141, DP_mult_208_n1140, DP_mult_208_n1139,
         DP_mult_208_n1138, DP_mult_208_n1137, DP_mult_208_n1136,
         DP_mult_208_n1135, DP_mult_208_n1134, DP_mult_208_n1133,
         DP_mult_208_n1132, DP_mult_208_n1131, DP_mult_208_n1130,
         DP_mult_208_n1129, DP_mult_208_n1128, DP_mult_208_n1127,
         DP_mult_208_n1126, DP_mult_208_n1125, DP_mult_208_n1124,
         DP_mult_208_n1123, DP_mult_208_n1122, DP_mult_208_n1121,
         DP_mult_208_n1120, DP_mult_208_n1119, DP_mult_208_n1118,
         DP_mult_208_n1117, DP_mult_208_n1116, DP_mult_208_n1115,
         DP_mult_208_n1114, DP_mult_208_n1113, DP_mult_208_n1112,
         DP_mult_208_n1111, DP_mult_208_n1110, DP_mult_208_n1109,
         DP_mult_208_n1108, DP_mult_208_n1107, DP_mult_208_n1106,
         DP_mult_208_n1105, DP_mult_208_n1104, DP_mult_208_n1103,
         DP_mult_208_n1102, DP_mult_208_n1101, DP_mult_208_n1100,
         DP_mult_208_n1099, DP_mult_208_n1098, DP_mult_208_n1097,
         DP_mult_208_n1096, DP_mult_208_n1095, DP_mult_208_n1094,
         DP_mult_208_n1093, DP_mult_208_n1092, DP_mult_208_n1091,
         DP_mult_208_n1090, DP_mult_208_n1089, DP_mult_208_n1088,
         DP_mult_208_n1087, DP_mult_208_n1086, DP_mult_208_n1085,
         DP_mult_208_n1084, DP_mult_208_n1083, DP_mult_208_n1082,
         DP_mult_208_n1081, DP_mult_208_n1080, DP_mult_208_n1079,
         DP_mult_208_n1078, DP_mult_208_n1077, DP_mult_208_n1076,
         DP_mult_208_n1075, DP_mult_208_n1074, DP_mult_208_n1073,
         DP_mult_208_n1072, DP_mult_208_n1071, DP_mult_208_n1070,
         DP_mult_208_n1069, DP_mult_208_n1068, DP_mult_208_n1067,
         DP_mult_208_n1066, DP_mult_208_n1065, DP_mult_208_n1064,
         DP_mult_208_n1063, DP_mult_208_n1062, DP_mult_208_n1061,
         DP_mult_208_n1060, DP_mult_208_n1059, DP_mult_208_n1058,
         DP_mult_208_n1057, DP_mult_208_n1056, DP_mult_208_n1055,
         DP_mult_208_n1054, DP_mult_208_n1053, DP_mult_208_n1052,
         DP_mult_208_n1051, DP_mult_208_n1050, DP_mult_208_n1049,
         DP_mult_208_n1048, DP_mult_208_n1047, DP_mult_208_n1046,
         DP_mult_208_n1045, DP_mult_208_n1044, DP_mult_208_n1043,
         DP_mult_208_n1042, DP_mult_208_n1041, DP_mult_208_n1040,
         DP_mult_208_n1039, DP_mult_208_n1038, DP_mult_208_n1037,
         DP_mult_208_n1036, DP_mult_208_n1035, DP_mult_208_n1034,
         DP_mult_208_n1033, DP_mult_208_n1032, DP_mult_208_n1031,
         DP_mult_208_n1030, DP_mult_208_n1029, DP_mult_208_n1028,
         DP_mult_208_n1027, DP_mult_208_n1026, DP_mult_208_n1025,
         DP_mult_208_n1024, DP_mult_208_n1023, DP_mult_208_n1022,
         DP_mult_208_n1021, DP_mult_208_n1020, DP_mult_208_n1019,
         DP_mult_208_n1018, DP_mult_208_n1017, DP_mult_208_n1016,
         DP_mult_208_n1015, DP_mult_208_n1014, DP_mult_208_n1013,
         DP_mult_208_n1012, DP_mult_208_n1011, DP_mult_208_n1010,
         DP_mult_208_n1009, DP_mult_208_n1008, DP_mult_208_n1007,
         DP_mult_208_n1006, DP_mult_208_n1005, DP_mult_208_n1004,
         DP_mult_208_n1003, DP_mult_208_n1002, DP_mult_208_n1001,
         DP_mult_208_n999, DP_mult_208_n998, DP_mult_208_n997,
         DP_mult_208_n996, DP_mult_208_n995, DP_mult_208_n994,
         DP_mult_208_n993, DP_mult_208_n992, DP_mult_208_n991,
         DP_mult_208_n990, DP_mult_208_n989, DP_mult_208_n988,
         DP_mult_208_n987, DP_mult_208_n986, DP_mult_208_n985,
         DP_mult_208_n984, DP_mult_208_n983, DP_mult_208_n982,
         DP_mult_208_n981, DP_mult_208_n980, DP_mult_208_n979,
         DP_mult_208_n978, DP_mult_208_n977, DP_mult_208_n976,
         DP_mult_208_n975, DP_mult_208_n974, DP_mult_208_n973,
         DP_mult_208_n972, DP_mult_208_n971, DP_mult_208_n970,
         DP_mult_208_n969, DP_mult_208_n968, DP_mult_208_n967,
         DP_mult_208_n966, DP_mult_208_n965, DP_mult_208_n964,
         DP_mult_208_n963, DP_mult_208_n962, DP_mult_208_n961,
         DP_mult_208_n959, DP_mult_208_n958, DP_mult_208_n957,
         DP_mult_208_n956, DP_mult_208_n955, DP_mult_208_n954,
         DP_mult_208_n953, DP_mult_208_n952, DP_mult_208_n951,
         DP_mult_208_n950, DP_mult_208_n949, DP_mult_208_n948,
         DP_mult_208_n947, DP_mult_208_n946, DP_mult_208_n945,
         DP_mult_208_n944, DP_mult_208_n943, DP_mult_208_n942,
         DP_mult_208_n941, DP_mult_208_n940, DP_mult_208_n939,
         DP_mult_208_n938, DP_mult_208_n937, DP_mult_208_n936,
         DP_mult_208_n935, DP_mult_208_n934, DP_mult_208_n933,
         DP_mult_208_n932, DP_mult_208_n931, DP_mult_208_n930,
         DP_mult_208_n929, DP_mult_208_n928, DP_mult_208_n927,
         DP_mult_208_n926, DP_mult_208_n925, DP_mult_208_n924,
         DP_mult_208_n923, DP_mult_208_n922, DP_mult_208_n921,
         DP_mult_208_n920, DP_mult_208_n919, DP_mult_208_n918,
         DP_mult_208_n917, DP_mult_208_n916, DP_mult_208_n915,
         DP_mult_208_n914, DP_mult_208_n913, DP_mult_208_n912,
         DP_mult_208_n911, DP_mult_208_n910, DP_mult_208_n909,
         DP_mult_208_n908, DP_mult_208_n907, DP_mult_208_n906,
         DP_mult_208_n905, DP_mult_208_n904, DP_mult_208_n903,
         DP_mult_208_n902, DP_mult_208_n901, DP_mult_208_n900,
         DP_mult_208_n899, DP_mult_208_n898, DP_mult_208_n897,
         DP_mult_208_n896, DP_mult_208_n895, DP_mult_208_n894,
         DP_mult_208_n893, DP_mult_208_n892, DP_mult_208_n891,
         DP_mult_208_n890, DP_mult_208_n889, DP_mult_208_n888,
         DP_mult_208_n887, DP_mult_208_n886, DP_mult_208_n885,
         DP_mult_208_n884, DP_mult_208_n883, DP_mult_208_n882,
         DP_mult_208_n881, DP_mult_208_n880, DP_mult_208_n879,
         DP_mult_208_n878, DP_mult_208_n877, DP_mult_208_n876,
         DP_mult_208_n875, DP_mult_208_n874, DP_mult_208_n873,
         DP_mult_208_n872, DP_mult_208_n871, DP_mult_208_n870,
         DP_mult_208_n869, DP_mult_208_n868, DP_mult_208_n867,
         DP_mult_208_n866, DP_mult_208_n865, DP_mult_208_n864,
         DP_mult_208_n863, DP_mult_208_n862, DP_mult_208_n861,
         DP_mult_208_n860, DP_mult_208_n859, DP_mult_208_n858,
         DP_mult_208_n857, DP_mult_208_n856, DP_mult_208_n855,
         DP_mult_208_n854, DP_mult_208_n853, DP_mult_208_n852,
         DP_mult_208_n851, DP_mult_208_n850, DP_mult_208_n849,
         DP_mult_208_n848, DP_mult_208_n847, DP_mult_208_n846,
         DP_mult_208_n845, DP_mult_208_n844, DP_mult_208_n843,
         DP_mult_208_n842, DP_mult_208_n841, DP_mult_208_n840,
         DP_mult_208_n839, DP_mult_208_n838, DP_mult_208_n837,
         DP_mult_208_n836, DP_mult_208_n835, DP_mult_208_n834,
         DP_mult_208_n833, DP_mult_208_n832, DP_mult_208_n831,
         DP_mult_208_n830, DP_mult_208_n829, DP_mult_208_n828,
         DP_mult_208_n827, DP_mult_208_n826, DP_mult_208_n825,
         DP_mult_208_n824, DP_mult_208_n823, DP_mult_208_n822,
         DP_mult_208_n821, DP_mult_208_n820, DP_mult_208_n819,
         DP_mult_208_n818, DP_mult_208_n817, DP_mult_208_n816,
         DP_mult_208_n815, DP_mult_208_n814, DP_mult_208_n813,
         DP_mult_208_n812, DP_mult_208_n811, DP_mult_208_n810,
         DP_mult_208_n809, DP_mult_208_n808, DP_mult_208_n807,
         DP_mult_208_n806, DP_mult_208_n805, DP_mult_208_n804,
         DP_mult_208_n803, DP_mult_208_n802, DP_mult_208_n801,
         DP_mult_208_n800, DP_mult_208_n799, DP_mult_208_n798,
         DP_mult_208_n797, DP_mult_208_n796, DP_mult_208_n795,
         DP_mult_208_n794, DP_mult_208_n793, DP_mult_208_n792,
         DP_mult_208_n791, DP_mult_208_n790, DP_mult_208_n789,
         DP_mult_208_n788, DP_mult_208_n787, DP_mult_208_n786,
         DP_mult_208_n785, DP_mult_208_n784, DP_mult_208_n783,
         DP_mult_208_n782, DP_mult_208_n781, DP_mult_208_n780,
         DP_mult_208_n779, DP_mult_208_n778, DP_mult_208_n777,
         DP_mult_208_n776, DP_mult_208_n775, DP_mult_208_n774,
         DP_mult_208_n773, DP_mult_208_n772, DP_mult_208_n771,
         DP_mult_208_n770, DP_mult_208_n769, DP_mult_208_n768,
         DP_mult_208_n767, DP_mult_208_n766, DP_mult_208_n765,
         DP_mult_208_n764, DP_mult_208_n763, DP_mult_208_n762,
         DP_mult_208_n761, DP_mult_208_n760, DP_mult_208_n759,
         DP_mult_208_n758, DP_mult_208_n757, DP_mult_208_n756,
         DP_mult_208_n755, DP_mult_208_n754, DP_mult_208_n753,
         DP_mult_208_n752, DP_mult_208_n751, DP_mult_208_n750,
         DP_mult_208_n749, DP_mult_208_n748, DP_mult_208_n747,
         DP_mult_208_n746, DP_mult_208_n745, DP_mult_208_n744,
         DP_mult_208_n743, DP_mult_208_n742, DP_mult_208_n741,
         DP_mult_208_n740, DP_mult_208_n739, DP_mult_208_n738,
         DP_mult_208_n737, DP_mult_208_n736, DP_mult_208_n735,
         DP_mult_208_n734, DP_mult_208_n733, DP_mult_208_n732,
         DP_mult_208_n731, DP_mult_208_n730, DP_mult_208_n729,
         DP_mult_208_n728, DP_mult_208_n727, DP_mult_208_n726,
         DP_mult_208_n725, DP_mult_208_n724, DP_mult_208_n723,
         DP_mult_208_n722, DP_mult_208_n721, DP_mult_208_n720,
         DP_mult_208_n719, DP_mult_208_n718, DP_mult_208_n717,
         DP_mult_208_n716, DP_mult_208_n715, DP_mult_208_n714,
         DP_mult_208_n713, DP_mult_208_n712, DP_mult_208_n711,
         DP_mult_208_n710, DP_mult_208_n709, DP_mult_208_n708,
         DP_mult_208_n707, DP_mult_208_n706, DP_mult_208_n705,
         DP_mult_208_n704, DP_mult_208_n703, DP_mult_208_n702,
         DP_mult_208_n701, DP_mult_208_n700, DP_mult_208_n699,
         DP_mult_208_n698, DP_mult_208_n697, DP_mult_208_n696,
         DP_mult_208_n695, DP_mult_208_n694, DP_mult_208_n693,
         DP_mult_208_n692, DP_mult_208_n691, DP_mult_208_n690,
         DP_mult_208_n689, DP_mult_208_n688, DP_mult_208_n687,
         DP_mult_208_n686, DP_mult_208_n685, DP_mult_208_n684,
         DP_mult_208_n683, DP_mult_208_n682, DP_mult_208_n681,
         DP_mult_208_n680, DP_mult_208_n679, DP_mult_208_n678,
         DP_mult_208_n677, DP_mult_208_n676, DP_mult_208_n675,
         DP_mult_208_n674, DP_mult_208_n672, DP_mult_208_n671,
         DP_mult_208_n670, DP_mult_208_n668, DP_mult_208_n667,
         DP_mult_208_n666, DP_mult_208_n663, DP_mult_208_n662,
         DP_mult_208_n661, DP_mult_208_n657, DP_mult_208_n646,
         DP_mult_208_n645, DP_mult_208_n644, DP_mult_208_n643,
         DP_mult_208_n638, DP_mult_208_n637, DP_mult_208_n636,
         DP_mult_208_n635, DP_mult_208_n634, DP_mult_208_n633,
         DP_mult_208_n632, DP_mult_208_n631, DP_mult_208_n630,
         DP_mult_208_n629, DP_mult_208_n628, DP_mult_208_n627,
         DP_mult_208_n626, DP_mult_208_n625, DP_mult_208_n620,
         DP_mult_208_n611, DP_mult_208_n610, DP_mult_208_n609,
         DP_mult_208_n600, DP_mult_208_n599, DP_mult_208_n598,
         DP_mult_208_n597, DP_mult_208_n596, DP_mult_208_n595,
         DP_mult_208_n594, DP_mult_208_n593, DP_mult_208_n592,
         DP_mult_208_n591, DP_mult_208_n590, DP_mult_208_n589,
         DP_mult_208_n588, DP_mult_208_n583, DP_mult_208_n582,
         DP_mult_208_n581, DP_mult_208_n572, DP_mult_208_n571,
         DP_mult_208_n570, DP_mult_208_n569, DP_mult_208_n568,
         DP_mult_208_n567, DP_mult_208_n566, DP_mult_208_n565,
         DP_mult_208_n564, DP_mult_208_n563, DP_mult_208_n562,
         DP_mult_208_n561, DP_mult_208_n560, DP_mult_208_n559,
         DP_mult_208_n558, DP_mult_208_n555, DP_mult_208_n554,
         DP_mult_208_n553, DP_mult_208_n552, DP_mult_208_n551,
         DP_mult_208_n550, DP_mult_208_n547, DP_mult_208_n546,
         DP_mult_208_n545, DP_mult_208_n544, DP_mult_208_n543,
         DP_mult_208_n542, DP_mult_208_n541, DP_mult_208_n540,
         DP_mult_208_n539, DP_mult_208_n538, DP_mult_208_n537,
         DP_mult_208_n536, DP_mult_208_n535, DP_mult_208_n534,
         DP_mult_208_n533, DP_mult_208_n532, DP_mult_208_n531,
         DP_mult_208_n526, DP_mult_208_n525, DP_mult_208_n524,
         DP_mult_208_n523, DP_mult_208_n522, DP_mult_208_n521,
         DP_mult_208_n520, DP_mult_208_n519, DP_mult_208_n517,
         DP_mult_208_n516, DP_mult_208_n515, DP_mult_208_n514,
         DP_mult_208_n513, DP_mult_208_n511, DP_mult_208_n508,
         DP_mult_208_n507, DP_mult_208_n506, DP_mult_208_n505,
         DP_mult_208_n504, DP_mult_208_n503, DP_mult_208_n502,
         DP_mult_208_n501, DP_mult_208_n499, DP_mult_208_n498,
         DP_mult_208_n497, DP_mult_208_n496, DP_mult_208_n495,
         DP_mult_208_n492, DP_mult_208_n491, DP_mult_208_n490,
         DP_mult_208_n489, DP_mult_208_n488, DP_mult_208_n487,
         DP_mult_208_n486, DP_mult_208_n483, DP_mult_208_n481,
         DP_mult_208_n480, DP_mult_208_n479, DP_mult_208_n478,
         DP_mult_208_n477, DP_mult_208_n476, DP_mult_208_n475,
         DP_mult_208_n474, DP_mult_208_n468, DP_mult_208_n467,
         DP_mult_208_n466, DP_mult_208_n465, DP_mult_208_n464,
         DP_mult_208_n463, DP_mult_208_n462, DP_mult_208_n461,
         DP_mult_208_n459, DP_mult_208_n457, DP_mult_208_n456,
         DP_mult_208_n455, DP_mult_208_n454, DP_mult_208_n453,
         DP_mult_208_n452, DP_mult_208_n451, DP_mult_208_n450,
         DP_mult_208_n448, DP_mult_208_n445, DP_mult_208_n439,
         DP_mult_208_n438, DP_mult_208_n437, DP_mult_208_n436,
         DP_mult_208_n435, DP_mult_208_n434, DP_mult_208_n432,
         DP_mult_208_n431, DP_mult_208_n430, DP_mult_208_n429,
         DP_mult_208_n428, DP_mult_208_n427, DP_mult_208_n426,
         DP_mult_208_n423, DP_mult_208_n422, DP_mult_208_n421,
         DP_mult_208_n420, DP_mult_208_n419, DP_mult_208_n418,
         DP_mult_208_n416, DP_mult_208_n412, DP_mult_208_n411,
         DP_mult_208_n410, DP_mult_208_n409, DP_mult_208_n407,
         DP_mult_208_n405, DP_mult_208_n402, DP_mult_208_n401,
         DP_mult_208_n400, DP_mult_208_n399, DP_mult_208_n398,
         DP_mult_208_n397, DP_mult_208_n396, DP_mult_208_n394,
         DP_mult_208_n390, DP_mult_208_n389, DP_mult_208_n388,
         DP_mult_208_n387, DP_mult_208_n384, DP_mult_208_n383,
         DP_mult_208_n382, DP_mult_208_n381, DP_mult_208_n380,
         DP_mult_208_n379, DP_mult_208_n378, DP_mult_208_n376,
         DP_mult_208_n372, DP_mult_208_n371, DP_mult_208_n370,
         DP_mult_208_n369, DP_mult_208_n367, DP_mult_208_n365,
         DP_mult_208_n364, DP_mult_208_n363, DP_mult_208_n362,
         DP_mult_208_n361, DP_mult_208_n360, DP_mult_208_n359,
         DP_mult_208_n356, DP_mult_208_n355, DP_mult_208_n354,
         DP_mult_208_n353, DP_mult_208_n352, DP_mult_208_n350,
         DP_mult_208_n348, DP_mult_208_n347, DP_mult_208_n346,
         DP_mult_208_n345, DP_mult_208_n344, DP_mult_208_n343,
         DP_mult_208_n342, DP_mult_208_n341, DP_mult_208_n339,
         DP_mult_208_n337, DP_mult_208_n336, DP_mult_208_n335,
         DP_mult_208_n334, DP_mult_208_n333, DP_mult_208_n332,
         DP_mult_208_n327, DP_mult_208_n326, DP_mult_208_n325,
         DP_mult_208_n320, DP_mult_208_n319, DP_mult_208_n318,
         DP_mult_208_n317, DP_mult_208_n316, DP_mult_208_n315,
         DP_mult_208_n314, DP_mult_208_n313, DP_mult_208_n312,
         DP_mult_208_n311, DP_mult_208_n310, DP_mult_208_n309,
         DP_mult_208_n308, DP_mult_208_n307, DP_mult_208_n306,
         DP_mult_208_n305, DP_mult_208_n304, DP_mult_208_n303,
         DP_mult_208_n302, DP_mult_208_n301, DP_mult_208_n277,
         DP_mult_208_n265, DP_mult_208_n251, DP_mult_209_n2317,
         DP_mult_209_n2316, DP_mult_209_n2315, DP_mult_209_n2314,
         DP_mult_209_n2313, DP_mult_209_n2312, DP_mult_209_n2311,
         DP_mult_209_n2310, DP_mult_209_n2309, DP_mult_209_n2308,
         DP_mult_209_n2307, DP_mult_209_n2306, DP_mult_209_n2305,
         DP_mult_209_n2304, DP_mult_209_n2303, DP_mult_209_n2302,
         DP_mult_209_n2301, DP_mult_209_n2300, DP_mult_209_n2299,
         DP_mult_209_n2298, DP_mult_209_n2297, DP_mult_209_n2296,
         DP_mult_209_n2295, DP_mult_209_n2294, DP_mult_209_n2293,
         DP_mult_209_n2292, DP_mult_209_n2291, DP_mult_209_n2290,
         DP_mult_209_n2289, DP_mult_209_n2288, DP_mult_209_n2287,
         DP_mult_209_n2286, DP_mult_209_n2285, DP_mult_209_n2284,
         DP_mult_209_n2283, DP_mult_209_n2282, DP_mult_209_n2281,
         DP_mult_209_n2280, DP_mult_209_n2279, DP_mult_209_n2278,
         DP_mult_209_n2277, DP_mult_209_n2276, DP_mult_209_n2275,
         DP_mult_209_n2274, DP_mult_209_n2273, DP_mult_209_n2272,
         DP_mult_209_n2271, DP_mult_209_n2270, DP_mult_209_n2269,
         DP_mult_209_n2268, DP_mult_209_n2267, DP_mult_209_n2266,
         DP_mult_209_n2265, DP_mult_209_n2264, DP_mult_209_n2263,
         DP_mult_209_n2262, DP_mult_209_n2261, DP_mult_209_n2260,
         DP_mult_209_n2259, DP_mult_209_n2258, DP_mult_209_n2257,
         DP_mult_209_n2256, DP_mult_209_n2255, DP_mult_209_n2254,
         DP_mult_209_n2253, DP_mult_209_n2252, DP_mult_209_n2251,
         DP_mult_209_n2250, DP_mult_209_n2249, DP_mult_209_n2248,
         DP_mult_209_n2247, DP_mult_209_n2246, DP_mult_209_n2245,
         DP_mult_209_n2244, DP_mult_209_n2243, DP_mult_209_n2242,
         DP_mult_209_n2241, DP_mult_209_n2240, DP_mult_209_n2239,
         DP_mult_209_n2238, DP_mult_209_n2237, DP_mult_209_n2236,
         DP_mult_209_n2235, DP_mult_209_n2234, DP_mult_209_n2233,
         DP_mult_209_n2232, DP_mult_209_n2231, DP_mult_209_n2230,
         DP_mult_209_n2229, DP_mult_209_n2228, DP_mult_209_n2227,
         DP_mult_209_n2226, DP_mult_209_n2225, DP_mult_209_n2224,
         DP_mult_209_n2223, DP_mult_209_n2222, DP_mult_209_n2221,
         DP_mult_209_n2220, DP_mult_209_n2219, DP_mult_209_n2218,
         DP_mult_209_n2217, DP_mult_209_n2216, DP_mult_209_n2215,
         DP_mult_209_n2214, DP_mult_209_n2213, DP_mult_209_n2212,
         DP_mult_209_n2211, DP_mult_209_n2210, DP_mult_209_n2209,
         DP_mult_209_n2208, DP_mult_209_n2207, DP_mult_209_n2206,
         DP_mult_209_n2205, DP_mult_209_n2204, DP_mult_209_n2203,
         DP_mult_209_n2202, DP_mult_209_n2201, DP_mult_209_n2200,
         DP_mult_209_n2199, DP_mult_209_n2198, DP_mult_209_n2197,
         DP_mult_209_n2196, DP_mult_209_n2195, DP_mult_209_n2194,
         DP_mult_209_n2193, DP_mult_209_n2192, DP_mult_209_n2191,
         DP_mult_209_n2190, DP_mult_209_n2189, DP_mult_209_n2188,
         DP_mult_209_n2187, DP_mult_209_n2186, DP_mult_209_n2185,
         DP_mult_209_n2184, DP_mult_209_n2183, DP_mult_209_n2182,
         DP_mult_209_n2181, DP_mult_209_n2180, DP_mult_209_n2179,
         DP_mult_209_n2178, DP_mult_209_n2177, DP_mult_209_n2176,
         DP_mult_209_n2175, DP_mult_209_n2174, DP_mult_209_n2173,
         DP_mult_209_n2172, DP_mult_209_n2171, DP_mult_209_n2170,
         DP_mult_209_n2169, DP_mult_209_n2168, DP_mult_209_n2167,
         DP_mult_209_n2166, DP_mult_209_n2165, DP_mult_209_n2164,
         DP_mult_209_n2163, DP_mult_209_n2162, DP_mult_209_n2161,
         DP_mult_209_n2160, DP_mult_209_n2159, DP_mult_209_n2158,
         DP_mult_209_n2157, DP_mult_209_n2156, DP_mult_209_n2155,
         DP_mult_209_n2154, DP_mult_209_n2153, DP_mult_209_n2152,
         DP_mult_209_n2151, DP_mult_209_n2150, DP_mult_209_n2149,
         DP_mult_209_n2148, DP_mult_209_n2147, DP_mult_209_n2146,
         DP_mult_209_n2145, DP_mult_209_n2144, DP_mult_209_n2143,
         DP_mult_209_n2142, DP_mult_209_n2141, DP_mult_209_n2140,
         DP_mult_209_n2139, DP_mult_209_n2138, DP_mult_209_n2137,
         DP_mult_209_n2136, DP_mult_209_n2135, DP_mult_209_n2134,
         DP_mult_209_n2133, DP_mult_209_n2132, DP_mult_209_n2131,
         DP_mult_209_n2130, DP_mult_209_n2129, DP_mult_209_n2128,
         DP_mult_209_n2127, DP_mult_209_n2126, DP_mult_209_n2125,
         DP_mult_209_n2124, DP_mult_209_n2123, DP_mult_209_n2122,
         DP_mult_209_n2121, DP_mult_209_n2120, DP_mult_209_n2119,
         DP_mult_209_n2118, DP_mult_209_n2117, DP_mult_209_n2116,
         DP_mult_209_n2115, DP_mult_209_n2114, DP_mult_209_n2113,
         DP_mult_209_n2112, DP_mult_209_n2111, DP_mult_209_n2110,
         DP_mult_209_n2109, DP_mult_209_n2108, DP_mult_209_n2107,
         DP_mult_209_n2106, DP_mult_209_n2105, DP_mult_209_n2104,
         DP_mult_209_n2103, DP_mult_209_n2102, DP_mult_209_n2101,
         DP_mult_209_n2100, DP_mult_209_n2099, DP_mult_209_n2098,
         DP_mult_209_n2097, DP_mult_209_n2096, DP_mult_209_n2095,
         DP_mult_209_n2094, DP_mult_209_n2093, DP_mult_209_n2092,
         DP_mult_209_n2091, DP_mult_209_n2090, DP_mult_209_n2089,
         DP_mult_209_n2088, DP_mult_209_n2087, DP_mult_209_n2086,
         DP_mult_209_n2085, DP_mult_209_n2084, DP_mult_209_n2083,
         DP_mult_209_n2082, DP_mult_209_n2081, DP_mult_209_n2080,
         DP_mult_209_n2079, DP_mult_209_n2078, DP_mult_209_n2077,
         DP_mult_209_n2076, DP_mult_209_n2075, DP_mult_209_n2074,
         DP_mult_209_n2073, DP_mult_209_n2072, DP_mult_209_n2071,
         DP_mult_209_n2070, DP_mult_209_n2069, DP_mult_209_n2068,
         DP_mult_209_n2067, DP_mult_209_n2066, DP_mult_209_n2065,
         DP_mult_209_n2064, DP_mult_209_n2063, DP_mult_209_n2062,
         DP_mult_209_n2061, DP_mult_209_n2060, DP_mult_209_n2059,
         DP_mult_209_n2058, DP_mult_209_n2057, DP_mult_209_n2056,
         DP_mult_209_n2055, DP_mult_209_n2054, DP_mult_209_n2053,
         DP_mult_209_n2052, DP_mult_209_n2051, DP_mult_209_n2050,
         DP_mult_209_n2049, DP_mult_209_n2048, DP_mult_209_n2047,
         DP_mult_209_n2046, DP_mult_209_n2045, DP_mult_209_n2044,
         DP_mult_209_n2043, DP_mult_209_n2042, DP_mult_209_n2041,
         DP_mult_209_n2040, DP_mult_209_n2039, DP_mult_209_n2038,
         DP_mult_209_n2037, DP_mult_209_n2036, DP_mult_209_n2035,
         DP_mult_209_n2034, DP_mult_209_n2033, DP_mult_209_n2032,
         DP_mult_209_n2031, DP_mult_209_n2030, DP_mult_209_n2029,
         DP_mult_209_n2028, DP_mult_209_n2027, DP_mult_209_n2026,
         DP_mult_209_n2025, DP_mult_209_n2024, DP_mult_209_n2023,
         DP_mult_209_n2022, DP_mult_209_n2021, DP_mult_209_n2020,
         DP_mult_209_n2019, DP_mult_209_n2018, DP_mult_209_n2017,
         DP_mult_209_n2016, DP_mult_209_n2015, DP_mult_209_n2014,
         DP_mult_209_n2013, DP_mult_209_n2012, DP_mult_209_n2011,
         DP_mult_209_n2010, DP_mult_209_n2009, DP_mult_209_n2008,
         DP_mult_209_n2007, DP_mult_209_n2006, DP_mult_209_n2005,
         DP_mult_209_n2004, DP_mult_209_n2003, DP_mult_209_n2002,
         DP_mult_209_n2001, DP_mult_209_n2000, DP_mult_209_n1999,
         DP_mult_209_n1998, DP_mult_209_n1997, DP_mult_209_n1996,
         DP_mult_209_n1995, DP_mult_209_n1994, DP_mult_209_n1993,
         DP_mult_209_n1992, DP_mult_209_n1991, DP_mult_209_n1990,
         DP_mult_209_n1989, DP_mult_209_n1988, DP_mult_209_n1987,
         DP_mult_209_n1986, DP_mult_209_n1985, DP_mult_209_n1984,
         DP_mult_209_n1983, DP_mult_209_n1982, DP_mult_209_n1981,
         DP_mult_209_n1980, DP_mult_209_n1979, DP_mult_209_n1978,
         DP_mult_209_n1977, DP_mult_209_n1976, DP_mult_209_n1975,
         DP_mult_209_n1974, DP_mult_209_n1973, DP_mult_209_n1972,
         DP_mult_209_n1971, DP_mult_209_n1970, DP_mult_209_n1969,
         DP_mult_209_n1968, DP_mult_209_n1967, DP_mult_209_n1966,
         DP_mult_209_n1965, DP_mult_209_n1964, DP_mult_209_n1963,
         DP_mult_209_n1962, DP_mult_209_n1961, DP_mult_209_n1960,
         DP_mult_209_n1959, DP_mult_209_n1958, DP_mult_209_n1957,
         DP_mult_209_n1956, DP_mult_209_n1955, DP_mult_209_n1954,
         DP_mult_209_n1953, DP_mult_209_n1952, DP_mult_209_n1951,
         DP_mult_209_n1950, DP_mult_209_n1949, DP_mult_209_n1948,
         DP_mult_209_n1947, DP_mult_209_n1946, DP_mult_209_n1945,
         DP_mult_209_n1944, DP_mult_209_n1943, DP_mult_209_n1942,
         DP_mult_209_n1941, DP_mult_209_n1940, DP_mult_209_n1939,
         DP_mult_209_n1938, DP_mult_209_n1937, DP_mult_209_n1936,
         DP_mult_209_n1935, DP_mult_209_n1934, DP_mult_209_n1933,
         DP_mult_209_n1932, DP_mult_209_n1931, DP_mult_209_n1930,
         DP_mult_209_n1929, DP_mult_209_n1817, DP_mult_209_n1816,
         DP_mult_209_n1815, DP_mult_209_n1814, DP_mult_209_n1813,
         DP_mult_209_n1812, DP_mult_209_n1811, DP_mult_209_n1810,
         DP_mult_209_n1809, DP_mult_209_n1808, DP_mult_209_n1807,
         DP_mult_209_n1806, DP_mult_209_n1781, DP_mult_209_n1780,
         DP_mult_209_n1779, DP_mult_209_n1778, DP_mult_209_n1777,
         DP_mult_209_n1776, DP_mult_209_n1775, DP_mult_209_n1774,
         DP_mult_209_n1773, DP_mult_209_n1772, DP_mult_209_n1771,
         DP_mult_209_n1770, DP_mult_209_n1769, DP_mult_209_n1768,
         DP_mult_209_n1767, DP_mult_209_n1766, DP_mult_209_n1765,
         DP_mult_209_n1764, DP_mult_209_n1763, DP_mult_209_n1762,
         DP_mult_209_n1761, DP_mult_209_n1760, DP_mult_209_n1759,
         DP_mult_209_n1758, DP_mult_209_n1757, DP_mult_209_n1756,
         DP_mult_209_n1755, DP_mult_209_n1754, DP_mult_209_n1753,
         DP_mult_209_n1752, DP_mult_209_n1751, DP_mult_209_n1750,
         DP_mult_209_n1749, DP_mult_209_n1748, DP_mult_209_n1747,
         DP_mult_209_n1746, DP_mult_209_n1745, DP_mult_209_n1744,
         DP_mult_209_n1743, DP_mult_209_n1742, DP_mult_209_n1741,
         DP_mult_209_n1740, DP_mult_209_n1739, DP_mult_209_n1738,
         DP_mult_209_n1737, DP_mult_209_n1736, DP_mult_209_n1735,
         DP_mult_209_n1734, DP_mult_209_n1733, DP_mult_209_n1732,
         DP_mult_209_n1731, DP_mult_209_n1730, DP_mult_209_n1729,
         DP_mult_209_n1728, DP_mult_209_n1727, DP_mult_209_n1726,
         DP_mult_209_n1725, DP_mult_209_n1724, DP_mult_209_n1723,
         DP_mult_209_n1722, DP_mult_209_n1721, DP_mult_209_n1720,
         DP_mult_209_n1719, DP_mult_209_n1718, DP_mult_209_n1717,
         DP_mult_209_n1716, DP_mult_209_n1715, DP_mult_209_n1714,
         DP_mult_209_n1713, DP_mult_209_n1712, DP_mult_209_n1711,
         DP_mult_209_n1710, DP_mult_209_n1709, DP_mult_209_n1708,
         DP_mult_209_n1707, DP_mult_209_n1706, DP_mult_209_n1705,
         DP_mult_209_n1704, DP_mult_209_n1703, DP_mult_209_n1702,
         DP_mult_209_n1701, DP_mult_209_n1700, DP_mult_209_n1699,
         DP_mult_209_n1698, DP_mult_209_n1697, DP_mult_209_n1696,
         DP_mult_209_n1695, DP_mult_209_n1694, DP_mult_209_n1693,
         DP_mult_209_n1692, DP_mult_209_n1691, DP_mult_209_n1690,
         DP_mult_209_n1689, DP_mult_209_n1688, DP_mult_209_n1687,
         DP_mult_209_n1686, DP_mult_209_n1685, DP_mult_209_n1684,
         DP_mult_209_n1683, DP_mult_209_n1682, DP_mult_209_n1681,
         DP_mult_209_n1680, DP_mult_209_n1679, DP_mult_209_n1678,
         DP_mult_209_n1677, DP_mult_209_n1676, DP_mult_209_n1675,
         DP_mult_209_n1674, DP_mult_209_n1673, DP_mult_209_n1672,
         DP_mult_209_n1671, DP_mult_209_n1670, DP_mult_209_n1669,
         DP_mult_209_n1668, DP_mult_209_n1667, DP_mult_209_n1666,
         DP_mult_209_n1665, DP_mult_209_n1664, DP_mult_209_n1663,
         DP_mult_209_n1662, DP_mult_209_n1661, DP_mult_209_n1660,
         DP_mult_209_n1659, DP_mult_209_n1658, DP_mult_209_n1657,
         DP_mult_209_n1656, DP_mult_209_n1655, DP_mult_209_n1654,
         DP_mult_209_n1653, DP_mult_209_n1652, DP_mult_209_n1651,
         DP_mult_209_n1650, DP_mult_209_n1649, DP_mult_209_n1648,
         DP_mult_209_n1647, DP_mult_209_n1646, DP_mult_209_n1645,
         DP_mult_209_n1644, DP_mult_209_n1643, DP_mult_209_n1642,
         DP_mult_209_n1641, DP_mult_209_n1640, DP_mult_209_n1639,
         DP_mult_209_n1638, DP_mult_209_n1637, DP_mult_209_n1636,
         DP_mult_209_n1635, DP_mult_209_n1634, DP_mult_209_n1633,
         DP_mult_209_n1632, DP_mult_209_n1631, DP_mult_209_n1630,
         DP_mult_209_n1629, DP_mult_209_n1628, DP_mult_209_n1627,
         DP_mult_209_n1626, DP_mult_209_n1625, DP_mult_209_n1624,
         DP_mult_209_n1623, DP_mult_209_n1622, DP_mult_209_n1621,
         DP_mult_209_n1620, DP_mult_209_n1619, DP_mult_209_n1618,
         DP_mult_209_n1617, DP_mult_209_n1616, DP_mult_209_n1615,
         DP_mult_209_n1614, DP_mult_209_n1613, DP_mult_209_n1612,
         DP_mult_209_n1611, DP_mult_209_n1610, DP_mult_209_n1609,
         DP_mult_209_n1608, DP_mult_209_n1607, DP_mult_209_n1606,
         DP_mult_209_n1605, DP_mult_209_n1604, DP_mult_209_n1603,
         DP_mult_209_n1602, DP_mult_209_n1601, DP_mult_209_n1600,
         DP_mult_209_n1599, DP_mult_209_n1598, DP_mult_209_n1597,
         DP_mult_209_n1596, DP_mult_209_n1595, DP_mult_209_n1594,
         DP_mult_209_n1593, DP_mult_209_n1592, DP_mult_209_n1591,
         DP_mult_209_n1590, DP_mult_209_n1589, DP_mult_209_n1588,
         DP_mult_209_n1587, DP_mult_209_n1586, DP_mult_209_n1585,
         DP_mult_209_n1584, DP_mult_209_n1583, DP_mult_209_n1582,
         DP_mult_209_n1581, DP_mult_209_n1580, DP_mult_209_n1579,
         DP_mult_209_n1578, DP_mult_209_n1577, DP_mult_209_n1576,
         DP_mult_209_n1575, DP_mult_209_n1574, DP_mult_209_n1573,
         DP_mult_209_n1572, DP_mult_209_n1571, DP_mult_209_n1570,
         DP_mult_209_n1569, DP_mult_209_n1568, DP_mult_209_n1567,
         DP_mult_209_n1566, DP_mult_209_n1565, DP_mult_209_n1564,
         DP_mult_209_n1563, DP_mult_209_n1562, DP_mult_209_n1561,
         DP_mult_209_n1560, DP_mult_209_n1559, DP_mult_209_n1558,
         DP_mult_209_n1557, DP_mult_209_n1556, DP_mult_209_n1555,
         DP_mult_209_n1554, DP_mult_209_n1553, DP_mult_209_n1552,
         DP_mult_209_n1551, DP_mult_209_n1550, DP_mult_209_n1549,
         DP_mult_209_n1548, DP_mult_209_n1547, DP_mult_209_n1546,
         DP_mult_209_n1545, DP_mult_209_n1544, DP_mult_209_n1543,
         DP_mult_209_n1542, DP_mult_209_n1541, DP_mult_209_n1540,
         DP_mult_209_n1539, DP_mult_209_n1538, DP_mult_209_n1537,
         DP_mult_209_n1536, DP_mult_209_n1535, DP_mult_209_n1534,
         DP_mult_209_n1533, DP_mult_209_n1532, DP_mult_209_n1531,
         DP_mult_209_n1530, DP_mult_209_n1529, DP_mult_209_n1528,
         DP_mult_209_n1527, DP_mult_209_n1526, DP_mult_209_n1525,
         DP_mult_209_n1524, DP_mult_209_n1523, DP_mult_209_n1522,
         DP_mult_209_n1521, DP_mult_209_n1520, DP_mult_209_n1519,
         DP_mult_209_n1518, DP_mult_209_n1517, DP_mult_209_n1516,
         DP_mult_209_n1515, DP_mult_209_n1514, DP_mult_209_n1513,
         DP_mult_209_n1512, DP_mult_209_n1511, DP_mult_209_n1510,
         DP_mult_209_n1509, DP_mult_209_n1508, DP_mult_209_n1507,
         DP_mult_209_n1506, DP_mult_209_n1505, DP_mult_209_n1504,
         DP_mult_209_n1503, DP_mult_209_n1502, DP_mult_209_n1501,
         DP_mult_209_n1500, DP_mult_209_n1499, DP_mult_209_n1498,
         DP_mult_209_n1497, DP_mult_209_n1496, DP_mult_209_n1495,
         DP_mult_209_n1494, DP_mult_209_n1493, DP_mult_209_n1492,
         DP_mult_209_n1491, DP_mult_209_n1490, DP_mult_209_n1489,
         DP_mult_209_n1488, DP_mult_209_n1487, DP_mult_209_n1486,
         DP_mult_209_n1485, DP_mult_209_n1484, DP_mult_209_n1483,
         DP_mult_209_n1482, DP_mult_209_n1481, DP_mult_209_n1480,
         DP_mult_209_n1479, DP_mult_209_n1478, DP_mult_209_n1477,
         DP_mult_209_n1476, DP_mult_209_n1475, DP_mult_209_n1474,
         DP_mult_209_n1473, DP_mult_209_n1472, DP_mult_209_n1471,
         DP_mult_209_n1470, DP_mult_209_n1469, DP_mult_209_n1468,
         DP_mult_209_n1467, DP_mult_209_n1466, DP_mult_209_n1465,
         DP_mult_209_n1464, DP_mult_209_n1463, DP_mult_209_n1462,
         DP_mult_209_n1461, DP_mult_209_n1460, DP_mult_209_n1459,
         DP_mult_209_n1458, DP_mult_209_n1457, DP_mult_209_n1456,
         DP_mult_209_n1455, DP_mult_209_n1454, DP_mult_209_n1453,
         DP_mult_209_n1452, DP_mult_209_n1451, DP_mult_209_n1450,
         DP_mult_209_n1449, DP_mult_209_n1448, DP_mult_209_n1447,
         DP_mult_209_n1446, DP_mult_209_n1445, DP_mult_209_n1444,
         DP_mult_209_n1443, DP_mult_209_n1442, DP_mult_209_n1441,
         DP_mult_209_n1440, DP_mult_209_n1439, DP_mult_209_n1438,
         DP_mult_209_n1437, DP_mult_209_n1436, DP_mult_209_n1435,
         DP_mult_209_n1434, DP_mult_209_n1433, DP_mult_209_n1432,
         DP_mult_209_n1431, DP_mult_209_n1430, DP_mult_209_n1429,
         DP_mult_209_n1428, DP_mult_209_n1427, DP_mult_209_n1426,
         DP_mult_209_n1425, DP_mult_209_n1424, DP_mult_209_n1423,
         DP_mult_209_n1422, DP_mult_209_n1421, DP_mult_209_n1420,
         DP_mult_209_n1419, DP_mult_209_n1418, DP_mult_209_n1417,
         DP_mult_209_n1416, DP_mult_209_n1415, DP_mult_209_n1414,
         DP_mult_209_n1413, DP_mult_209_n1412, DP_mult_209_n1411,
         DP_mult_209_n1410, DP_mult_209_n1409, DP_mult_209_n1408,
         DP_mult_209_n1407, DP_mult_209_n1406, DP_mult_209_n1405,
         DP_mult_209_n1404, DP_mult_209_n1403, DP_mult_209_n1402,
         DP_mult_209_n1401, DP_mult_209_n1400, DP_mult_209_n1399,
         DP_mult_209_n1398, DP_mult_209_n1397, DP_mult_209_n1396,
         DP_mult_209_n1395, DP_mult_209_n1394, DP_mult_209_n1393,
         DP_mult_209_n1392, DP_mult_209_n1391, DP_mult_209_n1390,
         DP_mult_209_n1389, DP_mult_209_n1388, DP_mult_209_n1387,
         DP_mult_209_n1386, DP_mult_209_n1385, DP_mult_209_n1384,
         DP_mult_209_n1383, DP_mult_209_n1382, DP_mult_209_n1381,
         DP_mult_209_n1380, DP_mult_209_n1379, DP_mult_209_n1378,
         DP_mult_209_n1377, DP_mult_209_n1376, DP_mult_209_n1375,
         DP_mult_209_n1374, DP_mult_209_n1373, DP_mult_209_n1372,
         DP_mult_209_n1371, DP_mult_209_n1370, DP_mult_209_n1369,
         DP_mult_209_n1368, DP_mult_209_n1367, DP_mult_209_n1366,
         DP_mult_209_n1365, DP_mult_209_n1364, DP_mult_209_n1363,
         DP_mult_209_n1362, DP_mult_209_n1361, DP_mult_209_n1360,
         DP_mult_209_n1359, DP_mult_209_n1358, DP_mult_209_n1357,
         DP_mult_209_n1356, DP_mult_209_n1355, DP_mult_209_n1354,
         DP_mult_209_n1353, DP_mult_209_n1352, DP_mult_209_n1351,
         DP_mult_209_n1350, DP_mult_209_n1349, DP_mult_209_n1348,
         DP_mult_209_n1347, DP_mult_209_n1346, DP_mult_209_n1345,
         DP_mult_209_n1344, DP_mult_209_n1343, DP_mult_209_n1342,
         DP_mult_209_n1341, DP_mult_209_n1340, DP_mult_209_n1339,
         DP_mult_209_n1338, DP_mult_209_n1337, DP_mult_209_n1336,
         DP_mult_209_n1335, DP_mult_209_n1334, DP_mult_209_n1333,
         DP_mult_209_n1332, DP_mult_209_n1331, DP_mult_209_n1330,
         DP_mult_209_n1329, DP_mult_209_n1328, DP_mult_209_n1327,
         DP_mult_209_n1326, DP_mult_209_n1325, DP_mult_209_n1324,
         DP_mult_209_n1323, DP_mult_209_n1322, DP_mult_209_n1321,
         DP_mult_209_n1320, DP_mult_209_n1319, DP_mult_209_n1318,
         DP_mult_209_n1317, DP_mult_209_n1316, DP_mult_209_n1315,
         DP_mult_209_n1314, DP_mult_209_n1313, DP_mult_209_n1312,
         DP_mult_209_n1311, DP_mult_209_n1310, DP_mult_209_n1309,
         DP_mult_209_n1308, DP_mult_209_n1307, DP_mult_209_n1306,
         DP_mult_209_n1305, DP_mult_209_n1304, DP_mult_209_n1303,
         DP_mult_209_n1302, DP_mult_209_n1301, DP_mult_209_n1300,
         DP_mult_209_n1299, DP_mult_209_n1298, DP_mult_209_n1297,
         DP_mult_209_n1296, DP_mult_209_n1295, DP_mult_209_n1294,
         DP_mult_209_n1293, DP_mult_209_n1292, DP_mult_209_n1291,
         DP_mult_209_n1290, DP_mult_209_n1289, DP_mult_209_n1288,
         DP_mult_209_n1287, DP_mult_209_n1286, DP_mult_209_n1285,
         DP_mult_209_n1284, DP_mult_209_n1283, DP_mult_209_n1282,
         DP_mult_209_n1281, DP_mult_209_n1280, DP_mult_209_n1279,
         DP_mult_209_n1278, DP_mult_209_n1277, DP_mult_209_n1276,
         DP_mult_209_n1275, DP_mult_209_n1274, DP_mult_209_n1273,
         DP_mult_209_n1272, DP_mult_209_n1271, DP_mult_209_n1270,
         DP_mult_209_n1269, DP_mult_209_n1268, DP_mult_209_n1267,
         DP_mult_209_n1266, DP_mult_209_n1265, DP_mult_209_n1264,
         DP_mult_209_n1263, DP_mult_209_n1262, DP_mult_209_n1261,
         DP_mult_209_n1260, DP_mult_209_n1259, DP_mult_209_n1258,
         DP_mult_209_n1257, DP_mult_209_n1256, DP_mult_209_n1255,
         DP_mult_209_n1254, DP_mult_209_n1253, DP_mult_209_n1252,
         DP_mult_209_n1251, DP_mult_209_n1250, DP_mult_209_n1249,
         DP_mult_209_n1248, DP_mult_209_n1247, DP_mult_209_n1246,
         DP_mult_209_n1245, DP_mult_209_n1244, DP_mult_209_n1243,
         DP_mult_209_n1242, DP_mult_209_n1241, DP_mult_209_n1240,
         DP_mult_209_n1239, DP_mult_209_n1238, DP_mult_209_n1237,
         DP_mult_209_n1236, DP_mult_209_n1235, DP_mult_209_n1234,
         DP_mult_209_n1233, DP_mult_209_n1232, DP_mult_209_n1231,
         DP_mult_209_n1230, DP_mult_209_n1229, DP_mult_209_n1228,
         DP_mult_209_n1227, DP_mult_209_n1226, DP_mult_209_n1225,
         DP_mult_209_n1224, DP_mult_209_n1223, DP_mult_209_n1222,
         DP_mult_209_n1221, DP_mult_209_n1220, DP_mult_209_n1219,
         DP_mult_209_n1218, DP_mult_209_n1217, DP_mult_209_n1216,
         DP_mult_209_n1215, DP_mult_209_n1214, DP_mult_209_n1213,
         DP_mult_209_n1212, DP_mult_209_n1211, DP_mult_209_n1210,
         DP_mult_209_n1209, DP_mult_209_n1208, DP_mult_209_n1207,
         DP_mult_209_n1206, DP_mult_209_n1205, DP_mult_209_n1204,
         DP_mult_209_n1203, DP_mult_209_n1202, DP_mult_209_n1201,
         DP_mult_209_n1200, DP_mult_209_n1199, DP_mult_209_n1198,
         DP_mult_209_n1197, DP_mult_209_n1196, DP_mult_209_n1195,
         DP_mult_209_n1194, DP_mult_209_n1193, DP_mult_209_n1192,
         DP_mult_209_n1191, DP_mult_209_n1190, DP_mult_209_n1189,
         DP_mult_209_n1188, DP_mult_209_n1187, DP_mult_209_n1186,
         DP_mult_209_n1185, DP_mult_209_n1184, DP_mult_209_n1183,
         DP_mult_209_n1182, DP_mult_209_n1181, DP_mult_209_n1180,
         DP_mult_209_n1179, DP_mult_209_n1178, DP_mult_209_n1177,
         DP_mult_209_n1176, DP_mult_209_n1175, DP_mult_209_n1174,
         DP_mult_209_n1173, DP_mult_209_n1172, DP_mult_209_n1171,
         DP_mult_209_n1170, DP_mult_209_n1169, DP_mult_209_n1168,
         DP_mult_209_n1167, DP_mult_209_n1166, DP_mult_209_n1165,
         DP_mult_209_n1164, DP_mult_209_n1163, DP_mult_209_n1162,
         DP_mult_209_n1161, DP_mult_209_n1160, DP_mult_209_n1159,
         DP_mult_209_n1158, DP_mult_209_n1157, DP_mult_209_n1156,
         DP_mult_209_n1155, DP_mult_209_n1154, DP_mult_209_n1153,
         DP_mult_209_n1152, DP_mult_209_n1151, DP_mult_209_n1150,
         DP_mult_209_n1149, DP_mult_209_n1148, DP_mult_209_n1147,
         DP_mult_209_n1146, DP_mult_209_n1145, DP_mult_209_n1144,
         DP_mult_209_n1143, DP_mult_209_n1142, DP_mult_209_n1141,
         DP_mult_209_n1140, DP_mult_209_n1139, DP_mult_209_n1138,
         DP_mult_209_n1137, DP_mult_209_n1136, DP_mult_209_n1135,
         DP_mult_209_n1134, DP_mult_209_n1133, DP_mult_209_n1132,
         DP_mult_209_n1131, DP_mult_209_n1130, DP_mult_209_n1129,
         DP_mult_209_n1128, DP_mult_209_n1127, DP_mult_209_n1126,
         DP_mult_209_n1125, DP_mult_209_n1124, DP_mult_209_n1123,
         DP_mult_209_n1122, DP_mult_209_n1121, DP_mult_209_n1120,
         DP_mult_209_n1119, DP_mult_209_n1118, DP_mult_209_n1117,
         DP_mult_209_n1116, DP_mult_209_n1115, DP_mult_209_n1114,
         DP_mult_209_n1113, DP_mult_209_n1112, DP_mult_209_n1111,
         DP_mult_209_n1110, DP_mult_209_n1109, DP_mult_209_n1108,
         DP_mult_209_n1107, DP_mult_209_n1106, DP_mult_209_n1105,
         DP_mult_209_n1104, DP_mult_209_n1103, DP_mult_209_n1102,
         DP_mult_209_n1101, DP_mult_209_n1100, DP_mult_209_n1099,
         DP_mult_209_n1098, DP_mult_209_n1097, DP_mult_209_n1096,
         DP_mult_209_n1095, DP_mult_209_n1094, DP_mult_209_n1093,
         DP_mult_209_n1092, DP_mult_209_n1091, DP_mult_209_n1090,
         DP_mult_209_n1089, DP_mult_209_n1088, DP_mult_209_n1087,
         DP_mult_209_n1086, DP_mult_209_n1085, DP_mult_209_n1084,
         DP_mult_209_n1083, DP_mult_209_n1082, DP_mult_209_n1081,
         DP_mult_209_n1080, DP_mult_209_n1079, DP_mult_209_n1078,
         DP_mult_209_n1077, DP_mult_209_n1076, DP_mult_209_n1075,
         DP_mult_209_n1074, DP_mult_209_n1073, DP_mult_209_n1072,
         DP_mult_209_n1071, DP_mult_209_n1070, DP_mult_209_n1069,
         DP_mult_209_n1068, DP_mult_209_n1067, DP_mult_209_n1066,
         DP_mult_209_n1065, DP_mult_209_n1064, DP_mult_209_n1063,
         DP_mult_209_n1062, DP_mult_209_n1061, DP_mult_209_n1060,
         DP_mult_209_n1059, DP_mult_209_n1058, DP_mult_209_n1057,
         DP_mult_209_n1056, DP_mult_209_n1055, DP_mult_209_n1054,
         DP_mult_209_n1053, DP_mult_209_n1052, DP_mult_209_n1051,
         DP_mult_209_n1050, DP_mult_209_n1049, DP_mult_209_n1048,
         DP_mult_209_n1047, DP_mult_209_n1046, DP_mult_209_n1045,
         DP_mult_209_n1044, DP_mult_209_n1043, DP_mult_209_n1042,
         DP_mult_209_n1041, DP_mult_209_n1040, DP_mult_209_n1039,
         DP_mult_209_n1038, DP_mult_209_n1037, DP_mult_209_n1036,
         DP_mult_209_n1035, DP_mult_209_n1034, DP_mult_209_n1033,
         DP_mult_209_n1032, DP_mult_209_n1031, DP_mult_209_n1030,
         DP_mult_209_n1029, DP_mult_209_n1028, DP_mult_209_n1027,
         DP_mult_209_n1026, DP_mult_209_n1025, DP_mult_209_n1024,
         DP_mult_209_n1023, DP_mult_209_n1022, DP_mult_209_n1021,
         DP_mult_209_n1020, DP_mult_209_n1019, DP_mult_209_n1018,
         DP_mult_209_n1017, DP_mult_209_n1016, DP_mult_209_n1015,
         DP_mult_209_n1014, DP_mult_209_n1013, DP_mult_209_n1012,
         DP_mult_209_n1011, DP_mult_209_n1010, DP_mult_209_n1009,
         DP_mult_209_n1008, DP_mult_209_n1007, DP_mult_209_n1006,
         DP_mult_209_n1005, DP_mult_209_n1004, DP_mult_209_n1003,
         DP_mult_209_n1002, DP_mult_209_n1001, DP_mult_209_n1000,
         DP_mult_209_n999, DP_mult_209_n998, DP_mult_209_n997,
         DP_mult_209_n996, DP_mult_209_n995, DP_mult_209_n994,
         DP_mult_209_n993, DP_mult_209_n992, DP_mult_209_n991,
         DP_mult_209_n990, DP_mult_209_n989, DP_mult_209_n988,
         DP_mult_209_n987, DP_mult_209_n986, DP_mult_209_n985,
         DP_mult_209_n984, DP_mult_209_n983, DP_mult_209_n982,
         DP_mult_209_n981, DP_mult_209_n980, DP_mult_209_n979,
         DP_mult_209_n978, DP_mult_209_n977, DP_mult_209_n976,
         DP_mult_209_n975, DP_mult_209_n974, DP_mult_209_n973,
         DP_mult_209_n972, DP_mult_209_n971, DP_mult_209_n970,
         DP_mult_209_n969, DP_mult_209_n968, DP_mult_209_n967,
         DP_mult_209_n966, DP_mult_209_n965, DP_mult_209_n964,
         DP_mult_209_n963, DP_mult_209_n962, DP_mult_209_n961,
         DP_mult_209_n960, DP_mult_209_n959, DP_mult_209_n958,
         DP_mult_209_n957, DP_mult_209_n956, DP_mult_209_n955,
         DP_mult_209_n954, DP_mult_209_n953, DP_mult_209_n952,
         DP_mult_209_n951, DP_mult_209_n950, DP_mult_209_n949,
         DP_mult_209_n948, DP_mult_209_n947, DP_mult_209_n946,
         DP_mult_209_n945, DP_mult_209_n944, DP_mult_209_n943,
         DP_mult_209_n942, DP_mult_209_n941, DP_mult_209_n940,
         DP_mult_209_n939, DP_mult_209_n938, DP_mult_209_n937,
         DP_mult_209_n936, DP_mult_209_n935, DP_mult_209_n934,
         DP_mult_209_n933, DP_mult_209_n932, DP_mult_209_n931,
         DP_mult_209_n930, DP_mult_209_n929, DP_mult_209_n928,
         DP_mult_209_n927, DP_mult_209_n926, DP_mult_209_n925,
         DP_mult_209_n924, DP_mult_209_n923, DP_mult_209_n922,
         DP_mult_209_n921, DP_mult_209_n920, DP_mult_209_n919,
         DP_mult_209_n918, DP_mult_209_n917, DP_mult_209_n916,
         DP_mult_209_n915, DP_mult_209_n914, DP_mult_209_n913,
         DP_mult_209_n912, DP_mult_209_n911, DP_mult_209_n910,
         DP_mult_209_n909, DP_mult_209_n908, DP_mult_209_n907,
         DP_mult_209_n906, DP_mult_209_n905, DP_mult_209_n904,
         DP_mult_209_n903, DP_mult_209_n902, DP_mult_209_n901,
         DP_mult_209_n900, DP_mult_209_n899, DP_mult_209_n898,
         DP_mult_209_n897, DP_mult_209_n896, DP_mult_209_n895,
         DP_mult_209_n894, DP_mult_209_n893, DP_mult_209_n892,
         DP_mult_209_n891, DP_mult_209_n890, DP_mult_209_n889,
         DP_mult_209_n888, DP_mult_209_n887, DP_mult_209_n886,
         DP_mult_209_n885, DP_mult_209_n884, DP_mult_209_n883,
         DP_mult_209_n882, DP_mult_209_n881, DP_mult_209_n880,
         DP_mult_209_n879, DP_mult_209_n878, DP_mult_209_n877,
         DP_mult_209_n876, DP_mult_209_n875, DP_mult_209_n874,
         DP_mult_209_n873, DP_mult_209_n872, DP_mult_209_n871,
         DP_mult_209_n870, DP_mult_209_n869, DP_mult_209_n868,
         DP_mult_209_n867, DP_mult_209_n866, DP_mult_209_n865,
         DP_mult_209_n864, DP_mult_209_n863, DP_mult_209_n862,
         DP_mult_209_n861, DP_mult_209_n860, DP_mult_209_n859,
         DP_mult_209_n858, DP_mult_209_n857, DP_mult_209_n856,
         DP_mult_209_n855, DP_mult_209_n854, DP_mult_209_n853,
         DP_mult_209_n852, DP_mult_209_n851, DP_mult_209_n850,
         DP_mult_209_n849, DP_mult_209_n848, DP_mult_209_n847,
         DP_mult_209_n846, DP_mult_209_n845, DP_mult_209_n844,
         DP_mult_209_n843, DP_mult_209_n841, DP_mult_209_n840,
         DP_mult_209_n839, DP_mult_209_n838, DP_mult_209_n837,
         DP_mult_209_n836, DP_mult_209_n835, DP_mult_209_n834,
         DP_mult_209_n833, DP_mult_209_n832, DP_mult_209_n831,
         DP_mult_209_n830, DP_mult_209_n829, DP_mult_209_n828,
         DP_mult_209_n827, DP_mult_209_n826, DP_mult_209_n825,
         DP_mult_209_n824, DP_mult_209_n823, DP_mult_209_n822,
         DP_mult_209_n821, DP_mult_209_n820, DP_mult_209_n819,
         DP_mult_209_n818, DP_mult_209_n817, DP_mult_209_n816,
         DP_mult_209_n815, DP_mult_209_n814, DP_mult_209_n813,
         DP_mult_209_n812, DP_mult_209_n811, DP_mult_209_n810,
         DP_mult_209_n809, DP_mult_209_n808, DP_mult_209_n807,
         DP_mult_209_n806, DP_mult_209_n805, DP_mult_209_n804,
         DP_mult_209_n803, DP_mult_209_n802, DP_mult_209_n801,
         DP_mult_209_n800, DP_mult_209_n799, DP_mult_209_n798,
         DP_mult_209_n797, DP_mult_209_n796, DP_mult_209_n795,
         DP_mult_209_n794, DP_mult_209_n793, DP_mult_209_n792,
         DP_mult_209_n791, DP_mult_209_n790, DP_mult_209_n789,
         DP_mult_209_n788, DP_mult_209_n787, DP_mult_209_n786,
         DP_mult_209_n785, DP_mult_209_n784, DP_mult_209_n783,
         DP_mult_209_n782, DP_mult_209_n781, DP_mult_209_n780,
         DP_mult_209_n779, DP_mult_209_n778, DP_mult_209_n777,
         DP_mult_209_n776, DP_mult_209_n775, DP_mult_209_n774,
         DP_mult_209_n773, DP_mult_209_n772, DP_mult_209_n771,
         DP_mult_209_n770, DP_mult_209_n769, DP_mult_209_n768,
         DP_mult_209_n767, DP_mult_209_n766, DP_mult_209_n765,
         DP_mult_209_n764, DP_mult_209_n763, DP_mult_209_n762,
         DP_mult_209_n761, DP_mult_209_n760, DP_mult_209_n759,
         DP_mult_209_n758, DP_mult_209_n757, DP_mult_209_n756,
         DP_mult_209_n755, DP_mult_209_n754, DP_mult_209_n753,
         DP_mult_209_n752, DP_mult_209_n751, DP_mult_209_n750,
         DP_mult_209_n749, DP_mult_209_n748, DP_mult_209_n747,
         DP_mult_209_n746, DP_mult_209_n745, DP_mult_209_n744,
         DP_mult_209_n743, DP_mult_209_n742, DP_mult_209_n741,
         DP_mult_209_n740, DP_mult_209_n739, DP_mult_209_n738,
         DP_mult_209_n737, DP_mult_209_n736, DP_mult_209_n735,
         DP_mult_209_n734, DP_mult_209_n733, DP_mult_209_n732,
         DP_mult_209_n731, DP_mult_209_n730, DP_mult_209_n729,
         DP_mult_209_n728, DP_mult_209_n727, DP_mult_209_n726,
         DP_mult_209_n725, DP_mult_209_n724, DP_mult_209_n723,
         DP_mult_209_n722, DP_mult_209_n721, DP_mult_209_n720,
         DP_mult_209_n719, DP_mult_209_n718, DP_mult_209_n717,
         DP_mult_209_n716, DP_mult_209_n715, DP_mult_209_n714,
         DP_mult_209_n713, DP_mult_209_n712, DP_mult_209_n711,
         DP_mult_209_n710, DP_mult_209_n709, DP_mult_209_n708,
         DP_mult_209_n707, DP_mult_209_n706, DP_mult_209_n705,
         DP_mult_209_n704, DP_mult_209_n703, DP_mult_209_n702,
         DP_mult_209_n701, DP_mult_209_n700, DP_mult_209_n699,
         DP_mult_209_n698, DP_mult_209_n697, DP_mult_209_n696,
         DP_mult_209_n695, DP_mult_209_n694, DP_mult_209_n693,
         DP_mult_209_n692, DP_mult_209_n691, DP_mult_209_n690,
         DP_mult_209_n689, DP_mult_209_n688, DP_mult_209_n687,
         DP_mult_209_n686, DP_mult_209_n685, DP_mult_209_n684,
         DP_mult_209_n683, DP_mult_209_n682, DP_mult_209_n681,
         DP_mult_209_n680, DP_mult_209_n679, DP_mult_209_n678,
         DP_mult_209_n677, DP_mult_209_n676, DP_mult_209_n675,
         DP_mult_209_n673, DP_mult_209_n671, DP_mult_209_n668,
         DP_mult_209_n667, DP_mult_209_n666, DP_mult_209_n663,
         DP_mult_209_n662, DP_mult_209_n661, DP_mult_209_n657,
         DP_mult_209_n646, DP_mult_209_n645, DP_mult_209_n644,
         DP_mult_209_n643, DP_mult_209_n638, DP_mult_209_n637,
         DP_mult_209_n636, DP_mult_209_n635, DP_mult_209_n634,
         DP_mult_209_n633, DP_mult_209_n632, DP_mult_209_n631,
         DP_mult_209_n630, DP_mult_209_n629, DP_mult_209_n628,
         DP_mult_209_n627, DP_mult_209_n626, DP_mult_209_n625,
         DP_mult_209_n620, DP_mult_209_n611, DP_mult_209_n610,
         DP_mult_209_n609, DP_mult_209_n600, DP_mult_209_n599,
         DP_mult_209_n598, DP_mult_209_n597, DP_mult_209_n596,
         DP_mult_209_n595, DP_mult_209_n594, DP_mult_209_n593,
         DP_mult_209_n592, DP_mult_209_n591, DP_mult_209_n590,
         DP_mult_209_n589, DP_mult_209_n588, DP_mult_209_n583,
         DP_mult_209_n582, DP_mult_209_n581, DP_mult_209_n572,
         DP_mult_209_n571, DP_mult_209_n570, DP_mult_209_n569,
         DP_mult_209_n568, DP_mult_209_n567, DP_mult_209_n566,
         DP_mult_209_n565, DP_mult_209_n564, DP_mult_209_n563,
         DP_mult_209_n562, DP_mult_209_n561, DP_mult_209_n560,
         DP_mult_209_n559, DP_mult_209_n558, DP_mult_209_n553,
         DP_mult_209_n552, DP_mult_209_n551, DP_mult_209_n550,
         DP_mult_209_n547, DP_mult_209_n546, DP_mult_209_n545,
         DP_mult_209_n544, DP_mult_209_n543, DP_mult_209_n542,
         DP_mult_209_n541, DP_mult_209_n540, DP_mult_209_n539,
         DP_mult_209_n538, DP_mult_209_n537, DP_mult_209_n536,
         DP_mult_209_n535, DP_mult_209_n534, DP_mult_209_n533,
         DP_mult_209_n532, DP_mult_209_n531, DP_mult_209_n526,
         DP_mult_209_n525, DP_mult_209_n524, DP_mult_209_n522,
         DP_mult_209_n521, DP_mult_209_n520, DP_mult_209_n519,
         DP_mult_209_n517, DP_mult_209_n516, DP_mult_209_n515,
         DP_mult_209_n514, DP_mult_209_n513, DP_mult_209_n512,
         DP_mult_209_n511, DP_mult_209_n508, DP_mult_209_n506,
         DP_mult_209_n505, DP_mult_209_n504, DP_mult_209_n503,
         DP_mult_209_n502, DP_mult_209_n501, DP_mult_209_n499,
         DP_mult_209_n498, DP_mult_209_n497, DP_mult_209_n496,
         DP_mult_209_n495, DP_mult_209_n492, DP_mult_209_n490,
         DP_mult_209_n489, DP_mult_209_n488, DP_mult_209_n487,
         DP_mult_209_n486, DP_mult_209_n483, DP_mult_209_n481,
         DP_mult_209_n480, DP_mult_209_n479, DP_mult_209_n478,
         DP_mult_209_n477, DP_mult_209_n476, DP_mult_209_n475,
         DP_mult_209_n474, DP_mult_209_n468, DP_mult_209_n467,
         DP_mult_209_n466, DP_mult_209_n465, DP_mult_209_n464,
         DP_mult_209_n463, DP_mult_209_n462, DP_mult_209_n461,
         DP_mult_209_n459, DP_mult_209_n457, DP_mult_209_n456,
         DP_mult_209_n455, DP_mult_209_n454, DP_mult_209_n453,
         DP_mult_209_n452, DP_mult_209_n451, DP_mult_209_n448,
         DP_mult_209_n445, DP_mult_209_n439, DP_mult_209_n438,
         DP_mult_209_n437, DP_mult_209_n436, DP_mult_209_n435,
         DP_mult_209_n434, DP_mult_209_n432, DP_mult_209_n431,
         DP_mult_209_n430, DP_mult_209_n429, DP_mult_209_n428,
         DP_mult_209_n427, DP_mult_209_n426, DP_mult_209_n423,
         DP_mult_209_n422, DP_mult_209_n421, DP_mult_209_n420,
         DP_mult_209_n419, DP_mult_209_n418, DP_mult_209_n416,
         DP_mult_209_n412, DP_mult_209_n411, DP_mult_209_n410,
         DP_mult_209_n409, DP_mult_209_n407, DP_mult_209_n405,
         DP_mult_209_n402, DP_mult_209_n401, DP_mult_209_n400,
         DP_mult_209_n399, DP_mult_209_n398, DP_mult_209_n397,
         DP_mult_209_n396, DP_mult_209_n394, DP_mult_209_n390,
         DP_mult_209_n389, DP_mult_209_n388, DP_mult_209_n387,
         DP_mult_209_n384, DP_mult_209_n383, DP_mult_209_n382,
         DP_mult_209_n381, DP_mult_209_n380, DP_mult_209_n379,
         DP_mult_209_n378, DP_mult_209_n376, DP_mult_209_n372,
         DP_mult_209_n371, DP_mult_209_n370, DP_mult_209_n369,
         DP_mult_209_n367, DP_mult_209_n365, DP_mult_209_n364,
         DP_mult_209_n363, DP_mult_209_n362, DP_mult_209_n361,
         DP_mult_209_n360, DP_mult_209_n359, DP_mult_209_n356,
         DP_mult_209_n355, DP_mult_209_n354, DP_mult_209_n353,
         DP_mult_209_n352, DP_mult_209_n350, DP_mult_209_n348,
         DP_mult_209_n347, DP_mult_209_n346, DP_mult_209_n345,
         DP_mult_209_n344, DP_mult_209_n343, DP_mult_209_n342,
         DP_mult_209_n341, DP_mult_209_n339, DP_mult_209_n337,
         DP_mult_209_n336, DP_mult_209_n335, DP_mult_209_n334,
         DP_mult_209_n333, DP_mult_209_n332, DP_mult_209_n327,
         DP_mult_209_n326, DP_mult_209_n325, DP_mult_209_n320,
         DP_mult_209_n319, DP_mult_209_n318, DP_mult_209_n317,
         DP_mult_209_n316, DP_mult_209_n315, DP_mult_209_n314,
         DP_mult_209_n313, DP_mult_209_n312, DP_mult_209_n311,
         DP_mult_209_n310, DP_mult_209_n309, DP_mult_209_n308,
         DP_mult_209_n307, DP_mult_209_n306, DP_mult_209_n305,
         DP_mult_209_n304, DP_mult_209_n303, DP_mult_209_n302,
         DP_mult_209_n301, DP_mult_209_n297, DP_mult_209_n283,
         DP_mult_209_n279, DP_mult_209_n277, DP_mult_209_n267,
         DP_mult_209_n259, DP_mult_209_n251, CU_n3, CU_n2, CU_n1,
         CU_nextState_0_, reg_delay_0_n6, reg_delay_0_n5, reg_delay_1_n4,
         reg_delay_1_n3;
  wire   [0:10] DP_y_out;
  wire   [0:23] DP_pipe13;
  wire   [0:23] DP_pipe0_coeff_pipe03;
  wire   [0:23] DP_pipe12;
  wire   [0:23] DP_pipe0_coeff_pipe02;
  wire   [0:23] DP_pipe11;
  wire   [0:23] DP_pipe0_coeff_pipe01;
  wire   [0:23] DP_pipe10;
  wire   [0:23] DP_pipe0_coeff_pipe00;
  wire   [0:23] DP_pipe03;
  wire   [0:23] DP_pipe02;
  wire   [0:23] DP_pipe01;
  wire   [0:23] DP_pipe00;
  wire   [0:23] DP_ret1;
  wire   [0:23] DP_sw1_coeff_ret1;
  wire   [0:23] DP_ret0;
  wire   [0:23] DP_sw0_coeff_ret0;
  wire   [0:23] DP_sw2;
  wire   [95:0] DP_coeffs_ff_int;
  wire   [47:0] DP_coeffs_fb_int;

  OAI21_X1 DP_U39 ( .B1(DP_n1), .B2(DP_n26), .A(DP_n25), .ZN(DP_y_out[10]) );
  INV_X1 DP_U38 ( .A(DP_y_10_), .ZN(DP_n26) );
  OAI21_X1 DP_U37 ( .B1(DP_n1), .B2(DP_n24), .A(DP_n25), .ZN(DP_y_out[9]) );
  INV_X1 DP_U36 ( .A(DP_y_9_), .ZN(DP_n24) );
  OAI21_X1 DP_U35 ( .B1(DP_n1), .B2(DP_n23), .A(DP_n25), .ZN(DP_y_out[8]) );
  INV_X1 DP_U34 ( .A(DP_y_8_), .ZN(DP_n23) );
  OAI21_X1 DP_U33 ( .B1(DP_n1), .B2(DP_n22), .A(DP_n25), .ZN(DP_y_out[7]) );
  INV_X1 DP_U32 ( .A(DP_y_7_), .ZN(DP_n22) );
  OAI21_X1 DP_U31 ( .B1(DP_n1), .B2(DP_n21), .A(DP_n25), .ZN(DP_y_out[6]) );
  INV_X1 DP_U30 ( .A(DP_y_6_), .ZN(DP_n21) );
  OAI21_X1 DP_U29 ( .B1(DP_n1), .B2(DP_n20), .A(DP_n25), .ZN(DP_y_out[5]) );
  INV_X1 DP_U28 ( .A(DP_y_5_), .ZN(DP_n20) );
  OAI21_X1 DP_U27 ( .B1(DP_n1), .B2(DP_n19), .A(DP_n25), .ZN(DP_y_out[4]) );
  INV_X1 DP_U26 ( .A(DP_y_4_), .ZN(DP_n19) );
  OAI21_X1 DP_U25 ( .B1(DP_n1), .B2(DP_n18), .A(DP_n25), .ZN(DP_y_out[3]) );
  INV_X1 DP_U24 ( .A(DP_y_3_), .ZN(DP_n18) );
  OAI21_X1 DP_U23 ( .B1(DP_n1), .B2(DP_n17), .A(DP_n25), .ZN(DP_y_out[2]) );
  INV_X1 DP_U22 ( .A(DP_y_2_), .ZN(DP_n17) );
  OAI21_X1 DP_U21 ( .B1(DP_n1), .B2(DP_n16), .A(DP_n25), .ZN(DP_y_out[1]) );
  INV_X1 DP_U20 ( .A(DP_y_1_), .ZN(DP_n16) );
  OAI21_X1 DP_U19 ( .B1(DP_n1), .B2(DP_n15), .A(DP_n25), .ZN(DP_y_out[0]) );
  INV_X1 DP_U18 ( .A(DP_y_23), .ZN(DP_n14) );
  INV_X1 DP_U17 ( .A(DP_y_0_), .ZN(DP_n15) );
  INV_X1 DP_U16 ( .A(DP_y_11_), .ZN(DP_n13) );
  BUF_X1 DP_U15 ( .A(rst_n), .Z(DP_n2) );
  BUF_X1 DP_U14 ( .A(DP_n2), .Z(DP_n6) );
  BUF_X1 DP_U13 ( .A(DP_n2), .Z(DP_n7) );
  BUF_X1 DP_U12 ( .A(DP_n2), .Z(DP_n8) );
  BUF_X1 DP_U11 ( .A(DP_n3), .Z(DP_n9) );
  BUF_X1 DP_U10 ( .A(DP_n3), .Z(DP_n11) );
  BUF_X1 DP_U9 ( .A(DP_n3), .Z(DP_n12) );
  BUF_X1 DP_U8 ( .A(DP_n2), .Z(DP_n4) );
  CLKBUF_X2 DP_U7 ( .A(DP_n2), .Z(DP_n5) );
  AND2_X2 DP_U6 ( .A1(DP_y_23), .A2(DP_n13), .ZN(DP_n1) );
  NAND2_X2 DP_U5 ( .A1(DP_n14), .A2(DP_y_11_), .ZN(DP_n25) );
  BUF_X1 DP_U4 ( .A(rst_n), .Z(DP_n3) );
  BUF_X2 DP_U3 ( .A(DP_n3), .Z(DP_n10) );
  MUX2_X1 DP_reg_in_U14 ( .A(DP_x_11_), .B(dIn[11]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n36) );
  MUX2_X1 DP_reg_in_U13 ( .A(DP_x_10_), .B(dIn[10]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n35) );
  MUX2_X1 DP_reg_in_U12 ( .A(DP_x_9_), .B(dIn[9]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n34) );
  MUX2_X1 DP_reg_in_U11 ( .A(DP_x_8_), .B(dIn[8]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n33) );
  MUX2_X1 DP_reg_in_U10 ( .A(DP_x_7_), .B(dIn[7]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n32) );
  MUX2_X1 DP_reg_in_U9 ( .A(DP_x_6_), .B(dIn[6]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n31) );
  MUX2_X1 DP_reg_in_U8 ( .A(DP_x_5_), .B(dIn[5]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n30) );
  MUX2_X1 DP_reg_in_U7 ( .A(DP_x_4_), .B(dIn[4]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n29) );
  MUX2_X1 DP_reg_in_U6 ( .A(DP_x_3_), .B(dIn[3]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n28) );
  MUX2_X1 DP_reg_in_U5 ( .A(DP_x_2_), .B(dIn[2]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n27) );
  MUX2_X1 DP_reg_in_U4 ( .A(DP_x_1_), .B(dIn[1]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n26) );
  MUX2_X1 DP_reg_in_U3 ( .A(DP_x_0_), .B(dIn[0]), .S(DP_reg_in_n13), .Z(
        DP_reg_in_n25) );
  BUF_X1 DP_reg_in_U2 ( .A(vIn), .Z(DP_reg_in_n13) );
  DFFR_X1 DP_reg_in_Q_reg_0_ ( .D(DP_reg_in_n25), .CK(clk), .RN(DP_n5), .Q(
        DP_x_0_) );
  DFFR_X1 DP_reg_in_Q_reg_1_ ( .D(DP_reg_in_n26), .CK(clk), .RN(DP_n5), .Q(
        DP_x_1_) );
  DFFR_X1 DP_reg_in_Q_reg_2_ ( .D(DP_reg_in_n27), .CK(clk), .RN(DP_n5), .Q(
        DP_x_2_) );
  DFFR_X1 DP_reg_in_Q_reg_3_ ( .D(DP_reg_in_n28), .CK(clk), .RN(DP_n5), .Q(
        DP_x_3_) );
  DFFR_X1 DP_reg_in_Q_reg_4_ ( .D(DP_reg_in_n29), .CK(clk), .RN(DP_n5), .Q(
        DP_x_4_) );
  DFFR_X1 DP_reg_in_Q_reg_5_ ( .D(DP_reg_in_n30), .CK(clk), .RN(DP_n5), .Q(
        DP_x_5_) );
  DFFR_X1 DP_reg_in_Q_reg_6_ ( .D(DP_reg_in_n31), .CK(clk), .RN(DP_n5), .Q(
        DP_x_6_) );
  DFFR_X1 DP_reg_in_Q_reg_7_ ( .D(DP_reg_in_n32), .CK(clk), .RN(DP_n5), .Q(
        DP_x_7_) );
  DFFR_X1 DP_reg_in_Q_reg_8_ ( .D(DP_reg_in_n33), .CK(clk), .RN(DP_n5), .Q(
        DP_x_8_) );
  DFFR_X1 DP_reg_in_Q_reg_9_ ( .D(DP_reg_in_n34), .CK(clk), .RN(DP_n5), .Q(
        DP_x_9_) );
  DFFR_X1 DP_reg_in_Q_reg_10_ ( .D(DP_reg_in_n35), .CK(clk), .RN(DP_n5), .Q(
        DP_x_10_) );
  DFFR_X1 DP_reg_in_Q_reg_11_ ( .D(DP_reg_in_n36), .CK(clk), .RN(DP_n5), .Q(
        DP_x_11_) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U49 ( .A(DP_reg_coeff_fb_i_1_n73), .B(
        coeffs_fb[47]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n72) );
  INV_X1 DP_reg_coeff_fb_i_1_U48 ( .A(DP_reg_coeff_fb_i_1_n48), .ZN(
        DP_reg_coeff_fb_i_1_n73) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U47 ( .A(DP_reg_coeff_fb_i_1_n39), .B(
        coeffs_fb[46]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n71) );
  INV_X1 DP_reg_coeff_fb_i_1_U46 ( .A(DP_reg_coeff_fb_i_1_n47), .ZN(
        DP_reg_coeff_fb_i_1_n39) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U45 ( .A(DP_reg_coeff_fb_i_1_n74), .B(
        coeffs_fb[45]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n70) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U44 ( .A(DP_reg_coeff_fb_i_1_n75), .B(
        coeffs_fb[44]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n69) );
  INV_X1 DP_reg_coeff_fb_i_1_U43 ( .A(DP_reg_coeff_fb_i_1_n45), .ZN(
        DP_coeffs_fb_int[3]) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U42 ( .A(DP_reg_coeff_fb_i_1_n76), .B(
        coeffs_fb[43]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n68) );
  INV_X1 DP_reg_coeff_fb_i_1_U41 ( .A(DP_reg_coeff_fb_i_1_n44), .ZN(
        DP_coeffs_fb_int[4]) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U40 ( .A(DP_reg_coeff_fb_i_1_n28), .B(
        coeffs_fb[42]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n67) );
  INV_X1 DP_reg_coeff_fb_i_1_U39 ( .A(DP_reg_coeff_fb_i_1_n43), .ZN(
        DP_reg_coeff_fb_i_1_n28) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U38 ( .A(DP_reg_coeff_fb_i_1_n77), .B(
        coeffs_fb[41]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n66) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U37 ( .A(DP_reg_coeff_fb_i_1_n26), .B(
        coeffs_fb[40]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n65) );
  INV_X1 DP_reg_coeff_fb_i_1_U36 ( .A(DP_reg_coeff_fb_i_1_n41), .ZN(
        DP_reg_coeff_fb_i_1_n26) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U35 ( .A(DP_reg_coeff_fb_i_1_n25), .B(
        coeffs_fb[39]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n64) );
  INV_X1 DP_reg_coeff_fb_i_1_U34 ( .A(DP_reg_coeff_fb_i_1_n40), .ZN(
        DP_reg_coeff_fb_i_1_n25) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U33 ( .A(DP_coeffs_fb_int[9]), .B(coeffs_fb[38]), 
        .S(DP_reg_coeff_fb_i_1_n14), .Z(DP_reg_coeff_fb_i_1_n63) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U32 ( .A(DP_reg_coeff_fb_i_1_n78), .B(
        coeffs_fb[37]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n62) );
  INV_X1 DP_reg_coeff_fb_i_1_U31 ( .A(DP_reg_coeff_fb_i_1_n38), .ZN(
        DP_coeffs_fb_int[10]) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U30 ( .A(DP_reg_coeff_fb_i_1_n23), .B(
        coeffs_fb[36]), .S(DP_reg_coeff_fb_i_1_n14), .Z(
        DP_reg_coeff_fb_i_1_n61) );
  INV_X1 DP_reg_coeff_fb_i_1_U29 ( .A(DP_reg_coeff_fb_i_1_n37), .ZN(
        DP_reg_coeff_fb_i_1_n23) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U28 ( .A(DP_reg_coeff_fb_i_1_n79), .B(
        coeffs_fb[35]), .S(DP_reg_coeff_fb_i_1_n13), .Z(
        DP_reg_coeff_fb_i_1_n60) );
  INV_X1 DP_reg_coeff_fb_i_1_U27 ( .A(DP_reg_coeff_fb_i_1_n36), .ZN(
        DP_coeffs_fb_int[12]) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U26 ( .A(DP_coeffs_fb_int[13]), .B(coeffs_fb[34]), .S(DP_reg_coeff_fb_i_1_n13), .Z(DP_reg_coeff_fb_i_1_n59) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U25 ( .A(DP_reg_coeff_fb_i_1_n21), .B(
        coeffs_fb[33]), .S(DP_reg_coeff_fb_i_1_n13), .Z(
        DP_reg_coeff_fb_i_1_n58) );
  INV_X1 DP_reg_coeff_fb_i_1_U24 ( .A(DP_reg_coeff_fb_i_1_n34), .ZN(
        DP_reg_coeff_fb_i_1_n21) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U23 ( .A(DP_coeffs_fb_int[15]), .B(coeffs_fb[32]), .S(DP_reg_coeff_fb_i_1_n13), .Z(DP_reg_coeff_fb_i_1_n57) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U22 ( .A(DP_reg_coeff_fb_i_1_n80), .B(
        coeffs_fb[31]), .S(DP_reg_coeff_fb_i_1_n13), .Z(
        DP_reg_coeff_fb_i_1_n56) );
  INV_X1 DP_reg_coeff_fb_i_1_U21 ( .A(DP_reg_coeff_fb_i_1_n32), .ZN(
        DP_coeffs_fb_int[16]) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U20 ( .A(DP_reg_coeff_fb_i_1_n81), .B(
        coeffs_fb[30]), .S(DP_reg_coeff_fb_i_1_n13), .Z(
        DP_reg_coeff_fb_i_1_n55) );
  INV_X1 DP_reg_coeff_fb_i_1_U19 ( .A(DP_reg_coeff_fb_i_1_n31), .ZN(
        DP_coeffs_fb_int[17]) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U18 ( .A(DP_reg_coeff_fb_i_1_n82), .B(
        coeffs_fb[29]), .S(DP_reg_coeff_fb_i_1_n13), .Z(
        DP_reg_coeff_fb_i_1_n54) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U17 ( .A(DP_reg_coeff_fb_i_1_n18), .B(
        coeffs_fb[28]), .S(DP_reg_coeff_fb_i_1_n13), .Z(
        DP_reg_coeff_fb_i_1_n53) );
  INV_X1 DP_reg_coeff_fb_i_1_U16 ( .A(DP_reg_coeff_fb_i_1_n29), .ZN(
        DP_reg_coeff_fb_i_1_n18) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U15 ( .A(DP_coeffs_fb_int[20]), .B(coeffs_fb[27]), .S(DP_reg_coeff_fb_i_1_n13), .Z(DP_reg_coeff_fb_i_1_n52) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U14 ( .A(DP_coeffs_fb_int[21]), .B(coeffs_fb[26]), .S(DP_reg_coeff_fb_i_1_n13), .Z(DP_reg_coeff_fb_i_1_n51) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U13 ( .A(DP_reg_coeff_fb_i_1_n83), .B(
        coeffs_fb[25]), .S(DP_reg_coeff_fb_i_1_n13), .Z(
        DP_reg_coeff_fb_i_1_n50) );
  MUX2_X1 DP_reg_coeff_fb_i_1_U12 ( .A(DP_coeffs_fb_int[23]), .B(coeffs_fb[24]), .S(DP_reg_coeff_fb_i_1_n13), .Z(DP_reg_coeff_fb_i_1_n49) );
  BUF_X1 DP_reg_coeff_fb_i_1_U11 ( .A(vIn), .Z(DP_reg_coeff_fb_i_1_n14) );
  BUF_X1 DP_reg_coeff_fb_i_1_U10 ( .A(vIn), .Z(DP_reg_coeff_fb_i_1_n13) );
  BUF_X1 DP_reg_coeff_fb_i_1_U9 ( .A(DP_n4), .Z(DP_reg_coeff_fb_i_1_n15) );
  BUF_X1 DP_reg_coeff_fb_i_1_U8 ( .A(DP_n4), .Z(DP_reg_coeff_fb_i_1_n16) );
  INV_X1 DP_reg_coeff_fb_i_1_U5 ( .A(DP_reg_coeff_fb_i_1_n3), .ZN(
        DP_coeffs_fb_int[18]) );
  INV_X1 DP_reg_coeff_fb_i_1_U4 ( .A(DP_reg_coeff_fb_i_1_n42), .ZN(
        DP_coeffs_fb_int[6]) );
  INV_X2 DP_reg_coeff_fb_i_1_U3 ( .A(DP_reg_coeff_fb_i_1_n46), .ZN(
        DP_coeffs_fb_int[2]) );
  INV_X1 DP_reg_coeff_fb_i_1_U2 ( .A(DP_reg_coeff_fb_i_1_n1), .ZN(
        DP_coeffs_fb_int[22]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_2_ ( .D(DP_reg_coeff_fb_i_1_n51), .CK(clk), 
        .RN(DP_n4), .Q(DP_coeffs_fb_int[21]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_5_ ( .D(DP_reg_coeff_fb_i_1_n54), .CK(clk), 
        .RN(DP_n4), .Q(DP_reg_coeff_fb_i_1_n82), .QN(DP_reg_coeff_fb_i_1_n3)
         );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_3_ ( .D(DP_reg_coeff_fb_i_1_n52), .CK(clk), 
        .RN(DP_n4), .Q(DP_coeffs_fb_int[20]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_1_ ( .D(DP_reg_coeff_fb_i_1_n50), .CK(clk), 
        .RN(DP_n4), .Q(DP_reg_coeff_fb_i_1_n83), .QN(DP_reg_coeff_fb_i_1_n1)
         );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_0_ ( .D(DP_reg_coeff_fb_i_1_n49), .CK(clk), 
        .RN(DP_n4), .Q(DP_coeffs_fb_int[23]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_8_ ( .D(DP_reg_coeff_fb_i_1_n57), .CK(clk), 
        .RN(DP_n4), .Q(DP_coeffs_fb_int[15]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_10_ ( .D(DP_reg_coeff_fb_i_1_n59), .CK(clk), .RN(DP_n4), .Q(DP_coeffs_fb_int[13]) );
  SDFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_14_ ( .D(1'b0), .SI(
        DP_reg_coeff_fb_i_1_n63), .SE(1'b1), .CK(clk), .RN(
        DP_reg_coeff_fb_i_1_n15), .Q(DP_coeffs_fb_int[9]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_4_ ( .D(DP_reg_coeff_fb_i_1_n53), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_1_n16), .Q(DP_coeffs_fb_int[19]), .QN(
        DP_reg_coeff_fb_i_1_n29) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_6_ ( .D(DP_reg_coeff_fb_i_1_n55), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_1_n16), .Q(DP_reg_coeff_fb_i_1_n81), .QN(
        DP_reg_coeff_fb_i_1_n31) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_7_ ( .D(DP_reg_coeff_fb_i_1_n56), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_1_n16), .Q(DP_reg_coeff_fb_i_1_n80), .QN(
        DP_reg_coeff_fb_i_1_n32) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_9_ ( .D(DP_reg_coeff_fb_i_1_n58), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_1_n16), .Q(DP_coeffs_fb_int[14]), .QN(
        DP_reg_coeff_fb_i_1_n34) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_11_ ( .D(DP_reg_coeff_fb_i_1_n60), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n16), .Q(DP_reg_coeff_fb_i_1_n79), .QN(
        DP_reg_coeff_fb_i_1_n36) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_12_ ( .D(DP_reg_coeff_fb_i_1_n61), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_coeffs_fb_int[11]), .QN(
        DP_reg_coeff_fb_i_1_n37) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_13_ ( .D(DP_reg_coeff_fb_i_1_n62), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_reg_coeff_fb_i_1_n78), .QN(
        DP_reg_coeff_fb_i_1_n38) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_15_ ( .D(DP_reg_coeff_fb_i_1_n64), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_coeffs_fb_int[8]), .QN(
        DP_reg_coeff_fb_i_1_n40) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_16_ ( .D(DP_reg_coeff_fb_i_1_n65), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_coeffs_fb_int[7]), .QN(
        DP_reg_coeff_fb_i_1_n41) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_17_ ( .D(DP_reg_coeff_fb_i_1_n66), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_reg_coeff_fb_i_1_n77), .QN(
        DP_reg_coeff_fb_i_1_n42) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_18_ ( .D(DP_reg_coeff_fb_i_1_n67), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_coeffs_fb_int[5]), .QN(
        DP_reg_coeff_fb_i_1_n43) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_19_ ( .D(DP_reg_coeff_fb_i_1_n68), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_reg_coeff_fb_i_1_n76), .QN(
        DP_reg_coeff_fb_i_1_n44) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_20_ ( .D(DP_reg_coeff_fb_i_1_n69), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_reg_coeff_fb_i_1_n75), .QN(
        DP_reg_coeff_fb_i_1_n45) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_21_ ( .D(DP_reg_coeff_fb_i_1_n70), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_reg_coeff_fb_i_1_n74), .QN(
        DP_reg_coeff_fb_i_1_n46) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_22_ ( .D(DP_reg_coeff_fb_i_1_n71), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_coeffs_fb_int[1]), .QN(
        DP_reg_coeff_fb_i_1_n47) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_23_ ( .D(DP_reg_coeff_fb_i_1_n72), .CK(clk), .RN(DP_reg_coeff_fb_i_1_n15), .Q(DP_coeffs_fb_int[0]), .QN(
        DP_reg_coeff_fb_i_1_n48) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U55 ( .A(DP_reg_coeff_fb_i_2_n78), .B(
        coeffs_fb[23]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n79) );
  INV_X1 DP_reg_coeff_fb_i_2_U54 ( .A(DP_reg_coeff_fb_i_2_n103), .ZN(
        DP_reg_coeff_fb_i_2_n78) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U53 ( .A(DP_reg_coeff_fb_i_2_n77), .B(
        coeffs_fb[22]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n80) );
  INV_X1 DP_reg_coeff_fb_i_2_U52 ( .A(DP_reg_coeff_fb_i_2_n104), .ZN(
        DP_reg_coeff_fb_i_2_n77) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U51 ( .A(DP_reg_coeff_fb_i_2_n76), .B(
        coeffs_fb[21]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n81) );
  INV_X1 DP_reg_coeff_fb_i_2_U50 ( .A(DP_reg_coeff_fb_i_2_n105), .ZN(
        DP_reg_coeff_fb_i_2_n76) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U49 ( .A(DP_reg_coeff_fb_i_2_n75), .B(
        coeffs_fb[20]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n82) );
  INV_X1 DP_reg_coeff_fb_i_2_U48 ( .A(DP_reg_coeff_fb_i_2_n106), .ZN(
        DP_reg_coeff_fb_i_2_n75) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U47 ( .A(DP_reg_coeff_fb_i_2_n125), .B(
        coeffs_fb[19]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n83) );
  INV_X1 DP_reg_coeff_fb_i_2_U46 ( .A(DP_reg_coeff_fb_i_2_n107), .ZN(
        DP_coeffs_fb_int[28]) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U45 ( .A(DP_reg_coeff_fb_i_2_n73), .B(
        coeffs_fb[18]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n84) );
  INV_X1 DP_reg_coeff_fb_i_2_U44 ( .A(DP_reg_coeff_fb_i_2_n108), .ZN(
        DP_reg_coeff_fb_i_2_n73) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U43 ( .A(DP_coeffs_fb_int[30]), .B(coeffs_fb[17]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n85) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U42 ( .A(DP_reg_coeff_fb_i_2_n42), .B(
        coeffs_fb[16]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n86) );
  INV_X1 DP_reg_coeff_fb_i_2_U41 ( .A(DP_reg_coeff_fb_i_2_n109), .ZN(
        DP_reg_coeff_fb_i_2_n42) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U40 ( .A(DP_reg_coeff_fb_i_2_n28), .B(
        coeffs_fb[15]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n87) );
  INV_X1 DP_reg_coeff_fb_i_2_U39 ( .A(DP_reg_coeff_fb_i_2_n110), .ZN(
        DP_reg_coeff_fb_i_2_n28) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U38 ( .A(DP_reg_coeff_fb_i_2_n24), .B(
        coeffs_fb[14]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n88) );
  INV_X1 DP_reg_coeff_fb_i_2_U37 ( .A(DP_reg_coeff_fb_i_2_n111), .ZN(
        DP_reg_coeff_fb_i_2_n24) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U36 ( .A(DP_reg_coeff_fb_i_2_n126), .B(
        coeffs_fb[13]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n89) );
  INV_X1 DP_reg_coeff_fb_i_2_U35 ( .A(DP_reg_coeff_fb_i_2_n112), .ZN(
        DP_coeffs_fb_int[34]) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U34 ( .A(DP_reg_coeff_fb_i_2_n22), .B(
        coeffs_fb[12]), .S(DP_reg_coeff_fb_i_2_n8), .Z(DP_reg_coeff_fb_i_2_n90) );
  INV_X1 DP_reg_coeff_fb_i_2_U33 ( .A(DP_reg_coeff_fb_i_2_n113), .ZN(
        DP_reg_coeff_fb_i_2_n22) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U32 ( .A(DP_reg_coeff_fb_i_2_n21), .B(
        coeffs_fb[11]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n91) );
  INV_X1 DP_reg_coeff_fb_i_2_U31 ( .A(DP_reg_coeff_fb_i_2_n114), .ZN(
        DP_reg_coeff_fb_i_2_n21) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U30 ( .A(DP_reg_coeff_fb_i_2_n20), .B(
        coeffs_fb[10]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n92) );
  INV_X1 DP_reg_coeff_fb_i_2_U29 ( .A(DP_reg_coeff_fb_i_2_n115), .ZN(
        DP_reg_coeff_fb_i_2_n20) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U28 ( .A(DP_reg_coeff_fb_i_2_n19), .B(
        coeffs_fb[9]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n93)
         );
  INV_X1 DP_reg_coeff_fb_i_2_U27 ( .A(DP_reg_coeff_fb_i_2_n116), .ZN(
        DP_reg_coeff_fb_i_2_n19) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U26 ( .A(DP_reg_coeff_fb_i_2_n18), .B(
        coeffs_fb[8]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n94)
         );
  INV_X1 DP_reg_coeff_fb_i_2_U25 ( .A(DP_reg_coeff_fb_i_2_n117), .ZN(
        DP_reg_coeff_fb_i_2_n18) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U24 ( .A(DP_reg_coeff_fb_i_2_n17), .B(
        coeffs_fb[7]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n95)
         );
  INV_X1 DP_reg_coeff_fb_i_2_U23 ( .A(DP_reg_coeff_fb_i_2_n118), .ZN(
        DP_reg_coeff_fb_i_2_n17) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U22 ( .A(DP_reg_coeff_fb_i_2_n16), .B(
        coeffs_fb[6]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n96)
         );
  INV_X1 DP_reg_coeff_fb_i_2_U21 ( .A(DP_reg_coeff_fb_i_2_n119), .ZN(
        DP_reg_coeff_fb_i_2_n16) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U20 ( .A(DP_reg_coeff_fb_i_2_n15), .B(
        coeffs_fb[5]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n97)
         );
  INV_X1 DP_reg_coeff_fb_i_2_U19 ( .A(DP_reg_coeff_fb_i_2_n120), .ZN(
        DP_reg_coeff_fb_i_2_n15) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U18 ( .A(DP_reg_coeff_fb_i_2_n14), .B(
        coeffs_fb[4]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n98)
         );
  INV_X1 DP_reg_coeff_fb_i_2_U17 ( .A(DP_reg_coeff_fb_i_2_n121), .ZN(
        DP_reg_coeff_fb_i_2_n14) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U16 ( .A(DP_coeffs_fb_int[44]), .B(coeffs_fb[3]), 
        .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n99) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U15 ( .A(DP_coeffs_fb_int[45]), .B(coeffs_fb[2]), 
        .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n100) );
  INV_X1 DP_reg_coeff_fb_i_2_U14 ( .A(DP_reg_coeff_fb_i_2_n122), .ZN(
        DP_coeffs_fb_int[45]) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U13 ( .A(DP_reg_coeff_fb_i_2_n12), .B(
        coeffs_fb[1]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n101) );
  INV_X1 DP_reg_coeff_fb_i_2_U12 ( .A(DP_reg_coeff_fb_i_2_n123), .ZN(
        DP_reg_coeff_fb_i_2_n12) );
  MUX2_X1 DP_reg_coeff_fb_i_2_U11 ( .A(DP_reg_coeff_fb_i_2_n11), .B(
        coeffs_fb[0]), .S(DP_reg_coeff_fb_i_2_n7), .Z(DP_reg_coeff_fb_i_2_n102) );
  INV_X1 DP_reg_coeff_fb_i_2_U10 ( .A(DP_reg_coeff_fb_i_2_n124), .ZN(
        DP_reg_coeff_fb_i_2_n11) );
  BUF_X1 DP_reg_coeff_fb_i_2_U9 ( .A(vIn), .Z(DP_reg_coeff_fb_i_2_n8) );
  BUF_X1 DP_reg_coeff_fb_i_2_U8 ( .A(vIn), .Z(DP_reg_coeff_fb_i_2_n7) );
  BUF_X1 DP_reg_coeff_fb_i_2_U7 ( .A(DP_n8), .Z(DP_reg_coeff_fb_i_2_n9) );
  BUF_X1 DP_reg_coeff_fb_i_2_U6 ( .A(DP_n8), .Z(DP_reg_coeff_fb_i_2_n10) );
  SDFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_17_ ( .D(1'b0), .SI(
        DP_reg_coeff_fb_i_2_n85), .SE(1'b1), .CK(clk), .RN(
        DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[30]) );
  SDFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_3_ ( .D(1'b0), .SI(
        DP_reg_coeff_fb_i_2_n99), .SE(1'b1), .CK(clk), .RN(
        DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[44]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_0_ ( .D(DP_reg_coeff_fb_i_2_n102), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[47]), .QN(
        DP_reg_coeff_fb_i_2_n124) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_1_ ( .D(DP_reg_coeff_fb_i_2_n101), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[46]), .QN(
        DP_reg_coeff_fb_i_2_n123) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_2_ ( .D(DP_reg_coeff_fb_i_2_n100), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n10), .QN(DP_reg_coeff_fb_i_2_n122) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_4_ ( .D(DP_reg_coeff_fb_i_2_n98), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[43]), .QN(
        DP_reg_coeff_fb_i_2_n121) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_5_ ( .D(DP_reg_coeff_fb_i_2_n97), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[42]), .QN(
        DP_reg_coeff_fb_i_2_n120) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_6_ ( .D(DP_reg_coeff_fb_i_2_n96), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[41]), .QN(
        DP_reg_coeff_fb_i_2_n119) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_7_ ( .D(DP_reg_coeff_fb_i_2_n95), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[40]), .QN(
        DP_reg_coeff_fb_i_2_n118) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_8_ ( .D(DP_reg_coeff_fb_i_2_n94), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[39]), .QN(
        DP_reg_coeff_fb_i_2_n117) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_9_ ( .D(DP_reg_coeff_fb_i_2_n93), .CK(clk), 
        .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[38]), .QN(
        DP_reg_coeff_fb_i_2_n116) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_10_ ( .D(DP_reg_coeff_fb_i_2_n92), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[37]), .QN(
        DP_reg_coeff_fb_i_2_n115) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_11_ ( .D(DP_reg_coeff_fb_i_2_n91), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n10), .Q(DP_coeffs_fb_int[36]), .QN(
        DP_reg_coeff_fb_i_2_n114) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_12_ ( .D(DP_reg_coeff_fb_i_2_n90), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[35]), .QN(
        DP_reg_coeff_fb_i_2_n113) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_13_ ( .D(DP_reg_coeff_fb_i_2_n89), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_reg_coeff_fb_i_2_n126), .QN(
        DP_reg_coeff_fb_i_2_n112) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_14_ ( .D(DP_reg_coeff_fb_i_2_n88), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[33]), .QN(
        DP_reg_coeff_fb_i_2_n111) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_15_ ( .D(DP_reg_coeff_fb_i_2_n87), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[32]), .QN(
        DP_reg_coeff_fb_i_2_n110) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_16_ ( .D(DP_reg_coeff_fb_i_2_n86), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[31]), .QN(
        DP_reg_coeff_fb_i_2_n109) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_18_ ( .D(DP_reg_coeff_fb_i_2_n84), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[29]), .QN(
        DP_reg_coeff_fb_i_2_n108) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_19_ ( .D(DP_reg_coeff_fb_i_2_n83), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_reg_coeff_fb_i_2_n125), .QN(
        DP_reg_coeff_fb_i_2_n107) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_20_ ( .D(DP_reg_coeff_fb_i_2_n82), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[27]), .QN(
        DP_reg_coeff_fb_i_2_n106) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_21_ ( .D(DP_reg_coeff_fb_i_2_n81), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[26]), .QN(
        DP_reg_coeff_fb_i_2_n105) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_22_ ( .D(DP_reg_coeff_fb_i_2_n80), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[25]), .QN(
        DP_reg_coeff_fb_i_2_n104) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_23_ ( .D(DP_reg_coeff_fb_i_2_n79), .CK(clk), .RN(DP_reg_coeff_fb_i_2_n9), .Q(DP_coeffs_fb_int[24]), .QN(
        DP_reg_coeff_fb_i_2_n103) );
  MUX2_X1 DP_reg_b_i_0_U53 ( .A(DP_reg_b_i_0_n77), .B(coeffs_ff[95]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n78) );
  INV_X1 DP_reg_b_i_0_U52 ( .A(DP_reg_b_i_0_n102), .ZN(DP_reg_b_i_0_n77) );
  MUX2_X1 DP_reg_b_i_0_U51 ( .A(DP_reg_b_i_0_n125), .B(coeffs_ff[94]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n79) );
  INV_X1 DP_reg_b_i_0_U50 ( .A(DP_reg_b_i_0_n103), .ZN(DP_coeffs_ff_int[1]) );
  MUX2_X1 DP_reg_b_i_0_U49 ( .A(DP_reg_b_i_0_n126), .B(coeffs_ff[93]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n80) );
  MUX2_X1 DP_reg_b_i_0_U48 ( .A(DP_reg_b_i_0_n3), .B(coeffs_ff[92]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n81) );
  INV_X1 DP_reg_b_i_0_U47 ( .A(DP_reg_b_i_0_n105), .ZN(DP_coeffs_ff_int[3]) );
  MUX2_X1 DP_reg_b_i_0_U46 ( .A(DP_reg_b_i_0_n73), .B(coeffs_ff[91]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n82) );
  INV_X1 DP_reg_b_i_0_U45 ( .A(DP_reg_b_i_0_n106), .ZN(DP_reg_b_i_0_n73) );
  MUX2_X1 DP_reg_b_i_0_U44 ( .A(DP_reg_b_i_0_n28), .B(coeffs_ff[90]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n83) );
  INV_X1 DP_reg_b_i_0_U43 ( .A(DP_reg_b_i_0_n107), .ZN(DP_reg_b_i_0_n28) );
  MUX2_X1 DP_reg_b_i_0_U42 ( .A(DP_reg_b_i_0_n127), .B(coeffs_ff[89]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n84) );
  INV_X1 DP_reg_b_i_0_U41 ( .A(DP_reg_b_i_0_n108), .ZN(DP_coeffs_ff_int[6]) );
  MUX2_X1 DP_reg_b_i_0_U40 ( .A(DP_reg_b_i_0_n23), .B(coeffs_ff[88]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n85) );
  INV_X1 DP_reg_b_i_0_U39 ( .A(DP_reg_b_i_0_n109), .ZN(DP_reg_b_i_0_n23) );
  MUX2_X1 DP_reg_b_i_0_U38 ( .A(DP_reg_b_i_0_n22), .B(coeffs_ff[87]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n86) );
  INV_X1 DP_reg_b_i_0_U37 ( .A(DP_reg_b_i_0_n110), .ZN(DP_reg_b_i_0_n22) );
  MUX2_X1 DP_reg_b_i_0_U36 ( .A(DP_reg_b_i_0_n21), .B(coeffs_ff[86]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n87) );
  INV_X1 DP_reg_b_i_0_U35 ( .A(DP_reg_b_i_0_n111), .ZN(DP_reg_b_i_0_n21) );
  MUX2_X1 DP_reg_b_i_0_U34 ( .A(DP_reg_b_i_0_n128), .B(coeffs_ff[85]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n88) );
  MUX2_X1 DP_reg_b_i_0_U33 ( .A(DP_reg_b_i_0_n19), .B(coeffs_ff[84]), .S(
        DP_reg_b_i_0_n5), .Z(DP_reg_b_i_0_n89) );
  INV_X1 DP_reg_b_i_0_U32 ( .A(DP_reg_b_i_0_n113), .ZN(DP_reg_b_i_0_n19) );
  MUX2_X1 DP_reg_b_i_0_U31 ( .A(DP_reg_b_i_0_n129), .B(coeffs_ff[83]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n90) );
  MUX2_X1 DP_reg_b_i_0_U30 ( .A(DP_reg_b_i_0_n17), .B(coeffs_ff[82]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n91) );
  INV_X1 DP_reg_b_i_0_U29 ( .A(DP_reg_b_i_0_n115), .ZN(DP_reg_b_i_0_n17) );
  MUX2_X1 DP_reg_b_i_0_U28 ( .A(DP_reg_b_i_0_n130), .B(coeffs_ff[81]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n92) );
  INV_X1 DP_reg_b_i_0_U27 ( .A(DP_reg_b_i_0_n116), .ZN(DP_coeffs_ff_int[14])
         );
  MUX2_X1 DP_reg_b_i_0_U26 ( .A(DP_reg_b_i_0_n15), .B(coeffs_ff[80]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n93) );
  INV_X1 DP_reg_b_i_0_U25 ( .A(DP_reg_b_i_0_n117), .ZN(DP_reg_b_i_0_n15) );
  MUX2_X1 DP_reg_b_i_0_U24 ( .A(DP_reg_b_i_0_n14), .B(coeffs_ff[79]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n94) );
  INV_X1 DP_reg_b_i_0_U23 ( .A(DP_reg_b_i_0_n118), .ZN(DP_reg_b_i_0_n14) );
  MUX2_X1 DP_reg_b_i_0_U22 ( .A(DP_reg_b_i_0_n13), .B(coeffs_ff[78]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n95) );
  INV_X1 DP_reg_b_i_0_U21 ( .A(DP_reg_b_i_0_n119), .ZN(DP_reg_b_i_0_n13) );
  MUX2_X1 DP_reg_b_i_0_U20 ( .A(DP_reg_b_i_0_n12), .B(coeffs_ff[77]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n96) );
  INV_X1 DP_reg_b_i_0_U19 ( .A(DP_reg_b_i_0_n120), .ZN(DP_reg_b_i_0_n12) );
  MUX2_X1 DP_reg_b_i_0_U18 ( .A(DP_reg_b_i_0_n11), .B(coeffs_ff[76]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n97) );
  INV_X1 DP_reg_b_i_0_U17 ( .A(DP_reg_b_i_0_n121), .ZN(DP_reg_b_i_0_n11) );
  MUX2_X1 DP_reg_b_i_0_U16 ( .A(DP_reg_b_i_0_n131), .B(coeffs_ff[75]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n98) );
  MUX2_X1 DP_reg_b_i_0_U15 ( .A(DP_reg_b_i_0_n10), .B(coeffs_ff[74]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n99) );
  INV_X1 DP_reg_b_i_0_U14 ( .A(DP_reg_b_i_0_n122), .ZN(DP_reg_b_i_0_n10) );
  MUX2_X1 DP_reg_b_i_0_U13 ( .A(DP_reg_b_i_0_n9), .B(coeffs_ff[73]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n100) );
  INV_X1 DP_reg_b_i_0_U12 ( .A(DP_reg_b_i_0_n123), .ZN(DP_reg_b_i_0_n9) );
  MUX2_X1 DP_reg_b_i_0_U11 ( .A(DP_reg_b_i_0_n8), .B(coeffs_ff[72]), .S(
        DP_reg_b_i_0_n4), .Z(DP_reg_b_i_0_n101) );
  INV_X1 DP_reg_b_i_0_U10 ( .A(DP_reg_b_i_0_n124), .ZN(DP_reg_b_i_0_n8) );
  BUF_X1 DP_reg_b_i_0_U9 ( .A(vIn), .Z(DP_reg_b_i_0_n5) );
  BUF_X1 DP_reg_b_i_0_U8 ( .A(vIn), .Z(DP_reg_b_i_0_n4) );
  BUF_X1 DP_reg_b_i_0_U7 ( .A(rst_n), .Z(DP_reg_b_i_0_n6) );
  BUF_X1 DP_reg_b_i_0_U6 ( .A(rst_n), .Z(DP_reg_b_i_0_n7) );
  INV_X2 DP_reg_b_i_0_U5 ( .A(DP_reg_b_i_0_n112), .ZN(DP_coeffs_ff_int[10]) );
  INV_X1 DP_reg_b_i_0_U4 ( .A(DP_reg_b_i_0_n1), .ZN(DP_coeffs_ff_int[20]) );
  INV_X1 DP_reg_b_i_0_U3 ( .A(DP_reg_b_i_0_n114), .ZN(DP_coeffs_ff_int[12]) );
  INV_X1 DP_reg_b_i_0_U2 ( .A(DP_reg_b_i_0_n104), .ZN(DP_coeffs_ff_int[2]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_3_ ( .D(DP_reg_b_i_0_n98), .CK(clk), .RN(rst_n), 
        .Q(DP_reg_b_i_0_n131), .QN(DP_reg_b_i_0_n1) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_0_ ( .D(DP_reg_b_i_0_n101), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[23]), .QN(DP_reg_b_i_0_n124) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_1_ ( .D(DP_reg_b_i_0_n100), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[22]), .QN(DP_reg_b_i_0_n123) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_2_ ( .D(DP_reg_b_i_0_n99), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[21]), .QN(DP_reg_b_i_0_n122) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_4_ ( .D(DP_reg_b_i_0_n97), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[19]), .QN(DP_reg_b_i_0_n121) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_5_ ( .D(DP_reg_b_i_0_n96), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[18]), .QN(DP_reg_b_i_0_n120) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_6_ ( .D(DP_reg_b_i_0_n95), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[17]), .QN(DP_reg_b_i_0_n119) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_7_ ( .D(DP_reg_b_i_0_n94), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[16]), .QN(DP_reg_b_i_0_n118) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_8_ ( .D(DP_reg_b_i_0_n93), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[15]), .QN(DP_reg_b_i_0_n117) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_9_ ( .D(DP_reg_b_i_0_n92), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_reg_b_i_0_n130), .QN(DP_reg_b_i_0_n116) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_10_ ( .D(DP_reg_b_i_0_n91), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_coeffs_ff_int[13]), .QN(DP_reg_b_i_0_n115) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_11_ ( .D(DP_reg_b_i_0_n90), .CK(clk), .RN(
        DP_reg_b_i_0_n7), .Q(DP_reg_b_i_0_n129), .QN(DP_reg_b_i_0_n114) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_12_ ( .D(DP_reg_b_i_0_n89), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_coeffs_ff_int[11]), .QN(DP_reg_b_i_0_n113) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_13_ ( .D(DP_reg_b_i_0_n88), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_reg_b_i_0_n128), .QN(DP_reg_b_i_0_n112) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_14_ ( .D(DP_reg_b_i_0_n87), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_coeffs_ff_int[9]), .QN(DP_reg_b_i_0_n111) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_15_ ( .D(DP_reg_b_i_0_n86), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_coeffs_ff_int[8]), .QN(DP_reg_b_i_0_n110) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_16_ ( .D(DP_reg_b_i_0_n85), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_coeffs_ff_int[7]), .QN(DP_reg_b_i_0_n109) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_17_ ( .D(DP_reg_b_i_0_n84), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_reg_b_i_0_n127), .QN(DP_reg_b_i_0_n108) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_18_ ( .D(DP_reg_b_i_0_n83), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_coeffs_ff_int[5]), .QN(DP_reg_b_i_0_n107) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_19_ ( .D(DP_reg_b_i_0_n82), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_coeffs_ff_int[4]), .QN(DP_reg_b_i_0_n106) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_20_ ( .D(DP_reg_b_i_0_n81), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_reg_b_i_0_n3), .QN(DP_reg_b_i_0_n105) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_21_ ( .D(DP_reg_b_i_0_n80), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_reg_b_i_0_n126), .QN(DP_reg_b_i_0_n104) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_22_ ( .D(DP_reg_b_i_0_n79), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_reg_b_i_0_n125), .QN(DP_reg_b_i_0_n103) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_23_ ( .D(DP_reg_b_i_0_n78), .CK(clk), .RN(
        DP_reg_b_i_0_n6), .Q(DP_coeffs_ff_int[0]), .QN(DP_reg_b_i_0_n102) );
  MUX2_X1 DP_reg_b_i_1_U55 ( .A(DP_reg_b_i_1_n78), .B(coeffs_ff[71]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n79) );
  INV_X1 DP_reg_b_i_1_U54 ( .A(DP_reg_b_i_1_n103), .ZN(DP_reg_b_i_1_n78) );
  MUX2_X1 DP_reg_b_i_1_U53 ( .A(DP_reg_b_i_1_n77), .B(coeffs_ff[70]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n80) );
  INV_X1 DP_reg_b_i_1_U52 ( .A(DP_reg_b_i_1_n104), .ZN(DP_reg_b_i_1_n77) );
  MUX2_X1 DP_reg_b_i_1_U51 ( .A(DP_reg_b_i_1_n125), .B(coeffs_ff[69]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n81) );
  INV_X1 DP_reg_b_i_1_U50 ( .A(DP_reg_b_i_1_n105), .ZN(DP_coeffs_ff_int[26])
         );
  MUX2_X1 DP_reg_b_i_1_U49 ( .A(DP_reg_b_i_1_n75), .B(coeffs_ff[68]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n82) );
  INV_X1 DP_reg_b_i_1_U48 ( .A(DP_reg_b_i_1_n106), .ZN(DP_reg_b_i_1_n75) );
  MUX2_X1 DP_reg_b_i_1_U47 ( .A(DP_reg_b_i_1_n74), .B(coeffs_ff[67]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n83) );
  INV_X1 DP_reg_b_i_1_U46 ( .A(DP_reg_b_i_1_n107), .ZN(DP_reg_b_i_1_n74) );
  MUX2_X1 DP_reg_b_i_1_U45 ( .A(DP_reg_b_i_1_n73), .B(coeffs_ff[66]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n84) );
  INV_X1 DP_reg_b_i_1_U44 ( .A(DP_reg_b_i_1_n108), .ZN(DP_reg_b_i_1_n73) );
  MUX2_X1 DP_reg_b_i_1_U43 ( .A(DP_coeffs_ff_int[30]), .B(coeffs_ff[65]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n85) );
  MUX2_X1 DP_reg_b_i_1_U42 ( .A(DP_reg_b_i_1_n42), .B(coeffs_ff[64]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n86) );
  INV_X1 DP_reg_b_i_1_U41 ( .A(DP_reg_b_i_1_n109), .ZN(DP_reg_b_i_1_n42) );
  MUX2_X1 DP_reg_b_i_1_U40 ( .A(DP_reg_b_i_1_n126), .B(coeffs_ff[63]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n87) );
  INV_X1 DP_reg_b_i_1_U39 ( .A(DP_reg_b_i_1_n110), .ZN(DP_coeffs_ff_int[32])
         );
  MUX2_X1 DP_reg_b_i_1_U38 ( .A(DP_reg_b_i_1_n24), .B(coeffs_ff[62]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n88) );
  INV_X1 DP_reg_b_i_1_U37 ( .A(DP_reg_b_i_1_n111), .ZN(DP_reg_b_i_1_n24) );
  MUX2_X1 DP_reg_b_i_1_U36 ( .A(DP_reg_b_i_1_n23), .B(coeffs_ff[61]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n89) );
  INV_X1 DP_reg_b_i_1_U35 ( .A(DP_reg_b_i_1_n112), .ZN(DP_reg_b_i_1_n23) );
  MUX2_X1 DP_reg_b_i_1_U34 ( .A(DP_reg_b_i_1_n22), .B(coeffs_ff[60]), .S(
        DP_reg_b_i_1_n8), .Z(DP_reg_b_i_1_n90) );
  INV_X1 DP_reg_b_i_1_U33 ( .A(DP_reg_b_i_1_n113), .ZN(DP_reg_b_i_1_n22) );
  MUX2_X1 DP_reg_b_i_1_U32 ( .A(DP_reg_b_i_1_n127), .B(coeffs_ff[59]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n91) );
  INV_X1 DP_reg_b_i_1_U31 ( .A(DP_reg_b_i_1_n114), .ZN(DP_coeffs_ff_int[36])
         );
  MUX2_X1 DP_reg_b_i_1_U30 ( .A(DP_reg_b_i_1_n20), .B(coeffs_ff[58]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n92) );
  INV_X1 DP_reg_b_i_1_U29 ( .A(DP_reg_b_i_1_n115), .ZN(DP_reg_b_i_1_n20) );
  MUX2_X1 DP_reg_b_i_1_U28 ( .A(DP_reg_b_i_1_n19), .B(coeffs_ff[57]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n93) );
  INV_X1 DP_reg_b_i_1_U27 ( .A(DP_reg_b_i_1_n116), .ZN(DP_reg_b_i_1_n19) );
  MUX2_X1 DP_reg_b_i_1_U26 ( .A(DP_reg_b_i_1_n18), .B(coeffs_ff[56]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n94) );
  INV_X1 DP_reg_b_i_1_U25 ( .A(DP_reg_b_i_1_n117), .ZN(DP_reg_b_i_1_n18) );
  MUX2_X1 DP_reg_b_i_1_U24 ( .A(DP_reg_b_i_1_n128), .B(coeffs_ff[55]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n95) );
  INV_X1 DP_reg_b_i_1_U23 ( .A(DP_reg_b_i_1_n118), .ZN(DP_coeffs_ff_int[40])
         );
  MUX2_X1 DP_reg_b_i_1_U22 ( .A(DP_reg_b_i_1_n16), .B(coeffs_ff[54]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n96) );
  INV_X1 DP_reg_b_i_1_U21 ( .A(DP_reg_b_i_1_n119), .ZN(DP_reg_b_i_1_n16) );
  MUX2_X1 DP_reg_b_i_1_U20 ( .A(DP_reg_b_i_1_n15), .B(coeffs_ff[53]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n97) );
  INV_X1 DP_reg_b_i_1_U19 ( .A(DP_reg_b_i_1_n120), .ZN(DP_reg_b_i_1_n15) );
  MUX2_X1 DP_reg_b_i_1_U18 ( .A(DP_reg_b_i_1_n14), .B(coeffs_ff[52]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n98) );
  INV_X1 DP_reg_b_i_1_U17 ( .A(DP_reg_b_i_1_n121), .ZN(DP_reg_b_i_1_n14) );
  MUX2_X1 DP_reg_b_i_1_U16 ( .A(DP_coeffs_ff_int[44]), .B(coeffs_ff[51]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n99) );
  MUX2_X1 DP_reg_b_i_1_U15 ( .A(DP_reg_b_i_1_n13), .B(coeffs_ff[50]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n100) );
  INV_X1 DP_reg_b_i_1_U14 ( .A(DP_reg_b_i_1_n122), .ZN(DP_reg_b_i_1_n13) );
  MUX2_X1 DP_reg_b_i_1_U13 ( .A(DP_reg_b_i_1_n12), .B(coeffs_ff[49]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n101) );
  INV_X1 DP_reg_b_i_1_U12 ( .A(DP_reg_b_i_1_n123), .ZN(DP_reg_b_i_1_n12) );
  MUX2_X1 DP_reg_b_i_1_U11 ( .A(DP_reg_b_i_1_n11), .B(coeffs_ff[48]), .S(
        DP_reg_b_i_1_n7), .Z(DP_reg_b_i_1_n102) );
  INV_X1 DP_reg_b_i_1_U10 ( .A(DP_reg_b_i_1_n124), .ZN(DP_reg_b_i_1_n11) );
  CLKBUF_X3 DP_reg_b_i_1_U9 ( .A(vIn), .Z(DP_reg_b_i_1_n7) );
  BUF_X1 DP_reg_b_i_1_U8 ( .A(vIn), .Z(DP_reg_b_i_1_n8) );
  BUF_X1 DP_reg_b_i_1_U7 ( .A(DP_n12), .Z(DP_reg_b_i_1_n9) );
  BUF_X1 DP_reg_b_i_1_U6 ( .A(DP_n12), .Z(DP_reg_b_i_1_n10) );
  SDFFR_X1 DP_reg_b_i_1_Q_reg_3_ ( .D(1'b0), .SI(DP_reg_b_i_1_n99), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[44]) );
  SDFFR_X1 DP_reg_b_i_1_Q_reg_17_ ( .D(1'b0), .SI(DP_reg_b_i_1_n85), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[30]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_0_ ( .D(DP_reg_b_i_1_n102), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[47]), .QN(DP_reg_b_i_1_n124) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_1_ ( .D(DP_reg_b_i_1_n101), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[46]), .QN(DP_reg_b_i_1_n123) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_2_ ( .D(DP_reg_b_i_1_n100), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[45]), .QN(DP_reg_b_i_1_n122) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_4_ ( .D(DP_reg_b_i_1_n98), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[43]), .QN(DP_reg_b_i_1_n121) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_5_ ( .D(DP_reg_b_i_1_n97), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[42]), .QN(DP_reg_b_i_1_n120) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_6_ ( .D(DP_reg_b_i_1_n96), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[41]), .QN(DP_reg_b_i_1_n119) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_7_ ( .D(DP_reg_b_i_1_n95), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_reg_b_i_1_n128), .QN(DP_reg_b_i_1_n118) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_8_ ( .D(DP_reg_b_i_1_n94), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[39]), .QN(DP_reg_b_i_1_n117) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_9_ ( .D(DP_reg_b_i_1_n93), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[38]), .QN(DP_reg_b_i_1_n116) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_10_ ( .D(DP_reg_b_i_1_n92), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_coeffs_ff_int[37]), .QN(DP_reg_b_i_1_n115) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_11_ ( .D(DP_reg_b_i_1_n91), .CK(clk), .RN(
        DP_reg_b_i_1_n10), .Q(DP_reg_b_i_1_n127), .QN(DP_reg_b_i_1_n114) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_12_ ( .D(DP_reg_b_i_1_n90), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[35]), .QN(DP_reg_b_i_1_n113) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_13_ ( .D(DP_reg_b_i_1_n89), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[34]), .QN(DP_reg_b_i_1_n112) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_14_ ( .D(DP_reg_b_i_1_n88), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[33]), .QN(DP_reg_b_i_1_n111) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_15_ ( .D(DP_reg_b_i_1_n87), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_reg_b_i_1_n126), .QN(DP_reg_b_i_1_n110) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_16_ ( .D(DP_reg_b_i_1_n86), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[31]), .QN(DP_reg_b_i_1_n109) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_18_ ( .D(DP_reg_b_i_1_n84), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[29]), .QN(DP_reg_b_i_1_n108) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_19_ ( .D(DP_reg_b_i_1_n83), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[28]), .QN(DP_reg_b_i_1_n107) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_20_ ( .D(DP_reg_b_i_1_n82), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[27]), .QN(DP_reg_b_i_1_n106) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_21_ ( .D(DP_reg_b_i_1_n81), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_reg_b_i_1_n125), .QN(DP_reg_b_i_1_n105) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_22_ ( .D(DP_reg_b_i_1_n80), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[25]), .QN(DP_reg_b_i_1_n104) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_23_ ( .D(DP_reg_b_i_1_n79), .CK(clk), .RN(
        DP_reg_b_i_1_n9), .Q(DP_coeffs_ff_int[24]), .QN(DP_reg_b_i_1_n103) );
  MUX2_X1 DP_reg_b_i_2_U53 ( .A(DP_reg_b_i_2_n76), .B(coeffs_ff[47]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n77) );
  INV_X1 DP_reg_b_i_2_U52 ( .A(DP_reg_b_i_2_n101), .ZN(DP_reg_b_i_2_n76) );
  MUX2_X1 DP_reg_b_i_2_U51 ( .A(DP_reg_b_i_2_n75), .B(coeffs_ff[46]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n78) );
  INV_X1 DP_reg_b_i_2_U50 ( .A(DP_reg_b_i_2_n102), .ZN(DP_reg_b_i_2_n75) );
  MUX2_X1 DP_reg_b_i_2_U49 ( .A(DP_reg_b_i_2_n74), .B(coeffs_ff[45]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n79) );
  INV_X1 DP_reg_b_i_2_U48 ( .A(DP_reg_b_i_2_n103), .ZN(DP_reg_b_i_2_n74) );
  MUX2_X1 DP_reg_b_i_2_U47 ( .A(DP_reg_b_i_2_n73), .B(coeffs_ff[44]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n80) );
  INV_X1 DP_reg_b_i_2_U46 ( .A(DP_reg_b_i_2_n104), .ZN(DP_reg_b_i_2_n73) );
  MUX2_X1 DP_reg_b_i_2_U45 ( .A(DP_reg_b_i_2_n124), .B(coeffs_ff[43]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n81) );
  MUX2_X1 DP_reg_b_i_2_U44 ( .A(DP_reg_b_i_2_n44), .B(coeffs_ff[42]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n82) );
  INV_X1 DP_reg_b_i_2_U43 ( .A(DP_reg_b_i_2_n105), .ZN(DP_reg_b_i_2_n44) );
  MUX2_X1 DP_reg_b_i_2_U42 ( .A(DP_reg_b_i_2_n125), .B(coeffs_ff[41]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n83) );
  MUX2_X1 DP_reg_b_i_2_U41 ( .A(DP_reg_b_i_2_n23), .B(coeffs_ff[40]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n84) );
  INV_X1 DP_reg_b_i_2_U40 ( .A(DP_reg_b_i_2_n107), .ZN(DP_reg_b_i_2_n23) );
  MUX2_X1 DP_reg_b_i_2_U39 ( .A(DP_reg_b_i_2_n22), .B(coeffs_ff[39]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n85) );
  INV_X1 DP_reg_b_i_2_U38 ( .A(DP_reg_b_i_2_n108), .ZN(DP_reg_b_i_2_n22) );
  MUX2_X1 DP_reg_b_i_2_U37 ( .A(DP_reg_b_i_2_n21), .B(coeffs_ff[38]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n86) );
  INV_X1 DP_reg_b_i_2_U36 ( .A(DP_reg_b_i_2_n109), .ZN(DP_reg_b_i_2_n21) );
  MUX2_X1 DP_reg_b_i_2_U35 ( .A(DP_reg_b_i_2_n126), .B(coeffs_ff[37]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n87) );
  INV_X1 DP_reg_b_i_2_U34 ( .A(DP_reg_b_i_2_n110), .ZN(DP_coeffs_ff_int[58])
         );
  MUX2_X1 DP_reg_b_i_2_U33 ( .A(DP_reg_b_i_2_n19), .B(coeffs_ff[36]), .S(
        DP_reg_b_i_2_n4), .Z(DP_reg_b_i_2_n88) );
  INV_X1 DP_reg_b_i_2_U32 ( .A(DP_reg_b_i_2_n111), .ZN(DP_reg_b_i_2_n19) );
  MUX2_X1 DP_reg_b_i_2_U31 ( .A(DP_reg_b_i_2_n18), .B(coeffs_ff[35]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n89) );
  INV_X1 DP_reg_b_i_2_U30 ( .A(DP_reg_b_i_2_n112), .ZN(DP_reg_b_i_2_n18) );
  MUX2_X1 DP_reg_b_i_2_U29 ( .A(DP_reg_b_i_2_n17), .B(coeffs_ff[34]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n90) );
  INV_X1 DP_reg_b_i_2_U28 ( .A(DP_reg_b_i_2_n113), .ZN(DP_reg_b_i_2_n17) );
  MUX2_X1 DP_reg_b_i_2_U27 ( .A(DP_reg_b_i_2_n127), .B(coeffs_ff[33]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n91) );
  INV_X1 DP_reg_b_i_2_U26 ( .A(DP_reg_b_i_2_n114), .ZN(DP_coeffs_ff_int[62])
         );
  MUX2_X1 DP_reg_b_i_2_U25 ( .A(DP_reg_b_i_2_n15), .B(coeffs_ff[32]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n92) );
  INV_X1 DP_reg_b_i_2_U24 ( .A(DP_reg_b_i_2_n115), .ZN(DP_reg_b_i_2_n15) );
  MUX2_X1 DP_reg_b_i_2_U23 ( .A(DP_reg_b_i_2_n128), .B(coeffs_ff[31]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n93) );
  INV_X1 DP_reg_b_i_2_U22 ( .A(DP_reg_b_i_2_n116), .ZN(DP_coeffs_ff_int[64])
         );
  MUX2_X1 DP_reg_b_i_2_U21 ( .A(DP_reg_b_i_2_n13), .B(coeffs_ff[30]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n94) );
  INV_X1 DP_reg_b_i_2_U20 ( .A(DP_reg_b_i_2_n117), .ZN(DP_reg_b_i_2_n13) );
  MUX2_X1 DP_reg_b_i_2_U19 ( .A(DP_reg_b_i_2_n129), .B(coeffs_ff[29]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n95) );
  INV_X1 DP_reg_b_i_2_U18 ( .A(DP_reg_b_i_2_n118), .ZN(DP_coeffs_ff_int[66])
         );
  MUX2_X1 DP_reg_b_i_2_U17 ( .A(DP_reg_b_i_2_n11), .B(coeffs_ff[28]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n96) );
  INV_X1 DP_reg_b_i_2_U16 ( .A(DP_reg_b_i_2_n119), .ZN(DP_reg_b_i_2_n11) );
  MUX2_X1 DP_reg_b_i_2_U15 ( .A(DP_reg_b_i_2_n130), .B(coeffs_ff[27]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n97) );
  INV_X1 DP_reg_b_i_2_U14 ( .A(DP_reg_b_i_2_n120), .ZN(DP_coeffs_ff_int[68])
         );
  MUX2_X1 DP_reg_b_i_2_U13 ( .A(DP_reg_b_i_2_n9), .B(coeffs_ff[26]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n98) );
  INV_X1 DP_reg_b_i_2_U12 ( .A(DP_reg_b_i_2_n121), .ZN(DP_reg_b_i_2_n9) );
  MUX2_X1 DP_reg_b_i_2_U11 ( .A(DP_reg_b_i_2_n8), .B(coeffs_ff[25]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n99) );
  INV_X1 DP_reg_b_i_2_U10 ( .A(DP_reg_b_i_2_n122), .ZN(DP_reg_b_i_2_n8) );
  MUX2_X1 DP_reg_b_i_2_U9 ( .A(DP_reg_b_i_2_n7), .B(coeffs_ff[24]), .S(
        DP_reg_b_i_2_n3), .Z(DP_reg_b_i_2_n100) );
  INV_X1 DP_reg_b_i_2_U8 ( .A(DP_reg_b_i_2_n123), .ZN(DP_reg_b_i_2_n7) );
  CLKBUF_X3 DP_reg_b_i_2_U7 ( .A(vIn), .Z(DP_reg_b_i_2_n3) );
  BUF_X1 DP_reg_b_i_2_U6 ( .A(vIn), .Z(DP_reg_b_i_2_n4) );
  BUF_X1 DP_reg_b_i_2_U5 ( .A(DP_n12), .Z(DP_reg_b_i_2_n5) );
  BUF_X1 DP_reg_b_i_2_U4 ( .A(DP_n12), .Z(DP_reg_b_i_2_n6) );
  INV_X1 DP_reg_b_i_2_U3 ( .A(DP_reg_b_i_2_n1), .ZN(DP_coeffs_ff_int[52]) );
  INV_X2 DP_reg_b_i_2_U2 ( .A(DP_reg_b_i_2_n106), .ZN(DP_coeffs_ff_int[54]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_19_ ( .D(DP_reg_b_i_2_n81), .CK(clk), .RN(DP_n12), 
        .Q(DP_reg_b_i_2_n124), .QN(DP_reg_b_i_2_n1) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_0_ ( .D(DP_reg_b_i_2_n100), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_coeffs_ff_int[71]), .QN(DP_reg_b_i_2_n123) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_1_ ( .D(DP_reg_b_i_2_n99), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_coeffs_ff_int[70]), .QN(DP_reg_b_i_2_n122) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_2_ ( .D(DP_reg_b_i_2_n98), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_coeffs_ff_int[69]), .QN(DP_reg_b_i_2_n121) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_3_ ( .D(DP_reg_b_i_2_n97), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_reg_b_i_2_n130), .QN(DP_reg_b_i_2_n120) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_4_ ( .D(DP_reg_b_i_2_n96), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_coeffs_ff_int[67]), .QN(DP_reg_b_i_2_n119) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_5_ ( .D(DP_reg_b_i_2_n95), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_reg_b_i_2_n129), .QN(DP_reg_b_i_2_n118) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_6_ ( .D(DP_reg_b_i_2_n94), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_coeffs_ff_int[65]), .QN(DP_reg_b_i_2_n117) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_7_ ( .D(DP_reg_b_i_2_n93), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_reg_b_i_2_n128), .QN(DP_reg_b_i_2_n116) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_8_ ( .D(DP_reg_b_i_2_n92), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_coeffs_ff_int[63]), .QN(DP_reg_b_i_2_n115) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_9_ ( .D(DP_reg_b_i_2_n91), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_reg_b_i_2_n127), .QN(DP_reg_b_i_2_n114) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_10_ ( .D(DP_reg_b_i_2_n90), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_coeffs_ff_int[61]), .QN(DP_reg_b_i_2_n113) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_11_ ( .D(DP_reg_b_i_2_n89), .CK(clk), .RN(
        DP_reg_b_i_2_n6), .Q(DP_coeffs_ff_int[60]), .QN(DP_reg_b_i_2_n112) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_12_ ( .D(DP_reg_b_i_2_n88), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[59]), .QN(DP_reg_b_i_2_n111) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_13_ ( .D(DP_reg_b_i_2_n87), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_reg_b_i_2_n126), .QN(DP_reg_b_i_2_n110) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_14_ ( .D(DP_reg_b_i_2_n86), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[57]), .QN(DP_reg_b_i_2_n109) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_15_ ( .D(DP_reg_b_i_2_n85), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[56]), .QN(DP_reg_b_i_2_n108) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_16_ ( .D(DP_reg_b_i_2_n84), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[55]), .QN(DP_reg_b_i_2_n107) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_17_ ( .D(DP_reg_b_i_2_n83), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_reg_b_i_2_n125), .QN(DP_reg_b_i_2_n106) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_18_ ( .D(DP_reg_b_i_2_n82), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[53]), .QN(DP_reg_b_i_2_n105) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_20_ ( .D(DP_reg_b_i_2_n80), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[51]), .QN(DP_reg_b_i_2_n104) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_21_ ( .D(DP_reg_b_i_2_n79), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[50]), .QN(DP_reg_b_i_2_n103) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_22_ ( .D(DP_reg_b_i_2_n78), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[49]), .QN(DP_reg_b_i_2_n102) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_23_ ( .D(DP_reg_b_i_2_n77), .CK(clk), .RN(
        DP_reg_b_i_2_n5), .Q(DP_coeffs_ff_int[48]), .QN(DP_reg_b_i_2_n101) );
  MUX2_X1 DP_reg_b_i_3_U55 ( .A(DP_reg_b_i_3_n78), .B(coeffs_ff[23]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n79) );
  INV_X1 DP_reg_b_i_3_U54 ( .A(DP_reg_b_i_3_n103), .ZN(DP_reg_b_i_3_n78) );
  MUX2_X1 DP_reg_b_i_3_U53 ( .A(DP_reg_b_i_3_n77), .B(coeffs_ff[22]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n80) );
  INV_X1 DP_reg_b_i_3_U52 ( .A(DP_reg_b_i_3_n104), .ZN(DP_reg_b_i_3_n77) );
  MUX2_X1 DP_reg_b_i_3_U51 ( .A(DP_reg_b_i_3_n126), .B(coeffs_ff[21]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n81) );
  INV_X1 DP_reg_b_i_3_U50 ( .A(DP_reg_b_i_3_n105), .ZN(DP_coeffs_ff_int[74])
         );
  MUX2_X1 DP_reg_b_i_3_U49 ( .A(DP_coeffs_ff_int[75]), .B(coeffs_ff[20]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n82) );
  INV_X1 DP_reg_b_i_3_U48 ( .A(DP_reg_b_i_3_n106), .ZN(DP_coeffs_ff_int[75])
         );
  MUX2_X1 DP_reg_b_i_3_U47 ( .A(DP_reg_b_i_3_n127), .B(coeffs_ff[19]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n83) );
  INV_X1 DP_reg_b_i_3_U46 ( .A(DP_reg_b_i_3_n107), .ZN(DP_coeffs_ff_int[76])
         );
  MUX2_X1 DP_reg_b_i_3_U45 ( .A(DP_reg_b_i_3_n73), .B(coeffs_ff[18]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n84) );
  INV_X1 DP_reg_b_i_3_U44 ( .A(DP_reg_b_i_3_n108), .ZN(DP_reg_b_i_3_n73) );
  MUX2_X1 DP_reg_b_i_3_U43 ( .A(DP_reg_b_i_3_n128), .B(coeffs_ff[17]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n85) );
  INV_X1 DP_reg_b_i_3_U42 ( .A(DP_reg_b_i_3_n109), .ZN(DP_coeffs_ff_int[78])
         );
  MUX2_X1 DP_reg_b_i_3_U41 ( .A(DP_reg_b_i_3_n24), .B(coeffs_ff[16]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n86) );
  INV_X1 DP_reg_b_i_3_U40 ( .A(DP_reg_b_i_3_n110), .ZN(DP_reg_b_i_3_n24) );
  MUX2_X1 DP_reg_b_i_3_U39 ( .A(DP_reg_b_i_3_n23), .B(coeffs_ff[15]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n87) );
  INV_X1 DP_reg_b_i_3_U38 ( .A(DP_reg_b_i_3_n111), .ZN(DP_reg_b_i_3_n23) );
  MUX2_X1 DP_reg_b_i_3_U37 ( .A(DP_reg_b_i_3_n22), .B(coeffs_ff[14]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n88) );
  INV_X1 DP_reg_b_i_3_U36 ( .A(DP_reg_b_i_3_n112), .ZN(DP_reg_b_i_3_n22) );
  MUX2_X1 DP_reg_b_i_3_U35 ( .A(DP_reg_b_i_3_n129), .B(coeffs_ff[13]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n89) );
  INV_X1 DP_reg_b_i_3_U34 ( .A(DP_reg_b_i_3_n113), .ZN(DP_coeffs_ff_int[82])
         );
  MUX2_X1 DP_reg_b_i_3_U33 ( .A(DP_reg_b_i_3_n20), .B(coeffs_ff[12]), .S(
        DP_reg_b_i_3_n6), .Z(DP_reg_b_i_3_n90) );
  INV_X1 DP_reg_b_i_3_U32 ( .A(DP_reg_b_i_3_n114), .ZN(DP_reg_b_i_3_n20) );
  MUX2_X1 DP_reg_b_i_3_U31 ( .A(DP_reg_b_i_3_n130), .B(coeffs_ff[11]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n91) );
  INV_X1 DP_reg_b_i_3_U30 ( .A(DP_reg_b_i_3_n115), .ZN(DP_coeffs_ff_int[84])
         );
  MUX2_X1 DP_reg_b_i_3_U29 ( .A(DP_reg_b_i_3_n18), .B(coeffs_ff[10]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n92) );
  INV_X1 DP_reg_b_i_3_U28 ( .A(DP_reg_b_i_3_n116), .ZN(DP_reg_b_i_3_n18) );
  MUX2_X1 DP_reg_b_i_3_U27 ( .A(DP_reg_b_i_3_n131), .B(coeffs_ff[9]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n93) );
  INV_X1 DP_reg_b_i_3_U26 ( .A(DP_reg_b_i_3_n117), .ZN(DP_coeffs_ff_int[86])
         );
  MUX2_X1 DP_reg_b_i_3_U25 ( .A(DP_reg_b_i_3_n16), .B(coeffs_ff[8]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n94) );
  INV_X1 DP_reg_b_i_3_U24 ( .A(DP_reg_b_i_3_n118), .ZN(DP_reg_b_i_3_n16) );
  MUX2_X1 DP_reg_b_i_3_U23 ( .A(DP_reg_b_i_3_n132), .B(coeffs_ff[7]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n95) );
  INV_X1 DP_reg_b_i_3_U22 ( .A(DP_reg_b_i_3_n119), .ZN(DP_coeffs_ff_int[88])
         );
  MUX2_X1 DP_reg_b_i_3_U21 ( .A(DP_reg_b_i_3_n14), .B(coeffs_ff[6]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n96) );
  INV_X1 DP_reg_b_i_3_U20 ( .A(DP_reg_b_i_3_n120), .ZN(DP_reg_b_i_3_n14) );
  MUX2_X1 DP_reg_b_i_3_U19 ( .A(DP_reg_b_i_3_n133), .B(coeffs_ff[5]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n97) );
  INV_X1 DP_reg_b_i_3_U18 ( .A(DP_reg_b_i_3_n121), .ZN(DP_coeffs_ff_int[90])
         );
  MUX2_X1 DP_reg_b_i_3_U17 ( .A(DP_reg_b_i_3_n12), .B(coeffs_ff[4]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n98) );
  INV_X1 DP_reg_b_i_3_U16 ( .A(DP_reg_b_i_3_n122), .ZN(DP_reg_b_i_3_n12) );
  MUX2_X1 DP_reg_b_i_3_U15 ( .A(DP_reg_b_i_3_n134), .B(coeffs_ff[3]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n99) );
  INV_X1 DP_reg_b_i_3_U14 ( .A(DP_reg_b_i_3_n123), .ZN(DP_coeffs_ff_int[92])
         );
  MUX2_X1 DP_reg_b_i_3_U13 ( .A(DP_reg_b_i_3_n10), .B(coeffs_ff[2]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n100) );
  INV_X1 DP_reg_b_i_3_U12 ( .A(DP_reg_b_i_3_n124), .ZN(DP_reg_b_i_3_n10) );
  MUX2_X1 DP_reg_b_i_3_U11 ( .A(DP_reg_b_i_3_n2), .B(coeffs_ff[1]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n101) );
  MUX2_X1 DP_reg_b_i_3_U10 ( .A(DP_reg_b_i_3_n9), .B(coeffs_ff[0]), .S(
        DP_reg_b_i_3_n5), .Z(DP_reg_b_i_3_n102) );
  INV_X1 DP_reg_b_i_3_U9 ( .A(DP_reg_b_i_3_n125), .ZN(DP_reg_b_i_3_n9) );
  BUF_X1 DP_reg_b_i_3_U8 ( .A(vIn), .Z(DP_reg_b_i_3_n6) );
  BUF_X1 DP_reg_b_i_3_U7 ( .A(vIn), .Z(DP_reg_b_i_3_n5) );
  BUF_X1 DP_reg_b_i_3_U6 ( .A(DP_n11), .Z(DP_reg_b_i_3_n7) );
  BUF_X1 DP_reg_b_i_3_U5 ( .A(DP_n11), .Z(DP_reg_b_i_3_n8) );
  INV_X1 DP_reg_b_i_3_U2 ( .A(DP_reg_b_i_3_n1), .ZN(DP_reg_b_i_3_n2) );
  SDFFR_X1 DP_reg_b_i_3_Q_reg_1_ ( .D(1'b0), .SI(DP_reg_b_i_3_n101), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_b_i_3_n8), .Q(DP_coeffs_ff_int[94]), .QN(
        DP_reg_b_i_3_n1) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_0_ ( .D(DP_reg_b_i_3_n102), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_coeffs_ff_int[95]), .QN(DP_reg_b_i_3_n125) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_2_ ( .D(DP_reg_b_i_3_n100), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_coeffs_ff_int[93]), .QN(DP_reg_b_i_3_n124) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_3_ ( .D(DP_reg_b_i_3_n99), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_reg_b_i_3_n134), .QN(DP_reg_b_i_3_n123) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_4_ ( .D(DP_reg_b_i_3_n98), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_coeffs_ff_int[91]), .QN(DP_reg_b_i_3_n122) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_5_ ( .D(DP_reg_b_i_3_n97), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_reg_b_i_3_n133), .QN(DP_reg_b_i_3_n121) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_6_ ( .D(DP_reg_b_i_3_n96), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_coeffs_ff_int[89]), .QN(DP_reg_b_i_3_n120) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_7_ ( .D(DP_reg_b_i_3_n95), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_reg_b_i_3_n132), .QN(DP_reg_b_i_3_n119) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_8_ ( .D(DP_reg_b_i_3_n94), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_coeffs_ff_int[87]), .QN(DP_reg_b_i_3_n118) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_9_ ( .D(DP_reg_b_i_3_n93), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_reg_b_i_3_n131), .QN(DP_reg_b_i_3_n117) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_10_ ( .D(DP_reg_b_i_3_n92), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_coeffs_ff_int[85]), .QN(DP_reg_b_i_3_n116) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_11_ ( .D(DP_reg_b_i_3_n91), .CK(clk), .RN(
        DP_reg_b_i_3_n8), .Q(DP_reg_b_i_3_n130), .QN(DP_reg_b_i_3_n115) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_12_ ( .D(DP_reg_b_i_3_n90), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_coeffs_ff_int[83]), .QN(DP_reg_b_i_3_n114) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_13_ ( .D(DP_reg_b_i_3_n89), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_reg_b_i_3_n129), .QN(DP_reg_b_i_3_n113) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_14_ ( .D(DP_reg_b_i_3_n88), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_coeffs_ff_int[81]), .QN(DP_reg_b_i_3_n112) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_15_ ( .D(DP_reg_b_i_3_n87), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_coeffs_ff_int[80]), .QN(DP_reg_b_i_3_n111) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_16_ ( .D(DP_reg_b_i_3_n86), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_coeffs_ff_int[79]), .QN(DP_reg_b_i_3_n110) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_17_ ( .D(DP_reg_b_i_3_n85), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_reg_b_i_3_n128), .QN(DP_reg_b_i_3_n109) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_18_ ( .D(DP_reg_b_i_3_n84), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_coeffs_ff_int[77]), .QN(DP_reg_b_i_3_n108) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_19_ ( .D(DP_reg_b_i_3_n83), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_reg_b_i_3_n127), .QN(DP_reg_b_i_3_n107) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_20_ ( .D(DP_reg_b_i_3_n82), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .QN(DP_reg_b_i_3_n106) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_21_ ( .D(DP_reg_b_i_3_n81), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_reg_b_i_3_n126), .QN(DP_reg_b_i_3_n105) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_22_ ( .D(DP_reg_b_i_3_n80), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_coeffs_ff_int[73]), .QN(DP_reg_b_i_3_n104) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_23_ ( .D(DP_reg_b_i_3_n79), .CK(clk), .RN(
        DP_reg_b_i_3_n7), .Q(DP_coeffs_ff_int[72]), .QN(DP_reg_b_i_3_n103) );
  MUX2_X1 DP_reg_sw0_U37 ( .A(DP_sw0_23_), .B(DP_w_23_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n41) );
  MUX2_X1 DP_reg_sw0_U36 ( .A(DP_sw0_22_), .B(DP_w_22_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n42) );
  MUX2_X1 DP_reg_sw0_U35 ( .A(DP_sw0_21_), .B(DP_w_21_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n43) );
  MUX2_X1 DP_reg_sw0_U34 ( .A(DP_sw0_20_), .B(DP_w_20_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n44) );
  MUX2_X1 DP_reg_sw0_U33 ( .A(DP_sw0_19_), .B(DP_w_19_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n45) );
  MUX2_X1 DP_reg_sw0_U32 ( .A(DP_sw0_18_), .B(DP_w_18_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n46) );
  MUX2_X1 DP_reg_sw0_U31 ( .A(DP_sw0_17_), .B(DP_w_17_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n47) );
  MUX2_X1 DP_reg_sw0_U30 ( .A(DP_sw0_16_), .B(DP_w_16_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n48) );
  MUX2_X1 DP_reg_sw0_U29 ( .A(DP_sw0_15_), .B(DP_w_15_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n65) );
  MUX2_X1 DP_reg_sw0_U28 ( .A(DP_sw0_14_), .B(DP_w_14_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n66) );
  MUX2_X1 DP_reg_sw0_U27 ( .A(DP_sw0_13_), .B(DP_w_13_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n67) );
  MUX2_X1 DP_reg_sw0_U26 ( .A(DP_reg_sw0_n22), .B(DP_w_12_), .S(DP_reg_sw0_n7), 
        .Z(DP_reg_sw0_n68) );
  INV_X1 DP_reg_sw0_U25 ( .A(DP_reg_sw0_n81), .ZN(DP_reg_sw0_n22) );
  MUX2_X1 DP_reg_sw0_U24 ( .A(DP_reg_sw0_n21), .B(DP_w_11_), .S(DP_reg_sw0_n6), 
        .Z(DP_reg_sw0_n69) );
  INV_X1 DP_reg_sw0_U23 ( .A(DP_reg_sw0_n82), .ZN(DP_reg_sw0_n21) );
  MUX2_X1 DP_reg_sw0_U22 ( .A(DP_sw0_10_), .B(DP_w_10_), .S(DP_reg_sw0_n6), 
        .Z(DP_reg_sw0_n70) );
  MUX2_X1 DP_reg_sw0_U21 ( .A(DP_reg_sw0_n19), .B(DP_w_9_), .S(DP_reg_sw0_n6), 
        .Z(DP_reg_sw0_n71) );
  INV_X1 DP_reg_sw0_U20 ( .A(DP_reg_sw0_n83), .ZN(DP_reg_sw0_n19) );
  MUX2_X1 DP_reg_sw0_U19 ( .A(DP_sw0_8_), .B(DP_w_8_), .S(DP_reg_sw0_n6), .Z(
        DP_reg_sw0_n72) );
  MUX2_X1 DP_reg_sw0_U18 ( .A(DP_reg_sw0_n17), .B(DP_w_7_), .S(DP_reg_sw0_n6), 
        .Z(DP_reg_sw0_n73) );
  INV_X1 DP_reg_sw0_U17 ( .A(DP_reg_sw0_n84), .ZN(DP_reg_sw0_n17) );
  MUX2_X1 DP_reg_sw0_U16 ( .A(DP_sw0_6_), .B(DP_w_6_), .S(DP_reg_sw0_n6), .Z(
        DP_reg_sw0_n74) );
  MUX2_X1 DP_reg_sw0_U15 ( .A(DP_reg_sw0_n15), .B(DP_w_5_), .S(DP_reg_sw0_n6), 
        .Z(DP_reg_sw0_n75) );
  INV_X1 DP_reg_sw0_U14 ( .A(DP_reg_sw0_n85), .ZN(DP_reg_sw0_n15) );
  MUX2_X1 DP_reg_sw0_U13 ( .A(DP_reg_sw0_n14), .B(DP_w_4_), .S(DP_reg_sw0_n6), 
        .Z(DP_reg_sw0_n76) );
  INV_X1 DP_reg_sw0_U12 ( .A(DP_reg_sw0_n86), .ZN(DP_reg_sw0_n14) );
  MUX2_X1 DP_reg_sw0_U11 ( .A(DP_sw0_3_), .B(DP_w_3_), .S(DP_reg_sw0_n6), .Z(
        DP_reg_sw0_n77) );
  MUX2_X1 DP_reg_sw0_U10 ( .A(DP_reg_sw0_n12), .B(DP_w_2_), .S(DP_reg_sw0_n6), 
        .Z(DP_reg_sw0_n78) );
  INV_X1 DP_reg_sw0_U9 ( .A(DP_reg_sw0_n87), .ZN(DP_reg_sw0_n12) );
  MUX2_X1 DP_reg_sw0_U8 ( .A(DP_sw0_1_), .B(DP_w_1_), .S(DP_reg_sw0_n6), .Z(
        DP_reg_sw0_n79) );
  MUX2_X1 DP_reg_sw0_U7 ( .A(DP_reg_sw0_n10), .B(DP_w_0_), .S(DP_reg_sw0_n6), 
        .Z(DP_reg_sw0_n80) );
  BUF_X1 DP_reg_sw0_U6 ( .A(DP_n11), .Z(DP_reg_sw0_n8) );
  BUF_X1 DP_reg_sw0_U5 ( .A(DP_n11), .Z(DP_reg_sw0_n9) );
  BUF_X1 DP_reg_sw0_U4 ( .A(sw_regs_en_int), .Z(DP_reg_sw0_n7) );
  BUF_X1 DP_reg_sw0_U3 ( .A(sw_regs_en_int), .Z(DP_reg_sw0_n6) );
  INV_X4 DP_reg_sw0_U2 ( .A(DP_reg_sw0_n3), .ZN(DP_sw0_0_) );
  DFFR_X2 DP_reg_sw0_Q_reg_22_ ( .D(DP_reg_sw0_n42), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_22_) );
  DFFR_X2 DP_reg_sw0_Q_reg_1_ ( .D(DP_reg_sw0_n79), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_1_) );
  DFFR_X1 DP_reg_sw0_Q_reg_0_ ( .D(DP_reg_sw0_n80), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_reg_sw0_n10), .QN(DP_reg_sw0_n3) );
  DFFR_X2 DP_reg_sw0_Q_reg_23_ ( .D(DP_reg_sw0_n41), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_23_) );
  DFFR_X1 DP_reg_sw0_Q_reg_2_ ( .D(DP_reg_sw0_n78), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_2_), .QN(DP_reg_sw0_n87) );
  DFFR_X1 DP_reg_sw0_Q_reg_3_ ( .D(DP_reg_sw0_n77), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_3_) );
  DFFR_X1 DP_reg_sw0_Q_reg_4_ ( .D(DP_reg_sw0_n76), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_4_), .QN(DP_reg_sw0_n86) );
  DFFR_X1 DP_reg_sw0_Q_reg_5_ ( .D(DP_reg_sw0_n75), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_5_), .QN(DP_reg_sw0_n85) );
  DFFR_X1 DP_reg_sw0_Q_reg_6_ ( .D(DP_reg_sw0_n74), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_6_) );
  DFFR_X1 DP_reg_sw0_Q_reg_7_ ( .D(DP_reg_sw0_n73), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_7_), .QN(DP_reg_sw0_n84) );
  DFFR_X1 DP_reg_sw0_Q_reg_8_ ( .D(DP_reg_sw0_n72), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_8_) );
  DFFR_X1 DP_reg_sw0_Q_reg_9_ ( .D(DP_reg_sw0_n71), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_9_), .QN(DP_reg_sw0_n83) );
  DFFR_X1 DP_reg_sw0_Q_reg_10_ ( .D(DP_reg_sw0_n70), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_10_) );
  DFFR_X1 DP_reg_sw0_Q_reg_11_ ( .D(DP_reg_sw0_n69), .CK(clk), .RN(
        DP_reg_sw0_n9), .Q(DP_sw0_11_), .QN(DP_reg_sw0_n82) );
  DFFR_X1 DP_reg_sw0_Q_reg_12_ ( .D(DP_reg_sw0_n68), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_12_), .QN(DP_reg_sw0_n81) );
  DFFR_X1 DP_reg_sw0_Q_reg_13_ ( .D(DP_reg_sw0_n67), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_13_) );
  DFFR_X1 DP_reg_sw0_Q_reg_14_ ( .D(DP_reg_sw0_n66), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_14_) );
  DFFR_X1 DP_reg_sw0_Q_reg_15_ ( .D(DP_reg_sw0_n65), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_15_) );
  DFFR_X1 DP_reg_sw0_Q_reg_16_ ( .D(DP_reg_sw0_n48), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_16_) );
  DFFR_X1 DP_reg_sw0_Q_reg_17_ ( .D(DP_reg_sw0_n47), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_17_) );
  DFFR_X1 DP_reg_sw0_Q_reg_18_ ( .D(DP_reg_sw0_n46), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_18_) );
  DFFR_X1 DP_reg_sw0_Q_reg_19_ ( .D(DP_reg_sw0_n45), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_19_) );
  DFFR_X1 DP_reg_sw0_Q_reg_20_ ( .D(DP_reg_sw0_n44), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_20_) );
  DFFR_X1 DP_reg_sw0_Q_reg_21_ ( .D(DP_reg_sw0_n43), .CK(clk), .RN(
        DP_reg_sw0_n8), .Q(DP_sw0_21_) );
  MUX2_X1 DP_reg_sw1_U48 ( .A(DP_reg_sw1_n45), .B(DP_sw0_23_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n73) );
  INV_X1 DP_reg_sw1_U47 ( .A(DP_reg_sw1_n97), .ZN(DP_reg_sw1_n45) );
  MUX2_X1 DP_reg_sw1_U46 ( .A(DP_reg_sw1_n33), .B(DP_sw0_22_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n74) );
  INV_X1 DP_reg_sw1_U45 ( .A(DP_reg_sw1_n98), .ZN(DP_reg_sw1_n33) );
  MUX2_X1 DP_reg_sw1_U44 ( .A(DP_reg_sw1_n31), .B(DP_sw0_21_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n75) );
  INV_X1 DP_reg_sw1_U43 ( .A(DP_reg_sw1_n99), .ZN(DP_reg_sw1_n31) );
  MUX2_X1 DP_reg_sw1_U42 ( .A(DP_sw1_20_), .B(DP_sw0_20_), .S(DP_reg_sw1_n4), 
        .Z(DP_reg_sw1_n76) );
  MUX2_X1 DP_reg_sw1_U41 ( .A(DP_reg_sw1_n27), .B(DP_sw0_19_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n77) );
  INV_X1 DP_reg_sw1_U40 ( .A(DP_reg_sw1_n100), .ZN(DP_reg_sw1_n27) );
  MUX2_X1 DP_reg_sw1_U39 ( .A(DP_reg_sw1_n25), .B(DP_sw0_18_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n78) );
  INV_X1 DP_reg_sw1_U38 ( .A(DP_reg_sw1_n101), .ZN(DP_reg_sw1_n25) );
  MUX2_X1 DP_reg_sw1_U37 ( .A(DP_reg_sw1_n24), .B(DP_sw0_17_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n79) );
  INV_X1 DP_reg_sw1_U36 ( .A(DP_reg_sw1_n102), .ZN(DP_reg_sw1_n24) );
  MUX2_X1 DP_reg_sw1_U35 ( .A(DP_reg_sw1_n23), .B(DP_sw0_16_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n80) );
  INV_X1 DP_reg_sw1_U34 ( .A(DP_reg_sw1_n103), .ZN(DP_reg_sw1_n23) );
  MUX2_X1 DP_reg_sw1_U33 ( .A(DP_reg_sw1_n22), .B(DP_sw0_15_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n81) );
  INV_X1 DP_reg_sw1_U32 ( .A(DP_reg_sw1_n104), .ZN(DP_reg_sw1_n22) );
  MUX2_X1 DP_reg_sw1_U31 ( .A(DP_reg_sw1_n21), .B(DP_sw0_14_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n82) );
  INV_X1 DP_reg_sw1_U30 ( .A(DP_reg_sw1_n105), .ZN(DP_reg_sw1_n21) );
  MUX2_X1 DP_reg_sw1_U29 ( .A(DP_reg_sw1_n20), .B(DP_sw0_13_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n83) );
  INV_X1 DP_reg_sw1_U28 ( .A(DP_reg_sw1_n106), .ZN(DP_reg_sw1_n20) );
  MUX2_X1 DP_reg_sw1_U27 ( .A(DP_reg_sw1_n19), .B(DP_sw0_12_), .S(
        DP_reg_sw1_n4), .Z(DP_reg_sw1_n84) );
  INV_X1 DP_reg_sw1_U26 ( .A(DP_reg_sw1_n107), .ZN(DP_reg_sw1_n19) );
  MUX2_X1 DP_reg_sw1_U25 ( .A(DP_reg_sw1_n18), .B(DP_sw0_11_), .S(
        DP_reg_sw1_n3), .Z(DP_reg_sw1_n85) );
  INV_X1 DP_reg_sw1_U24 ( .A(DP_reg_sw1_n108), .ZN(DP_reg_sw1_n18) );
  MUX2_X1 DP_reg_sw1_U23 ( .A(DP_reg_sw1_n17), .B(DP_sw0_10_), .S(
        DP_reg_sw1_n3), .Z(DP_reg_sw1_n86) );
  INV_X1 DP_reg_sw1_U22 ( .A(DP_reg_sw1_n109), .ZN(DP_reg_sw1_n17) );
  MUX2_X1 DP_reg_sw1_U21 ( .A(DP_reg_sw1_n16), .B(DP_sw0_9_), .S(DP_reg_sw1_n3), .Z(DP_reg_sw1_n87) );
  INV_X1 DP_reg_sw1_U20 ( .A(DP_reg_sw1_n110), .ZN(DP_reg_sw1_n16) );
  MUX2_X1 DP_reg_sw1_U19 ( .A(DP_sw1_8_), .B(DP_sw0_8_), .S(DP_reg_sw1_n3), 
        .Z(DP_reg_sw1_n88) );
  MUX2_X1 DP_reg_sw1_U18 ( .A(DP_reg_sw1_n14), .B(DP_sw0_7_), .S(DP_reg_sw1_n3), .Z(DP_reg_sw1_n89) );
  INV_X1 DP_reg_sw1_U17 ( .A(DP_reg_sw1_n111), .ZN(DP_reg_sw1_n14) );
  MUX2_X1 DP_reg_sw1_U16 ( .A(DP_sw1_6_), .B(DP_sw0_6_), .S(DP_reg_sw1_n3), 
        .Z(DP_reg_sw1_n90) );
  MUX2_X1 DP_reg_sw1_U15 ( .A(DP_reg_sw1_n12), .B(DP_sw0_5_), .S(DP_reg_sw1_n3), .Z(DP_reg_sw1_n91) );
  INV_X1 DP_reg_sw1_U14 ( .A(DP_reg_sw1_n112), .ZN(DP_reg_sw1_n12) );
  MUX2_X1 DP_reg_sw1_U13 ( .A(DP_sw1_4_), .B(DP_sw0_4_), .S(DP_reg_sw1_n3), 
        .Z(DP_reg_sw1_n92) );
  MUX2_X1 DP_reg_sw1_U12 ( .A(DP_reg_sw1_n10), .B(DP_sw0_3_), .S(DP_reg_sw1_n3), .Z(DP_reg_sw1_n93) );
  INV_X1 DP_reg_sw1_U11 ( .A(DP_reg_sw1_n113), .ZN(DP_reg_sw1_n10) );
  MUX2_X1 DP_reg_sw1_U10 ( .A(DP_sw1_2_), .B(DP_sw0_2_), .S(DP_reg_sw1_n3), 
        .Z(DP_reg_sw1_n94) );
  MUX2_X1 DP_reg_sw1_U9 ( .A(DP_reg_sw1_n8), .B(DP_sw0_1_), .S(DP_reg_sw1_n3), 
        .Z(DP_reg_sw1_n95) );
  INV_X1 DP_reg_sw1_U8 ( .A(DP_reg_sw1_n114), .ZN(DP_reg_sw1_n8) );
  MUX2_X1 DP_reg_sw1_U7 ( .A(DP_reg_sw1_n7), .B(DP_sw0_0_), .S(DP_reg_sw1_n3), 
        .Z(DP_reg_sw1_n96) );
  BUF_X1 DP_reg_sw1_U6 ( .A(DP_n10), .Z(DP_reg_sw1_n5) );
  BUF_X1 DP_reg_sw1_U5 ( .A(DP_n10), .Z(DP_reg_sw1_n6) );
  BUF_X1 DP_reg_sw1_U4 ( .A(sw_regs_en_int), .Z(DP_reg_sw1_n4) );
  BUF_X1 DP_reg_sw1_U3 ( .A(sw_regs_en_int), .Z(DP_reg_sw1_n3) );
  INV_X4 DP_reg_sw1_U2 ( .A(DP_reg_sw1_n1), .ZN(DP_sw1_0_) );
  DFFR_X1 DP_reg_sw1_Q_reg_0_ ( .D(DP_reg_sw1_n96), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_reg_sw1_n7), .QN(DP_reg_sw1_n1) );
  DFFR_X1 DP_reg_sw1_Q_reg_1_ ( .D(DP_reg_sw1_n95), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_1_), .QN(DP_reg_sw1_n114) );
  DFFR_X1 DP_reg_sw1_Q_reg_2_ ( .D(DP_reg_sw1_n94), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_2_) );
  DFFR_X1 DP_reg_sw1_Q_reg_3_ ( .D(DP_reg_sw1_n93), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_3_), .QN(DP_reg_sw1_n113) );
  DFFR_X1 DP_reg_sw1_Q_reg_4_ ( .D(DP_reg_sw1_n92), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_4_) );
  DFFR_X1 DP_reg_sw1_Q_reg_5_ ( .D(DP_reg_sw1_n91), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_5_), .QN(DP_reg_sw1_n112) );
  DFFR_X1 DP_reg_sw1_Q_reg_6_ ( .D(DP_reg_sw1_n90), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_6_) );
  DFFR_X1 DP_reg_sw1_Q_reg_7_ ( .D(DP_reg_sw1_n89), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_7_), .QN(DP_reg_sw1_n111) );
  DFFR_X1 DP_reg_sw1_Q_reg_8_ ( .D(DP_reg_sw1_n88), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_8_) );
  DFFR_X1 DP_reg_sw1_Q_reg_9_ ( .D(DP_reg_sw1_n87), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_9_), .QN(DP_reg_sw1_n110) );
  DFFR_X1 DP_reg_sw1_Q_reg_10_ ( .D(DP_reg_sw1_n86), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_10_), .QN(DP_reg_sw1_n109) );
  DFFR_X1 DP_reg_sw1_Q_reg_11_ ( .D(DP_reg_sw1_n85), .CK(clk), .RN(
        DP_reg_sw1_n6), .Q(DP_sw1_11_), .QN(DP_reg_sw1_n108) );
  DFFR_X1 DP_reg_sw1_Q_reg_12_ ( .D(DP_reg_sw1_n84), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_12_), .QN(DP_reg_sw1_n107) );
  DFFR_X1 DP_reg_sw1_Q_reg_13_ ( .D(DP_reg_sw1_n83), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_13_), .QN(DP_reg_sw1_n106) );
  DFFR_X1 DP_reg_sw1_Q_reg_14_ ( .D(DP_reg_sw1_n82), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_14_), .QN(DP_reg_sw1_n105) );
  DFFR_X1 DP_reg_sw1_Q_reg_15_ ( .D(DP_reg_sw1_n81), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_15_), .QN(DP_reg_sw1_n104) );
  DFFR_X1 DP_reg_sw1_Q_reg_16_ ( .D(DP_reg_sw1_n80), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_16_), .QN(DP_reg_sw1_n103) );
  DFFR_X1 DP_reg_sw1_Q_reg_17_ ( .D(DP_reg_sw1_n79), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_17_), .QN(DP_reg_sw1_n102) );
  DFFR_X1 DP_reg_sw1_Q_reg_18_ ( .D(DP_reg_sw1_n78), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_18_), .QN(DP_reg_sw1_n101) );
  DFFR_X1 DP_reg_sw1_Q_reg_19_ ( .D(DP_reg_sw1_n77), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_19_), .QN(DP_reg_sw1_n100) );
  DFFR_X1 DP_reg_sw1_Q_reg_20_ ( .D(DP_reg_sw1_n76), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_20_) );
  DFFR_X1 DP_reg_sw1_Q_reg_21_ ( .D(DP_reg_sw1_n75), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_21_), .QN(DP_reg_sw1_n99) );
  DFFR_X1 DP_reg_sw1_Q_reg_22_ ( .D(DP_reg_sw1_n74), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_22_), .QN(DP_reg_sw1_n98) );
  DFFR_X1 DP_reg_sw1_Q_reg_23_ ( .D(DP_reg_sw1_n73), .CK(clk), .RN(
        DP_reg_sw1_n5), .Q(DP_sw1_23_), .QN(DP_reg_sw1_n97) );
  MUX2_X1 DP_reg_sw2_U27 ( .A(DP_sw2[23]), .B(DP_sw1_23_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n27) );
  MUX2_X1 DP_reg_sw2_U26 ( .A(DP_sw2[22]), .B(DP_sw1_22_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n28) );
  MUX2_X1 DP_reg_sw2_U25 ( .A(DP_sw2[21]), .B(DP_sw1_21_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n29) );
  MUX2_X1 DP_reg_sw2_U24 ( .A(DP_sw2[20]), .B(DP_sw1_20_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n30) );
  MUX2_X1 DP_reg_sw2_U23 ( .A(DP_sw2[19]), .B(DP_sw1_19_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n31) );
  MUX2_X1 DP_reg_sw2_U22 ( .A(DP_sw2[18]), .B(DP_sw1_18_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n32) );
  MUX2_X1 DP_reg_sw2_U21 ( .A(DP_sw2[17]), .B(DP_sw1_17_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n33) );
  MUX2_X1 DP_reg_sw2_U20 ( .A(DP_sw2[16]), .B(DP_sw1_16_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n34) );
  MUX2_X1 DP_reg_sw2_U19 ( .A(DP_sw2[15]), .B(DP_sw1_15_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n35) );
  MUX2_X1 DP_reg_sw2_U18 ( .A(DP_sw2[14]), .B(DP_sw1_14_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n36) );
  MUX2_X1 DP_reg_sw2_U17 ( .A(DP_sw2[13]), .B(DP_sw1_13_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n37) );
  MUX2_X1 DP_reg_sw2_U16 ( .A(DP_sw2[12]), .B(DP_sw1_12_), .S(DP_reg_sw2_n26), 
        .Z(DP_reg_sw2_n38) );
  MUX2_X1 DP_reg_sw2_U15 ( .A(DP_sw2[11]), .B(DP_sw1_11_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n39) );
  MUX2_X1 DP_reg_sw2_U14 ( .A(DP_sw2[10]), .B(DP_sw1_10_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n40) );
  MUX2_X1 DP_reg_sw2_U13 ( .A(DP_sw2[9]), .B(DP_sw1_9_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n41) );
  MUX2_X1 DP_reg_sw2_U12 ( .A(DP_sw2[8]), .B(DP_sw1_8_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n42) );
  MUX2_X1 DP_reg_sw2_U11 ( .A(DP_sw2[7]), .B(DP_sw1_7_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n43) );
  MUX2_X1 DP_reg_sw2_U10 ( .A(DP_sw2[6]), .B(DP_sw1_6_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n44) );
  MUX2_X1 DP_reg_sw2_U9 ( .A(DP_sw2[5]), .B(DP_sw1_5_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n45) );
  MUX2_X1 DP_reg_sw2_U8 ( .A(DP_sw2[4]), .B(DP_sw1_4_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n46) );
  MUX2_X1 DP_reg_sw2_U7 ( .A(DP_sw2[3]), .B(DP_sw1_3_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n47) );
  MUX2_X1 DP_reg_sw2_U6 ( .A(DP_sw2[2]), .B(DP_sw1_2_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n48) );
  MUX2_X1 DP_reg_sw2_U5 ( .A(DP_sw2[1]), .B(DP_sw1_1_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n51) );
  MUX2_X1 DP_reg_sw2_U4 ( .A(DP_sw2[0]), .B(DP_sw1_0_), .S(DP_reg_sw2_n25), 
        .Z(DP_reg_sw2_n52) );
  BUF_X1 DP_reg_sw2_U3 ( .A(sw_regs_en_int), .Z(DP_reg_sw2_n26) );
  BUF_X1 DP_reg_sw2_U2 ( .A(sw_regs_en_int), .Z(DP_reg_sw2_n25) );
  DFFR_X1 DP_reg_sw2_Q_reg_2_ ( .D(DP_reg_sw2_n48), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[2]) );
  DFFR_X1 DP_reg_sw2_Q_reg_4_ ( .D(DP_reg_sw2_n46), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[4]) );
  DFFR_X1 DP_reg_sw2_Q_reg_6_ ( .D(DP_reg_sw2_n44), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[6]) );
  DFFR_X1 DP_reg_sw2_Q_reg_8_ ( .D(DP_reg_sw2_n42), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[8]) );
  DFFR_X1 DP_reg_sw2_Q_reg_20_ ( .D(DP_reg_sw2_n30), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[20]) );
  DFFR_X1 DP_reg_sw2_Q_reg_10_ ( .D(DP_reg_sw2_n40), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[10]) );
  DFFR_X1 DP_reg_sw2_Q_reg_12_ ( .D(DP_reg_sw2_n38), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[12]) );
  DFFR_X1 DP_reg_sw2_Q_reg_14_ ( .D(DP_reg_sw2_n36), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[14]) );
  DFFR_X1 DP_reg_sw2_Q_reg_16_ ( .D(DP_reg_sw2_n34), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[16]) );
  DFFR_X1 DP_reg_sw2_Q_reg_18_ ( .D(DP_reg_sw2_n32), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[18]) );
  DFFR_X1 DP_reg_sw2_Q_reg_22_ ( .D(DP_reg_sw2_n28), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[22]) );
  DFFR_X1 DP_reg_sw2_Q_reg_1_ ( .D(DP_reg_sw2_n51), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[1]) );
  DFFR_X1 DP_reg_sw2_Q_reg_3_ ( .D(DP_reg_sw2_n47), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[3]) );
  DFFR_X1 DP_reg_sw2_Q_reg_5_ ( .D(DP_reg_sw2_n45), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[5]) );
  DFFR_X1 DP_reg_sw2_Q_reg_7_ ( .D(DP_reg_sw2_n43), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[7]) );
  DFFR_X1 DP_reg_sw2_Q_reg_9_ ( .D(DP_reg_sw2_n41), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[9]) );
  DFFR_X1 DP_reg_sw2_Q_reg_11_ ( .D(DP_reg_sw2_n39), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[11]) );
  DFFR_X1 DP_reg_sw2_Q_reg_13_ ( .D(DP_reg_sw2_n37), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[13]) );
  DFFR_X1 DP_reg_sw2_Q_reg_15_ ( .D(DP_reg_sw2_n35), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[15]) );
  DFFR_X1 DP_reg_sw2_Q_reg_17_ ( .D(DP_reg_sw2_n33), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[17]) );
  DFFR_X1 DP_reg_sw2_Q_reg_19_ ( .D(DP_reg_sw2_n31), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[19]) );
  DFFR_X1 DP_reg_sw2_Q_reg_21_ ( .D(DP_reg_sw2_n29), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[21]) );
  DFFR_X1 DP_reg_sw2_Q_reg_23_ ( .D(DP_reg_sw2_n27), .CK(clk), .RN(DP_n10), 
        .Q(DP_sw2[23]) );
  DFFR_X1 DP_reg_sw2_Q_reg_0_ ( .D(DP_reg_sw2_n52), .CK(clk), .RN(DP_n10), .Q(
        DP_sw2[0]) );
  NAND2_X1 DP_reg_ret0_U52 ( .A1(DP_reg_ret0_n76), .A2(DP_reg_ret0_n75), .ZN(
        DP_reg_ret0_n77) );
  NAND2_X1 DP_reg_ret0_U51 ( .A1(DP_ret0[23]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n75) );
  NAND2_X1 DP_reg_ret0_U50 ( .A1(DP_sw0_coeff_ret0[23]), .A2(1'b1), .ZN(
        DP_reg_ret0_n76) );
  NAND2_X1 DP_reg_ret0_U49 ( .A1(DP_reg_ret0_n47), .A2(DP_reg_ret0_n48), .ZN(
        DP_reg_ret0_n78) );
  NAND2_X1 DP_reg_ret0_U48 ( .A1(DP_sw0_coeff_ret0[22]), .A2(1'b1), .ZN(
        DP_reg_ret0_n47) );
  NAND2_X1 DP_reg_ret0_U47 ( .A1(DP_ret0[22]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n48) );
  NAND2_X1 DP_reg_ret0_U46 ( .A1(DP_reg_ret0_n44), .A2(DP_reg_ret0_n45), .ZN(
        DP_reg_ret0_n79) );
  NAND2_X1 DP_reg_ret0_U45 ( .A1(DP_sw0_coeff_ret0[21]), .A2(1'b1), .ZN(
        DP_reg_ret0_n44) );
  NAND2_X1 DP_reg_ret0_U44 ( .A1(DP_ret0[21]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n45) );
  NAND2_X1 DP_reg_ret0_U43 ( .A1(DP_reg_ret0_n41), .A2(DP_reg_ret0_n42), .ZN(
        DP_reg_ret0_n80) );
  NAND2_X1 DP_reg_ret0_U42 ( .A1(DP_sw0_coeff_ret0[20]), .A2(1'b1), .ZN(
        DP_reg_ret0_n41) );
  NAND2_X1 DP_reg_ret0_U41 ( .A1(DP_ret0[20]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n42) );
  NAND2_X1 DP_reg_ret0_U40 ( .A1(DP_reg_ret0_n38), .A2(DP_reg_ret0_n39), .ZN(
        DP_reg_ret0_n81) );
  NAND2_X1 DP_reg_ret0_U39 ( .A1(DP_sw0_coeff_ret0[19]), .A2(1'b1), .ZN(
        DP_reg_ret0_n38) );
  NAND2_X1 DP_reg_ret0_U38 ( .A1(DP_ret0[19]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n39) );
  NAND2_X1 DP_reg_ret0_U37 ( .A1(DP_reg_ret0_n35), .A2(DP_reg_ret0_n36), .ZN(
        DP_reg_ret0_n82) );
  NAND2_X1 DP_reg_ret0_U36 ( .A1(DP_sw0_coeff_ret0[18]), .A2(1'b1), .ZN(
        DP_reg_ret0_n35) );
  NAND2_X1 DP_reg_ret0_U35 ( .A1(DP_ret0[18]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n36) );
  NAND2_X1 DP_reg_ret0_U34 ( .A1(DP_reg_ret0_n32), .A2(DP_reg_ret0_n33), .ZN(
        DP_reg_ret0_n83) );
  NAND2_X1 DP_reg_ret0_U33 ( .A1(DP_sw0_coeff_ret0[17]), .A2(1'b1), .ZN(
        DP_reg_ret0_n32) );
  NAND2_X1 DP_reg_ret0_U32 ( .A1(DP_ret0[17]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n33) );
  NAND2_X1 DP_reg_ret0_U31 ( .A1(DP_reg_ret0_n29), .A2(DP_reg_ret0_n30), .ZN(
        DP_reg_ret0_n84) );
  NAND2_X1 DP_reg_ret0_U30 ( .A1(DP_sw0_coeff_ret0[16]), .A2(1'b1), .ZN(
        DP_reg_ret0_n29) );
  NAND2_X1 DP_reg_ret0_U29 ( .A1(DP_ret0[16]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n30) );
  NAND2_X1 DP_reg_ret0_U28 ( .A1(DP_reg_ret0_n26), .A2(DP_reg_ret0_n27), .ZN(
        DP_reg_ret0_n85) );
  NAND2_X1 DP_reg_ret0_U27 ( .A1(DP_sw0_coeff_ret0[15]), .A2(1'b1), .ZN(
        DP_reg_ret0_n26) );
  NAND2_X1 DP_reg_ret0_U26 ( .A1(DP_ret0[15]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n27) );
  NAND2_X1 DP_reg_ret0_U25 ( .A1(DP_reg_ret0_n23), .A2(DP_reg_ret0_n24), .ZN(
        DP_reg_ret0_n86) );
  NAND2_X1 DP_reg_ret0_U24 ( .A1(DP_sw0_coeff_ret0[14]), .A2(1'b1), .ZN(
        DP_reg_ret0_n23) );
  NAND2_X1 DP_reg_ret0_U23 ( .A1(DP_ret0[14]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n24) );
  NAND2_X1 DP_reg_ret0_U22 ( .A1(DP_reg_ret0_n20), .A2(DP_reg_ret0_n21), .ZN(
        DP_reg_ret0_n87) );
  NAND2_X1 DP_reg_ret0_U21 ( .A1(DP_sw0_coeff_ret0[13]), .A2(1'b1), .ZN(
        DP_reg_ret0_n20) );
  NAND2_X1 DP_reg_ret0_U20 ( .A1(DP_ret0[13]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n21) );
  NAND2_X1 DP_reg_ret0_U19 ( .A1(DP_reg_ret0_n18), .A2(DP_reg_ret0_n17), .ZN(
        DP_reg_ret0_n88) );
  NAND2_X1 DP_reg_ret0_U18 ( .A1(DP_ret0[12]), .A2(DP_reg_ret0_n73), .ZN(
        DP_reg_ret0_n17) );
  INV_X1 DP_reg_ret0_U17 ( .A(1'b1), .ZN(DP_reg_ret0_n73) );
  NAND2_X1 DP_reg_ret0_U16 ( .A1(DP_sw0_coeff_ret0[12]), .A2(1'b1), .ZN(
        DP_reg_ret0_n18) );
  MUX2_X1 DP_reg_ret0_U15 ( .A(DP_ret0[11]), .B(DP_sw0_coeff_ret0[11]), .S(
        1'b1), .Z(DP_reg_ret0_n89) );
  MUX2_X1 DP_reg_ret0_U14 ( .A(DP_ret0[10]), .B(DP_sw0_coeff_ret0[10]), .S(
        1'b1), .Z(DP_reg_ret0_n90) );
  MUX2_X1 DP_reg_ret0_U13 ( .A(DP_ret0[9]), .B(DP_sw0_coeff_ret0[9]), .S(1'b1), 
        .Z(DP_reg_ret0_n91) );
  MUX2_X1 DP_reg_ret0_U12 ( .A(DP_ret0[8]), .B(DP_sw0_coeff_ret0[8]), .S(1'b1), 
        .Z(DP_reg_ret0_n92) );
  MUX2_X1 DP_reg_ret0_U11 ( .A(DP_ret0[7]), .B(DP_sw0_coeff_ret0[7]), .S(1'b1), 
        .Z(DP_reg_ret0_n93) );
  MUX2_X1 DP_reg_ret0_U10 ( .A(DP_ret0[6]), .B(DP_sw0_coeff_ret0[6]), .S(1'b1), 
        .Z(DP_reg_ret0_n94) );
  MUX2_X1 DP_reg_ret0_U9 ( .A(DP_ret0[5]), .B(DP_sw0_coeff_ret0[5]), .S(1'b1), 
        .Z(DP_reg_ret0_n95) );
  MUX2_X1 DP_reg_ret0_U8 ( .A(DP_ret0[4]), .B(DP_sw0_coeff_ret0[4]), .S(1'b1), 
        .Z(DP_reg_ret0_n96) );
  MUX2_X1 DP_reg_ret0_U7 ( .A(DP_ret0[3]), .B(DP_sw0_coeff_ret0[3]), .S(1'b1), 
        .Z(DP_reg_ret0_n97) );
  MUX2_X1 DP_reg_ret0_U6 ( .A(DP_ret0[2]), .B(DP_sw0_coeff_ret0[2]), .S(1'b1), 
        .Z(DP_reg_ret0_n98) );
  MUX2_X1 DP_reg_ret0_U5 ( .A(DP_ret0[1]), .B(DP_sw0_coeff_ret0[1]), .S(1'b1), 
        .Z(DP_reg_ret0_n99) );
  MUX2_X1 DP_reg_ret0_U4 ( .A(DP_ret0[0]), .B(DP_sw0_coeff_ret0[0]), .S(1'b1), 
        .Z(DP_reg_ret0_n100) );
  BUF_X1 DP_reg_ret0_U3 ( .A(DP_n9), .Z(DP_reg_ret0_n5) );
  BUF_X1 DP_reg_ret0_U2 ( .A(DP_n9), .Z(DP_reg_ret0_n6) );
  DFFR_X1 DP_reg_ret0_Q_reg_3_ ( .D(DP_reg_ret0_n97), .CK(clk), .RN(DP_n9), 
        .Q(DP_ret0[3]) );
  DFFR_X1 DP_reg_ret0_Q_reg_0_ ( .D(DP_reg_ret0_n100), .CK(clk), .RN(DP_n9), 
        .Q(DP_ret0[0]) );
  DFFR_X1 DP_reg_ret0_Q_reg_1_ ( .D(DP_reg_ret0_n99), .CK(clk), .RN(DP_n9), 
        .Q(DP_ret0[1]) );
  DFFR_X1 DP_reg_ret0_Q_reg_21_ ( .D(DP_reg_ret0_n79), .CK(clk), .RN(DP_n9), 
        .Q(DP_ret0[21]) );
  DFFR_X1 DP_reg_ret0_Q_reg_2_ ( .D(DP_reg_ret0_n98), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[2]) );
  DFFR_X1 DP_reg_ret0_Q_reg_4_ ( .D(DP_reg_ret0_n96), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[4]) );
  DFFR_X1 DP_reg_ret0_Q_reg_5_ ( .D(DP_reg_ret0_n95), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[5]) );
  DFFR_X1 DP_reg_ret0_Q_reg_6_ ( .D(DP_reg_ret0_n94), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[6]) );
  DFFR_X1 DP_reg_ret0_Q_reg_7_ ( .D(DP_reg_ret0_n93), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[7]) );
  DFFR_X1 DP_reg_ret0_Q_reg_8_ ( .D(DP_reg_ret0_n92), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[8]) );
  DFFR_X1 DP_reg_ret0_Q_reg_9_ ( .D(DP_reg_ret0_n91), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[9]) );
  DFFR_X1 DP_reg_ret0_Q_reg_10_ ( .D(DP_reg_ret0_n90), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[10]) );
  DFFR_X1 DP_reg_ret0_Q_reg_11_ ( .D(DP_reg_ret0_n89), .CK(clk), .RN(
        DP_reg_ret0_n6), .Q(DP_ret0[11]) );
  DFFR_X1 DP_reg_ret0_Q_reg_12_ ( .D(DP_reg_ret0_n88), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[12]) );
  DFFR_X1 DP_reg_ret0_Q_reg_13_ ( .D(DP_reg_ret0_n87), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[13]) );
  DFFR_X1 DP_reg_ret0_Q_reg_14_ ( .D(DP_reg_ret0_n86), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[14]) );
  DFFR_X1 DP_reg_ret0_Q_reg_15_ ( .D(DP_reg_ret0_n85), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[15]) );
  DFFR_X1 DP_reg_ret0_Q_reg_16_ ( .D(DP_reg_ret0_n84), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[16]) );
  DFFR_X1 DP_reg_ret0_Q_reg_17_ ( .D(DP_reg_ret0_n83), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[17]) );
  DFFR_X1 DP_reg_ret0_Q_reg_18_ ( .D(DP_reg_ret0_n82), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[18]) );
  DFFR_X1 DP_reg_ret0_Q_reg_19_ ( .D(DP_reg_ret0_n81), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[19]) );
  DFFR_X1 DP_reg_ret0_Q_reg_20_ ( .D(DP_reg_ret0_n80), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[20]) );
  DFFR_X1 DP_reg_ret0_Q_reg_22_ ( .D(DP_reg_ret0_n78), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[22]) );
  DFFR_X1 DP_reg_ret0_Q_reg_23_ ( .D(DP_reg_ret0_n77), .CK(clk), .RN(
        DP_reg_ret0_n5), .Q(DP_ret0[23]) );
  NAND2_X1 DP_reg_ret1_U52 ( .A1(DP_reg_ret1_n79), .A2(DP_reg_ret1_n78), .ZN(
        DP_reg_ret1_n80) );
  NAND2_X1 DP_reg_ret1_U51 ( .A1(DP_ret1[23]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n78) );
  NAND2_X1 DP_reg_ret1_U50 ( .A1(DP_sw1_coeff_ret1[23]), .A2(1'b1), .ZN(
        DP_reg_ret1_n79) );
  NAND2_X1 DP_reg_ret1_U49 ( .A1(DP_reg_ret1_n74), .A2(DP_reg_ret1_n75), .ZN(
        DP_reg_ret1_n81) );
  NAND2_X1 DP_reg_ret1_U48 ( .A1(DP_sw1_coeff_ret1[22]), .A2(1'b1), .ZN(
        DP_reg_ret1_n74) );
  NAND2_X1 DP_reg_ret1_U47 ( .A1(DP_ret1[22]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n75) );
  NAND2_X1 DP_reg_ret1_U46 ( .A1(DP_reg_ret1_n47), .A2(DP_reg_ret1_n48), .ZN(
        DP_reg_ret1_n82) );
  NAND2_X1 DP_reg_ret1_U45 ( .A1(DP_sw1_coeff_ret1[21]), .A2(1'b1), .ZN(
        DP_reg_ret1_n47) );
  NAND2_X1 DP_reg_ret1_U44 ( .A1(DP_ret1[21]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n48) );
  NAND2_X1 DP_reg_ret1_U43 ( .A1(DP_reg_ret1_n44), .A2(DP_reg_ret1_n45), .ZN(
        DP_reg_ret1_n83) );
  NAND2_X1 DP_reg_ret1_U42 ( .A1(DP_sw1_coeff_ret1[20]), .A2(1'b1), .ZN(
        DP_reg_ret1_n44) );
  NAND2_X1 DP_reg_ret1_U41 ( .A1(DP_ret1[20]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n45) );
  NAND2_X1 DP_reg_ret1_U40 ( .A1(DP_reg_ret1_n41), .A2(DP_reg_ret1_n42), .ZN(
        DP_reg_ret1_n84) );
  NAND2_X1 DP_reg_ret1_U39 ( .A1(DP_sw1_coeff_ret1[19]), .A2(1'b1), .ZN(
        DP_reg_ret1_n41) );
  NAND2_X1 DP_reg_ret1_U38 ( .A1(DP_ret1[19]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n42) );
  NAND2_X1 DP_reg_ret1_U37 ( .A1(DP_reg_ret1_n38), .A2(DP_reg_ret1_n39), .ZN(
        DP_reg_ret1_n85) );
  NAND2_X1 DP_reg_ret1_U36 ( .A1(DP_sw1_coeff_ret1[18]), .A2(1'b1), .ZN(
        DP_reg_ret1_n38) );
  NAND2_X1 DP_reg_ret1_U35 ( .A1(DP_ret1[18]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n39) );
  NAND2_X1 DP_reg_ret1_U34 ( .A1(DP_reg_ret1_n35), .A2(DP_reg_ret1_n36), .ZN(
        DP_reg_ret1_n86) );
  NAND2_X1 DP_reg_ret1_U33 ( .A1(DP_sw1_coeff_ret1[17]), .A2(1'b1), .ZN(
        DP_reg_ret1_n35) );
  NAND2_X1 DP_reg_ret1_U32 ( .A1(DP_ret1[17]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n36) );
  NAND2_X1 DP_reg_ret1_U31 ( .A1(DP_reg_ret1_n32), .A2(DP_reg_ret1_n33), .ZN(
        DP_reg_ret1_n87) );
  NAND2_X1 DP_reg_ret1_U30 ( .A1(DP_sw1_coeff_ret1[16]), .A2(1'b1), .ZN(
        DP_reg_ret1_n32) );
  NAND2_X1 DP_reg_ret1_U29 ( .A1(DP_ret1[16]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n33) );
  NAND2_X1 DP_reg_ret1_U28 ( .A1(DP_reg_ret1_n29), .A2(DP_reg_ret1_n30), .ZN(
        DP_reg_ret1_n88) );
  NAND2_X1 DP_reg_ret1_U27 ( .A1(DP_sw1_coeff_ret1[15]), .A2(1'b1), .ZN(
        DP_reg_ret1_n29) );
  NAND2_X1 DP_reg_ret1_U26 ( .A1(DP_ret1[15]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n30) );
  NAND2_X1 DP_reg_ret1_U25 ( .A1(DP_reg_ret1_n26), .A2(DP_reg_ret1_n27), .ZN(
        DP_reg_ret1_n89) );
  NAND2_X1 DP_reg_ret1_U24 ( .A1(DP_sw1_coeff_ret1[14]), .A2(1'b1), .ZN(
        DP_reg_ret1_n26) );
  NAND2_X1 DP_reg_ret1_U23 ( .A1(DP_ret1[14]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n27) );
  NAND2_X1 DP_reg_ret1_U22 ( .A1(DP_reg_ret1_n23), .A2(DP_reg_ret1_n24), .ZN(
        DP_reg_ret1_n90) );
  NAND2_X1 DP_reg_ret1_U21 ( .A1(DP_sw1_coeff_ret1[13]), .A2(1'b1), .ZN(
        DP_reg_ret1_n23) );
  NAND2_X1 DP_reg_ret1_U20 ( .A1(DP_ret1[13]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n24) );
  NAND2_X1 DP_reg_ret1_U19 ( .A1(DP_reg_ret1_n21), .A2(DP_reg_ret1_n20), .ZN(
        DP_reg_ret1_n91) );
  NAND2_X1 DP_reg_ret1_U18 ( .A1(DP_ret1[12]), .A2(DP_reg_ret1_n76), .ZN(
        DP_reg_ret1_n20) );
  INV_X1 DP_reg_ret1_U17 ( .A(1'b1), .ZN(DP_reg_ret1_n76) );
  NAND2_X1 DP_reg_ret1_U16 ( .A1(DP_sw1_coeff_ret1[12]), .A2(1'b1), .ZN(
        DP_reg_ret1_n21) );
  MUX2_X1 DP_reg_ret1_U15 ( .A(DP_ret1[11]), .B(DP_sw1_coeff_ret1[11]), .S(
        1'b1), .Z(DP_reg_ret1_n92) );
  MUX2_X1 DP_reg_ret1_U14 ( .A(DP_ret1[10]), .B(DP_sw1_coeff_ret1[10]), .S(
        1'b1), .Z(DP_reg_ret1_n93) );
  MUX2_X1 DP_reg_ret1_U13 ( .A(DP_ret1[9]), .B(DP_sw1_coeff_ret1[9]), .S(1'b1), 
        .Z(DP_reg_ret1_n94) );
  MUX2_X1 DP_reg_ret1_U12 ( .A(DP_ret1[8]), .B(DP_sw1_coeff_ret1[8]), .S(1'b1), 
        .Z(DP_reg_ret1_n95) );
  MUX2_X1 DP_reg_ret1_U11 ( .A(DP_ret1[7]), .B(DP_sw1_coeff_ret1[7]), .S(1'b1), 
        .Z(DP_reg_ret1_n96) );
  MUX2_X1 DP_reg_ret1_U10 ( .A(DP_ret1[6]), .B(DP_sw1_coeff_ret1[6]), .S(1'b1), 
        .Z(DP_reg_ret1_n97) );
  MUX2_X1 DP_reg_ret1_U9 ( .A(DP_ret1[5]), .B(DP_sw1_coeff_ret1[5]), .S(1'b1), 
        .Z(DP_reg_ret1_n98) );
  MUX2_X1 DP_reg_ret1_U8 ( .A(DP_ret1[4]), .B(DP_sw1_coeff_ret1[4]), .S(1'b1), 
        .Z(DP_reg_ret1_n99) );
  MUX2_X1 DP_reg_ret1_U7 ( .A(DP_ret1[3]), .B(DP_sw1_coeff_ret1[3]), .S(1'b1), 
        .Z(DP_reg_ret1_n100) );
  MUX2_X1 DP_reg_ret1_U6 ( .A(DP_ret1[2]), .B(DP_sw1_coeff_ret1[2]), .S(1'b1), 
        .Z(DP_reg_ret1_n101) );
  MUX2_X1 DP_reg_ret1_U5 ( .A(DP_ret1[1]), .B(DP_sw1_coeff_ret1[1]), .S(1'b1), 
        .Z(DP_reg_ret1_n102) );
  MUX2_X1 DP_reg_ret1_U4 ( .A(DP_ret1[0]), .B(DP_sw1_coeff_ret1[0]), .S(1'b1), 
        .Z(DP_reg_ret1_n103) );
  BUF_X1 DP_reg_ret1_U3 ( .A(DP_n9), .Z(DP_reg_ret1_n5) );
  BUF_X1 DP_reg_ret1_U2 ( .A(DP_n9), .Z(DP_reg_ret1_n6) );
  DFFR_X1 DP_reg_ret1_Q_reg_16_ ( .D(DP_reg_ret1_n87), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[16]) );
  DFFR_X1 DP_reg_ret1_Q_reg_19_ ( .D(DP_reg_ret1_n84), .CK(clk), .RN(DP_n9), 
        .Q(DP_ret1[19]) );
  DFFR_X1 DP_reg_ret1_Q_reg_17_ ( .D(DP_reg_ret1_n86), .CK(clk), .RN(DP_n9), 
        .Q(DP_ret1[17]) );
  DFFR_X1 DP_reg_ret1_Q_reg_22_ ( .D(DP_reg_ret1_n81), .CK(clk), .RN(DP_n9), 
        .Q(DP_ret1[22]) );
  DFFR_X1 DP_reg_ret1_Q_reg_0_ ( .D(DP_reg_ret1_n103), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[0]) );
  DFFR_X1 DP_reg_ret1_Q_reg_1_ ( .D(DP_reg_ret1_n102), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[1]) );
  DFFR_X1 DP_reg_ret1_Q_reg_2_ ( .D(DP_reg_ret1_n101), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[2]) );
  DFFR_X1 DP_reg_ret1_Q_reg_3_ ( .D(DP_reg_ret1_n100), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[3]) );
  DFFR_X1 DP_reg_ret1_Q_reg_4_ ( .D(DP_reg_ret1_n99), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[4]) );
  DFFR_X1 DP_reg_ret1_Q_reg_5_ ( .D(DP_reg_ret1_n98), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[5]) );
  DFFR_X1 DP_reg_ret1_Q_reg_6_ ( .D(DP_reg_ret1_n97), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[6]) );
  DFFR_X1 DP_reg_ret1_Q_reg_7_ ( .D(DP_reg_ret1_n96), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[7]) );
  DFFR_X1 DP_reg_ret1_Q_reg_8_ ( .D(DP_reg_ret1_n95), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[8]) );
  DFFR_X1 DP_reg_ret1_Q_reg_9_ ( .D(DP_reg_ret1_n94), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[9]) );
  DFFR_X1 DP_reg_ret1_Q_reg_10_ ( .D(DP_reg_ret1_n93), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[10]) );
  DFFR_X1 DP_reg_ret1_Q_reg_11_ ( .D(DP_reg_ret1_n92), .CK(clk), .RN(
        DP_reg_ret1_n6), .Q(DP_ret1[11]) );
  DFFR_X1 DP_reg_ret1_Q_reg_12_ ( .D(DP_reg_ret1_n91), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[12]) );
  DFFR_X1 DP_reg_ret1_Q_reg_13_ ( .D(DP_reg_ret1_n90), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[13]) );
  DFFR_X1 DP_reg_ret1_Q_reg_14_ ( .D(DP_reg_ret1_n89), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[14]) );
  DFFR_X1 DP_reg_ret1_Q_reg_15_ ( .D(DP_reg_ret1_n88), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[15]) );
  DFFR_X1 DP_reg_ret1_Q_reg_18_ ( .D(DP_reg_ret1_n85), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[18]) );
  DFFR_X1 DP_reg_ret1_Q_reg_20_ ( .D(DP_reg_ret1_n83), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[20]) );
  DFFR_X1 DP_reg_ret1_Q_reg_21_ ( .D(DP_reg_ret1_n82), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[21]) );
  DFFR_X1 DP_reg_ret1_Q_reg_23_ ( .D(DP_reg_ret1_n80), .CK(clk), .RN(
        DP_reg_ret1_n5), .Q(DP_ret1[23]) );
  MUX2_X1 DP_reg_pipe00_U35 ( .A(DP_pipe00[23]), .B(DP_w_23_), .S(1'b1), .Z(
        DP_reg_pipe00_n36) );
  MUX2_X1 DP_reg_pipe00_U34 ( .A(DP_pipe00[22]), .B(DP_w_22_), .S(1'b1), .Z(
        DP_reg_pipe00_n37) );
  MUX2_X1 DP_reg_pipe00_U33 ( .A(DP_pipe00[21]), .B(DP_w_21_), .S(1'b1), .Z(
        DP_reg_pipe00_n38) );
  MUX2_X1 DP_reg_pipe00_U32 ( .A(DP_pipe00[20]), .B(DP_w_20_), .S(1'b1), .Z(
        DP_reg_pipe00_n39) );
  MUX2_X1 DP_reg_pipe00_U31 ( .A(DP_pipe00[19]), .B(DP_w_19_), .S(1'b1), .Z(
        DP_reg_pipe00_n40) );
  MUX2_X1 DP_reg_pipe00_U30 ( .A(DP_pipe00[18]), .B(DP_w_18_), .S(1'b1), .Z(
        DP_reg_pipe00_n41) );
  MUX2_X1 DP_reg_pipe00_U29 ( .A(DP_pipe00[17]), .B(DP_w_17_), .S(1'b1), .Z(
        DP_reg_pipe00_n42) );
  MUX2_X1 DP_reg_pipe00_U28 ( .A(DP_pipe00[16]), .B(DP_w_16_), .S(1'b1), .Z(
        DP_reg_pipe00_n43) );
  MUX2_X1 DP_reg_pipe00_U27 ( .A(DP_pipe00[15]), .B(DP_w_15_), .S(1'b1), .Z(
        DP_reg_pipe00_n44) );
  MUX2_X1 DP_reg_pipe00_U26 ( .A(DP_pipe00[14]), .B(DP_w_14_), .S(1'b1), .Z(
        DP_reg_pipe00_n45) );
  MUX2_X1 DP_reg_pipe00_U25 ( .A(DP_pipe00[13]), .B(DP_w_13_), .S(1'b1), .Z(
        DP_reg_pipe00_n46) );
  MUX2_X1 DP_reg_pipe00_U24 ( .A(DP_pipe00[12]), .B(DP_w_12_), .S(1'b1), .Z(
        DP_reg_pipe00_n47) );
  MUX2_X1 DP_reg_pipe00_U23 ( .A(DP_pipe00[11]), .B(DP_w_11_), .S(1'b1), .Z(
        DP_reg_pipe00_n48) );
  MUX2_X1 DP_reg_pipe00_U22 ( .A(DP_pipe00[10]), .B(DP_w_10_), .S(1'b1), .Z(
        DP_reg_pipe00_n60) );
  MUX2_X1 DP_reg_pipe00_U21 ( .A(DP_pipe00[9]), .B(DP_w_9_), .S(1'b1), .Z(
        DP_reg_pipe00_n61) );
  MUX2_X1 DP_reg_pipe00_U20 ( .A(DP_reg_pipe00_n14), .B(DP_w_8_), .S(1'b1), 
        .Z(DP_reg_pipe00_n62) );
  INV_X1 DP_reg_pipe00_U19 ( .A(DP_reg_pipe00_n71), .ZN(DP_reg_pipe00_n14) );
  MUX2_X1 DP_reg_pipe00_U18 ( .A(DP_reg_pipe00_n13), .B(DP_w_7_), .S(1'b1), 
        .Z(DP_reg_pipe00_n63) );
  INV_X1 DP_reg_pipe00_U17 ( .A(DP_reg_pipe00_n72), .ZN(DP_reg_pipe00_n13) );
  MUX2_X1 DP_reg_pipe00_U16 ( .A(DP_reg_pipe00_n12), .B(DP_w_6_), .S(1'b1), 
        .Z(DP_reg_pipe00_n64) );
  INV_X1 DP_reg_pipe00_U15 ( .A(DP_reg_pipe00_n73), .ZN(DP_reg_pipe00_n12) );
  MUX2_X1 DP_reg_pipe00_U14 ( .A(DP_reg_pipe00_n11), .B(DP_w_5_), .S(1'b1), 
        .Z(DP_reg_pipe00_n65) );
  INV_X1 DP_reg_pipe00_U13 ( .A(DP_reg_pipe00_n74), .ZN(DP_reg_pipe00_n11) );
  MUX2_X1 DP_reg_pipe00_U12 ( .A(DP_reg_pipe00_n10), .B(DP_w_4_), .S(1'b1), 
        .Z(DP_reg_pipe00_n66) );
  INV_X1 DP_reg_pipe00_U11 ( .A(DP_reg_pipe00_n75), .ZN(DP_reg_pipe00_n10) );
  MUX2_X1 DP_reg_pipe00_U10 ( .A(DP_reg_pipe00_n9), .B(DP_w_3_), .S(1'b1), .Z(
        DP_reg_pipe00_n67) );
  INV_X1 DP_reg_pipe00_U9 ( .A(DP_reg_pipe00_n76), .ZN(DP_reg_pipe00_n9) );
  MUX2_X1 DP_reg_pipe00_U8 ( .A(DP_reg_pipe00_n8), .B(DP_w_2_), .S(1'b1), .Z(
        DP_reg_pipe00_n68) );
  INV_X1 DP_reg_pipe00_U7 ( .A(DP_reg_pipe00_n77), .ZN(DP_reg_pipe00_n8) );
  MUX2_X1 DP_reg_pipe00_U6 ( .A(DP_reg_pipe00_n7), .B(DP_w_1_), .S(1'b1), .Z(
        DP_reg_pipe00_n69) );
  INV_X1 DP_reg_pipe00_U5 ( .A(DP_reg_pipe00_n78), .ZN(DP_reg_pipe00_n7) );
  MUX2_X1 DP_reg_pipe00_U4 ( .A(DP_pipe00[0]), .B(DP_w_0_), .S(1'b1), .Z(
        DP_reg_pipe00_n70) );
  BUF_X1 DP_reg_pipe00_U3 ( .A(DP_n8), .Z(DP_reg_pipe00_n4) );
  BUF_X1 DP_reg_pipe00_U2 ( .A(DP_n8), .Z(DP_reg_pipe00_n5) );
  DFFR_X2 DP_reg_pipe00_Q_reg_0_ ( .D(DP_reg_pipe00_n70), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[0]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_11_ ( .D(DP_reg_pipe00_n48), .CK(clk), .RN(DP_n8), .Q(DP_pipe00[11]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_9_ ( .D(DP_reg_pipe00_n61), .CK(clk), .RN(DP_n8), 
        .Q(DP_pipe00[9]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_1_ ( .D(DP_reg_pipe00_n69), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[1]), .QN(DP_reg_pipe00_n78) );
  DFFR_X1 DP_reg_pipe00_Q_reg_2_ ( .D(DP_reg_pipe00_n68), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[2]), .QN(DP_reg_pipe00_n77) );
  DFFR_X1 DP_reg_pipe00_Q_reg_3_ ( .D(DP_reg_pipe00_n67), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[3]), .QN(DP_reg_pipe00_n76) );
  DFFR_X1 DP_reg_pipe00_Q_reg_4_ ( .D(DP_reg_pipe00_n66), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[4]), .QN(DP_reg_pipe00_n75) );
  DFFR_X1 DP_reg_pipe00_Q_reg_5_ ( .D(DP_reg_pipe00_n65), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[5]), .QN(DP_reg_pipe00_n74) );
  DFFR_X1 DP_reg_pipe00_Q_reg_6_ ( .D(DP_reg_pipe00_n64), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[6]), .QN(DP_reg_pipe00_n73) );
  DFFR_X1 DP_reg_pipe00_Q_reg_7_ ( .D(DP_reg_pipe00_n63), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[7]), .QN(DP_reg_pipe00_n72) );
  DFFR_X1 DP_reg_pipe00_Q_reg_8_ ( .D(DP_reg_pipe00_n62), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[8]), .QN(DP_reg_pipe00_n71) );
  DFFR_X1 DP_reg_pipe00_Q_reg_10_ ( .D(DP_reg_pipe00_n60), .CK(clk), .RN(
        DP_reg_pipe00_n5), .Q(DP_pipe00[10]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_12_ ( .D(DP_reg_pipe00_n47), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[12]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_13_ ( .D(DP_reg_pipe00_n46), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[13]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_14_ ( .D(DP_reg_pipe00_n45), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[14]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_15_ ( .D(DP_reg_pipe00_n44), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[15]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_16_ ( .D(DP_reg_pipe00_n43), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[16]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_17_ ( .D(DP_reg_pipe00_n42), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[17]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_18_ ( .D(DP_reg_pipe00_n41), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[18]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_19_ ( .D(DP_reg_pipe00_n40), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[19]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_20_ ( .D(DP_reg_pipe00_n39), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[20]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_21_ ( .D(DP_reg_pipe00_n38), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[21]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_22_ ( .D(DP_reg_pipe00_n37), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[22]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_23_ ( .D(DP_reg_pipe00_n36), .CK(clk), .RN(
        DP_reg_pipe00_n4), .Q(DP_pipe00[23]) );
  MUX2_X1 DP_reg_pipe01_U46 ( .A(DP_reg_pipe01_n29), .B(DP_sw0_23_), .S(1'b1), 
        .Z(DP_reg_pipe01_n36) );
  INV_X1 DP_reg_pipe01_U45 ( .A(DP_reg_pipe01_n93), .ZN(DP_reg_pipe01_n29) );
  MUX2_X1 DP_reg_pipe01_U44 ( .A(DP_reg_pipe01_n27), .B(DP_sw0_22_), .S(1'b1), 
        .Z(DP_reg_pipe01_n38) );
  INV_X1 DP_reg_pipe01_U43 ( .A(DP_reg_pipe01_n94), .ZN(DP_reg_pipe01_n27) );
  MUX2_X1 DP_reg_pipe01_U42 ( .A(DP_reg_pipe01_n25), .B(DP_sw0_21_), .S(1'b1), 
        .Z(DP_reg_pipe01_n71) );
  INV_X1 DP_reg_pipe01_U41 ( .A(DP_reg_pipe01_n95), .ZN(DP_reg_pipe01_n25) );
  MUX2_X1 DP_reg_pipe01_U40 ( .A(DP_reg_pipe01_n24), .B(DP_sw0_20_), .S(1'b1), 
        .Z(DP_reg_pipe01_n72) );
  INV_X1 DP_reg_pipe01_U39 ( .A(DP_reg_pipe01_n96), .ZN(DP_reg_pipe01_n24) );
  MUX2_X1 DP_reg_pipe01_U38 ( .A(DP_reg_pipe01_n23), .B(DP_sw0_19_), .S(1'b1), 
        .Z(DP_reg_pipe01_n73) );
  INV_X1 DP_reg_pipe01_U37 ( .A(DP_reg_pipe01_n97), .ZN(DP_reg_pipe01_n23) );
  MUX2_X1 DP_reg_pipe01_U36 ( .A(DP_reg_pipe01_n22), .B(DP_sw0_18_), .S(1'b1), 
        .Z(DP_reg_pipe01_n74) );
  INV_X1 DP_reg_pipe01_U35 ( .A(DP_reg_pipe01_n98), .ZN(DP_reg_pipe01_n22) );
  MUX2_X1 DP_reg_pipe01_U34 ( .A(DP_reg_pipe01_n21), .B(DP_sw0_17_), .S(1'b1), 
        .Z(DP_reg_pipe01_n75) );
  INV_X1 DP_reg_pipe01_U33 ( .A(DP_reg_pipe01_n99), .ZN(DP_reg_pipe01_n21) );
  MUX2_X1 DP_reg_pipe01_U32 ( .A(DP_reg_pipe01_n20), .B(DP_sw0_16_), .S(1'b1), 
        .Z(DP_reg_pipe01_n76) );
  INV_X1 DP_reg_pipe01_U31 ( .A(DP_reg_pipe01_n100), .ZN(DP_reg_pipe01_n20) );
  MUX2_X1 DP_reg_pipe01_U30 ( .A(DP_reg_pipe01_n19), .B(DP_sw0_15_), .S(1'b1), 
        .Z(DP_reg_pipe01_n77) );
  INV_X1 DP_reg_pipe01_U29 ( .A(DP_reg_pipe01_n101), .ZN(DP_reg_pipe01_n19) );
  MUX2_X1 DP_reg_pipe01_U28 ( .A(DP_reg_pipe01_n18), .B(DP_sw0_14_), .S(1'b1), 
        .Z(DP_reg_pipe01_n78) );
  INV_X1 DP_reg_pipe01_U27 ( .A(DP_reg_pipe01_n102), .ZN(DP_reg_pipe01_n18) );
  MUX2_X1 DP_reg_pipe01_U26 ( .A(DP_pipe01[13]), .B(DP_sw0_13_), .S(1'b1), .Z(
        DP_reg_pipe01_n79) );
  MUX2_X1 DP_reg_pipe01_U25 ( .A(DP_reg_pipe01_n17), .B(DP_sw0_12_), .S(1'b1), 
        .Z(DP_reg_pipe01_n80) );
  INV_X1 DP_reg_pipe01_U24 ( .A(DP_reg_pipe01_n103), .ZN(DP_reg_pipe01_n17) );
  MUX2_X1 DP_reg_pipe01_U23 ( .A(DP_pipe01[11]), .B(DP_sw0_11_), .S(1'b1), .Z(
        DP_reg_pipe01_n81) );
  MUX2_X1 DP_reg_pipe01_U22 ( .A(DP_reg_pipe01_n16), .B(DP_sw0_10_), .S(1'b1), 
        .Z(DP_reg_pipe01_n82) );
  INV_X1 DP_reg_pipe01_U21 ( .A(DP_reg_pipe01_n104), .ZN(DP_reg_pipe01_n16) );
  MUX2_X1 DP_reg_pipe01_U20 ( .A(DP_reg_pipe01_n15), .B(DP_sw0_9_), .S(1'b1), 
        .Z(DP_reg_pipe01_n83) );
  INV_X1 DP_reg_pipe01_U19 ( .A(DP_reg_pipe01_n105), .ZN(DP_reg_pipe01_n15) );
  MUX2_X1 DP_reg_pipe01_U18 ( .A(DP_reg_pipe01_n14), .B(DP_sw0_8_), .S(1'b1), 
        .Z(DP_reg_pipe01_n84) );
  INV_X1 DP_reg_pipe01_U17 ( .A(DP_reg_pipe01_n106), .ZN(DP_reg_pipe01_n14) );
  MUX2_X1 DP_reg_pipe01_U16 ( .A(DP_reg_pipe01_n13), .B(DP_sw0_7_), .S(1'b1), 
        .Z(DP_reg_pipe01_n85) );
  INV_X1 DP_reg_pipe01_U15 ( .A(DP_reg_pipe01_n107), .ZN(DP_reg_pipe01_n13) );
  MUX2_X1 DP_reg_pipe01_U14 ( .A(DP_reg_pipe01_n12), .B(DP_sw0_6_), .S(1'b1), 
        .Z(DP_reg_pipe01_n86) );
  INV_X1 DP_reg_pipe01_U13 ( .A(DP_reg_pipe01_n108), .ZN(DP_reg_pipe01_n12) );
  MUX2_X1 DP_reg_pipe01_U12 ( .A(DP_reg_pipe01_n11), .B(DP_sw0_5_), .S(1'b1), 
        .Z(DP_reg_pipe01_n87) );
  INV_X1 DP_reg_pipe01_U11 ( .A(DP_reg_pipe01_n109), .ZN(DP_reg_pipe01_n11) );
  MUX2_X1 DP_reg_pipe01_U10 ( .A(DP_pipe01[4]), .B(DP_sw0_4_), .S(1'b1), .Z(
        DP_reg_pipe01_n88) );
  MUX2_X1 DP_reg_pipe01_U9 ( .A(DP_reg_pipe01_n9), .B(DP_sw0_3_), .S(1'b1), 
        .Z(DP_reg_pipe01_n89) );
  INV_X1 DP_reg_pipe01_U8 ( .A(DP_reg_pipe01_n110), .ZN(DP_reg_pipe01_n9) );
  MUX2_X1 DP_reg_pipe01_U7 ( .A(DP_pipe01[2]), .B(DP_sw0_2_), .S(1'b1), .Z(
        DP_reg_pipe01_n90) );
  MUX2_X1 DP_reg_pipe01_U6 ( .A(DP_reg_pipe01_n7), .B(DP_sw0_1_), .S(1'b1), 
        .Z(DP_reg_pipe01_n91) );
  INV_X1 DP_reg_pipe01_U5 ( .A(DP_reg_pipe01_n111), .ZN(DP_reg_pipe01_n7) );
  MUX2_X1 DP_reg_pipe01_U4 ( .A(DP_pipe01[0]), .B(DP_sw0_0_), .S(1'b1), .Z(
        DP_reg_pipe01_n92) );
  BUF_X1 DP_reg_pipe01_U3 ( .A(DP_n7), .Z(DP_reg_pipe01_n4) );
  BUF_X1 DP_reg_pipe01_U2 ( .A(DP_n7), .Z(DP_reg_pipe01_n5) );
  DFFR_X2 DP_reg_pipe01_Q_reg_0_ ( .D(DP_reg_pipe01_n92), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[0]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_13_ ( .D(DP_reg_pipe01_n79), .CK(clk), .RN(DP_n7), .Q(DP_pipe01[13]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_11_ ( .D(DP_reg_pipe01_n81), .CK(clk), .RN(DP_n7), .Q(DP_pipe01[11]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_1_ ( .D(DP_reg_pipe01_n91), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[1]), .QN(DP_reg_pipe01_n111) );
  DFFR_X1 DP_reg_pipe01_Q_reg_2_ ( .D(DP_reg_pipe01_n90), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[2]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_3_ ( .D(DP_reg_pipe01_n89), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[3]), .QN(DP_reg_pipe01_n110) );
  DFFR_X1 DP_reg_pipe01_Q_reg_4_ ( .D(DP_reg_pipe01_n88), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[4]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_5_ ( .D(DP_reg_pipe01_n87), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[5]), .QN(DP_reg_pipe01_n109) );
  DFFR_X1 DP_reg_pipe01_Q_reg_6_ ( .D(DP_reg_pipe01_n86), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[6]), .QN(DP_reg_pipe01_n108) );
  DFFR_X1 DP_reg_pipe01_Q_reg_7_ ( .D(DP_reg_pipe01_n85), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[7]), .QN(DP_reg_pipe01_n107) );
  DFFR_X1 DP_reg_pipe01_Q_reg_8_ ( .D(DP_reg_pipe01_n84), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[8]), .QN(DP_reg_pipe01_n106) );
  DFFR_X1 DP_reg_pipe01_Q_reg_9_ ( .D(DP_reg_pipe01_n83), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[9]), .QN(DP_reg_pipe01_n105) );
  DFFR_X1 DP_reg_pipe01_Q_reg_10_ ( .D(DP_reg_pipe01_n82), .CK(clk), .RN(
        DP_reg_pipe01_n5), .Q(DP_pipe01[10]), .QN(DP_reg_pipe01_n104) );
  DFFR_X1 DP_reg_pipe01_Q_reg_12_ ( .D(DP_reg_pipe01_n80), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[12]), .QN(DP_reg_pipe01_n103) );
  DFFR_X1 DP_reg_pipe01_Q_reg_14_ ( .D(DP_reg_pipe01_n78), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[14]), .QN(DP_reg_pipe01_n102) );
  DFFR_X1 DP_reg_pipe01_Q_reg_15_ ( .D(DP_reg_pipe01_n77), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[15]), .QN(DP_reg_pipe01_n101) );
  DFFR_X1 DP_reg_pipe01_Q_reg_16_ ( .D(DP_reg_pipe01_n76), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[16]), .QN(DP_reg_pipe01_n100) );
  DFFR_X1 DP_reg_pipe01_Q_reg_17_ ( .D(DP_reg_pipe01_n75), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[17]), .QN(DP_reg_pipe01_n99) );
  DFFR_X1 DP_reg_pipe01_Q_reg_18_ ( .D(DP_reg_pipe01_n74), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[18]), .QN(DP_reg_pipe01_n98) );
  DFFR_X1 DP_reg_pipe01_Q_reg_19_ ( .D(DP_reg_pipe01_n73), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[19]), .QN(DP_reg_pipe01_n97) );
  DFFR_X1 DP_reg_pipe01_Q_reg_20_ ( .D(DP_reg_pipe01_n72), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[20]), .QN(DP_reg_pipe01_n96) );
  DFFR_X1 DP_reg_pipe01_Q_reg_21_ ( .D(DP_reg_pipe01_n71), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[21]), .QN(DP_reg_pipe01_n95) );
  DFFR_X1 DP_reg_pipe01_Q_reg_22_ ( .D(DP_reg_pipe01_n38), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[22]), .QN(DP_reg_pipe01_n94) );
  DFFR_X1 DP_reg_pipe01_Q_reg_23_ ( .D(DP_reg_pipe01_n36), .CK(clk), .RN(
        DP_reg_pipe01_n4), .Q(DP_pipe01[23]), .QN(DP_reg_pipe01_n93) );
  MUX2_X1 DP_reg_pipe02_U47 ( .A(DP_reg_pipe02_n32), .B(DP_sw1_23_), .S(1'b1), 
        .Z(DP_reg_pipe02_n39) );
  INV_X1 DP_reg_pipe02_U46 ( .A(DP_reg_pipe02_n95), .ZN(DP_reg_pipe02_n32) );
  MUX2_X1 DP_reg_pipe02_U45 ( .A(DP_reg_pipe02_n27), .B(DP_sw1_22_), .S(1'b1), 
        .Z(DP_reg_pipe02_n72) );
  INV_X1 DP_reg_pipe02_U44 ( .A(DP_reg_pipe02_n96), .ZN(DP_reg_pipe02_n27) );
  MUX2_X1 DP_reg_pipe02_U43 ( .A(DP_reg_pipe02_n25), .B(DP_sw1_21_), .S(1'b1), 
        .Z(DP_reg_pipe02_n73) );
  INV_X1 DP_reg_pipe02_U42 ( .A(DP_reg_pipe02_n97), .ZN(DP_reg_pipe02_n25) );
  MUX2_X1 DP_reg_pipe02_U41 ( .A(DP_reg_pipe02_n24), .B(DP_sw1_20_), .S(1'b1), 
        .Z(DP_reg_pipe02_n74) );
  INV_X1 DP_reg_pipe02_U40 ( .A(DP_reg_pipe02_n98), .ZN(DP_reg_pipe02_n24) );
  MUX2_X1 DP_reg_pipe02_U39 ( .A(DP_reg_pipe02_n23), .B(DP_sw1_19_), .S(1'b1), 
        .Z(DP_reg_pipe02_n75) );
  INV_X1 DP_reg_pipe02_U38 ( .A(DP_reg_pipe02_n99), .ZN(DP_reg_pipe02_n23) );
  MUX2_X1 DP_reg_pipe02_U37 ( .A(DP_reg_pipe02_n22), .B(DP_sw1_18_), .S(1'b1), 
        .Z(DP_reg_pipe02_n76) );
  INV_X1 DP_reg_pipe02_U36 ( .A(DP_reg_pipe02_n100), .ZN(DP_reg_pipe02_n22) );
  MUX2_X1 DP_reg_pipe02_U35 ( .A(DP_reg_pipe02_n21), .B(DP_sw1_17_), .S(1'b1), 
        .Z(DP_reg_pipe02_n77) );
  INV_X1 DP_reg_pipe02_U34 ( .A(DP_reg_pipe02_n101), .ZN(DP_reg_pipe02_n21) );
  MUX2_X1 DP_reg_pipe02_U33 ( .A(DP_reg_pipe02_n20), .B(DP_sw1_16_), .S(1'b1), 
        .Z(DP_reg_pipe02_n78) );
  INV_X1 DP_reg_pipe02_U32 ( .A(DP_reg_pipe02_n102), .ZN(DP_reg_pipe02_n20) );
  MUX2_X1 DP_reg_pipe02_U31 ( .A(DP_reg_pipe02_n19), .B(DP_sw1_15_), .S(1'b1), 
        .Z(DP_reg_pipe02_n79) );
  INV_X1 DP_reg_pipe02_U30 ( .A(DP_reg_pipe02_n103), .ZN(DP_reg_pipe02_n19) );
  MUX2_X1 DP_reg_pipe02_U29 ( .A(DP_pipe02[14]), .B(DP_sw1_14_), .S(1'b1), .Z(
        DP_reg_pipe02_n80) );
  MUX2_X1 DP_reg_pipe02_U28 ( .A(DP_reg_pipe02_n17), .B(DP_sw1_13_), .S(1'b1), 
        .Z(DP_reg_pipe02_n81) );
  INV_X1 DP_reg_pipe02_U27 ( .A(DP_reg_pipe02_n104), .ZN(DP_reg_pipe02_n17) );
  MUX2_X1 DP_reg_pipe02_U26 ( .A(DP_reg_pipe02_n16), .B(DP_sw1_12_), .S(1'b1), 
        .Z(DP_reg_pipe02_n82) );
  INV_X1 DP_reg_pipe02_U25 ( .A(DP_reg_pipe02_n105), .ZN(DP_reg_pipe02_n16) );
  MUX2_X1 DP_reg_pipe02_U24 ( .A(DP_reg_pipe02_n15), .B(DP_sw1_11_), .S(1'b1), 
        .Z(DP_reg_pipe02_n83) );
  INV_X1 DP_reg_pipe02_U23 ( .A(DP_reg_pipe02_n106), .ZN(DP_reg_pipe02_n15) );
  MUX2_X1 DP_reg_pipe02_U22 ( .A(DP_reg_pipe02_n14), .B(DP_sw1_10_), .S(1'b1), 
        .Z(DP_reg_pipe02_n84) );
  INV_X1 DP_reg_pipe02_U21 ( .A(DP_reg_pipe02_n107), .ZN(DP_reg_pipe02_n14) );
  MUX2_X1 DP_reg_pipe02_U20 ( .A(DP_reg_pipe02_n13), .B(DP_sw1_9_), .S(1'b1), 
        .Z(DP_reg_pipe02_n85) );
  INV_X1 DP_reg_pipe02_U19 ( .A(DP_reg_pipe02_n108), .ZN(DP_reg_pipe02_n13) );
  MUX2_X1 DP_reg_pipe02_U18 ( .A(DP_reg_pipe02_n12), .B(DP_sw1_8_), .S(1'b1), 
        .Z(DP_reg_pipe02_n86) );
  INV_X1 DP_reg_pipe02_U17 ( .A(DP_reg_pipe02_n109), .ZN(DP_reg_pipe02_n12) );
  MUX2_X1 DP_reg_pipe02_U16 ( .A(DP_pipe02[7]), .B(DP_sw1_7_), .S(1'b1), .Z(
        DP_reg_pipe02_n87) );
  MUX2_X1 DP_reg_pipe02_U15 ( .A(DP_reg_pipe02_n10), .B(DP_sw1_6_), .S(1'b1), 
        .Z(DP_reg_pipe02_n88) );
  INV_X1 DP_reg_pipe02_U14 ( .A(DP_reg_pipe02_n110), .ZN(DP_reg_pipe02_n10) );
  MUX2_X1 DP_reg_pipe02_U13 ( .A(DP_reg_pipe02_n9), .B(DP_sw1_5_), .S(1'b1), 
        .Z(DP_reg_pipe02_n89) );
  INV_X1 DP_reg_pipe02_U12 ( .A(DP_reg_pipe02_n111), .ZN(DP_reg_pipe02_n9) );
  MUX2_X1 DP_reg_pipe02_U11 ( .A(DP_reg_pipe02_n8), .B(DP_sw1_4_), .S(1'b1), 
        .Z(DP_reg_pipe02_n90) );
  INV_X1 DP_reg_pipe02_U10 ( .A(DP_reg_pipe02_n112), .ZN(DP_reg_pipe02_n8) );
  MUX2_X1 DP_reg_pipe02_U9 ( .A(DP_reg_pipe02_n7), .B(DP_sw1_3_), .S(1'b1), 
        .Z(DP_reg_pipe02_n91) );
  INV_X1 DP_reg_pipe02_U8 ( .A(DP_reg_pipe02_n113), .ZN(DP_reg_pipe02_n7) );
  MUX2_X1 DP_reg_pipe02_U7 ( .A(DP_pipe02[2]), .B(DP_sw1_2_), .S(1'b1), .Z(
        DP_reg_pipe02_n92) );
  MUX2_X1 DP_reg_pipe02_U6 ( .A(DP_reg_pipe02_n5), .B(DP_sw1_1_), .S(1'b1), 
        .Z(DP_reg_pipe02_n93) );
  INV_X1 DP_reg_pipe02_U5 ( .A(DP_reg_pipe02_n114), .ZN(DP_reg_pipe02_n5) );
  MUX2_X1 DP_reg_pipe02_U4 ( .A(DP_pipe02[0]), .B(DP_sw1_0_), .S(1'b1), .Z(
        DP_reg_pipe02_n94) );
  BUF_X1 DP_reg_pipe02_U3 ( .A(DP_n7), .Z(DP_reg_pipe02_n2) );
  BUF_X1 DP_reg_pipe02_U2 ( .A(DP_n7), .Z(DP_reg_pipe02_n3) );
  DFFR_X2 DP_reg_pipe02_Q_reg_0_ ( .D(DP_reg_pipe02_n94), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[0]) );
  DFFR_X1 DP_reg_pipe02_Q_reg_1_ ( .D(DP_reg_pipe02_n93), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[1]), .QN(DP_reg_pipe02_n114) );
  DFFR_X1 DP_reg_pipe02_Q_reg_2_ ( .D(DP_reg_pipe02_n92), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[2]) );
  DFFR_X1 DP_reg_pipe02_Q_reg_3_ ( .D(DP_reg_pipe02_n91), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[3]), .QN(DP_reg_pipe02_n113) );
  DFFR_X1 DP_reg_pipe02_Q_reg_4_ ( .D(DP_reg_pipe02_n90), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[4]), .QN(DP_reg_pipe02_n112) );
  DFFR_X1 DP_reg_pipe02_Q_reg_5_ ( .D(DP_reg_pipe02_n89), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[5]), .QN(DP_reg_pipe02_n111) );
  DFFR_X1 DP_reg_pipe02_Q_reg_6_ ( .D(DP_reg_pipe02_n88), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[6]), .QN(DP_reg_pipe02_n110) );
  DFFR_X1 DP_reg_pipe02_Q_reg_7_ ( .D(DP_reg_pipe02_n87), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[7]) );
  DFFR_X1 DP_reg_pipe02_Q_reg_8_ ( .D(DP_reg_pipe02_n86), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[8]), .QN(DP_reg_pipe02_n109) );
  DFFR_X1 DP_reg_pipe02_Q_reg_9_ ( .D(DP_reg_pipe02_n85), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[9]), .QN(DP_reg_pipe02_n108) );
  DFFR_X1 DP_reg_pipe02_Q_reg_10_ ( .D(DP_reg_pipe02_n84), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[10]), .QN(DP_reg_pipe02_n107) );
  DFFR_X1 DP_reg_pipe02_Q_reg_11_ ( .D(DP_reg_pipe02_n83), .CK(clk), .RN(
        DP_reg_pipe02_n3), .Q(DP_pipe02[11]), .QN(DP_reg_pipe02_n106) );
  DFFR_X1 DP_reg_pipe02_Q_reg_12_ ( .D(DP_reg_pipe02_n82), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[12]), .QN(DP_reg_pipe02_n105) );
  DFFR_X1 DP_reg_pipe02_Q_reg_13_ ( .D(DP_reg_pipe02_n81), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[13]), .QN(DP_reg_pipe02_n104) );
  DFFR_X1 DP_reg_pipe02_Q_reg_14_ ( .D(DP_reg_pipe02_n80), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[14]) );
  DFFR_X1 DP_reg_pipe02_Q_reg_15_ ( .D(DP_reg_pipe02_n79), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[15]), .QN(DP_reg_pipe02_n103) );
  DFFR_X1 DP_reg_pipe02_Q_reg_16_ ( .D(DP_reg_pipe02_n78), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[16]), .QN(DP_reg_pipe02_n102) );
  DFFR_X1 DP_reg_pipe02_Q_reg_17_ ( .D(DP_reg_pipe02_n77), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[17]), .QN(DP_reg_pipe02_n101) );
  DFFR_X1 DP_reg_pipe02_Q_reg_18_ ( .D(DP_reg_pipe02_n76), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[18]), .QN(DP_reg_pipe02_n100) );
  DFFR_X1 DP_reg_pipe02_Q_reg_19_ ( .D(DP_reg_pipe02_n75), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[19]), .QN(DP_reg_pipe02_n99) );
  DFFR_X1 DP_reg_pipe02_Q_reg_20_ ( .D(DP_reg_pipe02_n74), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[20]), .QN(DP_reg_pipe02_n98) );
  DFFR_X1 DP_reg_pipe02_Q_reg_21_ ( .D(DP_reg_pipe02_n73), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[21]), .QN(DP_reg_pipe02_n97) );
  DFFR_X1 DP_reg_pipe02_Q_reg_22_ ( .D(DP_reg_pipe02_n72), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[22]), .QN(DP_reg_pipe02_n96) );
  DFFR_X1 DP_reg_pipe02_Q_reg_23_ ( .D(DP_reg_pipe02_n39), .CK(clk), .RN(
        DP_reg_pipe02_n2), .Q(DP_pipe02[23]), .QN(DP_reg_pipe02_n95) );
  MUX2_X1 DP_reg_pipe03_U47 ( .A(DP_reg_pipe03_n34), .B(DP_sw2[23]), .S(1'b1), 
        .Z(DP_reg_pipe03_n39) );
  INV_X1 DP_reg_pipe03_U46 ( .A(DP_reg_pipe03_n95), .ZN(DP_reg_pipe03_n34) );
  MUX2_X1 DP_reg_pipe03_U45 ( .A(DP_reg_pipe03_n33), .B(DP_sw2[22]), .S(1'b1), 
        .Z(DP_reg_pipe03_n72) );
  INV_X1 DP_reg_pipe03_U44 ( .A(DP_reg_pipe03_n96), .ZN(DP_reg_pipe03_n33) );
  MUX2_X1 DP_reg_pipe03_U43 ( .A(DP_reg_pipe03_n27), .B(DP_sw2[21]), .S(1'b1), 
        .Z(DP_reg_pipe03_n73) );
  INV_X1 DP_reg_pipe03_U42 ( .A(DP_reg_pipe03_n97), .ZN(DP_reg_pipe03_n27) );
  MUX2_X1 DP_reg_pipe03_U41 ( .A(DP_reg_pipe03_n25), .B(DP_sw2[20]), .S(1'b1), 
        .Z(DP_reg_pipe03_n74) );
  INV_X1 DP_reg_pipe03_U40 ( .A(DP_reg_pipe03_n98), .ZN(DP_reg_pipe03_n25) );
  MUX2_X1 DP_reg_pipe03_U39 ( .A(DP_reg_pipe03_n24), .B(DP_sw2[19]), .S(1'b1), 
        .Z(DP_reg_pipe03_n75) );
  INV_X1 DP_reg_pipe03_U38 ( .A(DP_reg_pipe03_n99), .ZN(DP_reg_pipe03_n24) );
  MUX2_X1 DP_reg_pipe03_U37 ( .A(DP_reg_pipe03_n23), .B(DP_sw2[18]), .S(1'b1), 
        .Z(DP_reg_pipe03_n76) );
  INV_X1 DP_reg_pipe03_U36 ( .A(DP_reg_pipe03_n100), .ZN(DP_reg_pipe03_n23) );
  MUX2_X1 DP_reg_pipe03_U35 ( .A(DP_reg_pipe03_n22), .B(DP_sw2[17]), .S(1'b1), 
        .Z(DP_reg_pipe03_n77) );
  INV_X1 DP_reg_pipe03_U34 ( .A(DP_reg_pipe03_n101), .ZN(DP_reg_pipe03_n22) );
  MUX2_X1 DP_reg_pipe03_U33 ( .A(DP_reg_pipe03_n21), .B(DP_sw2[16]), .S(1'b1), 
        .Z(DP_reg_pipe03_n78) );
  INV_X1 DP_reg_pipe03_U32 ( .A(DP_reg_pipe03_n102), .ZN(DP_reg_pipe03_n21) );
  MUX2_X1 DP_reg_pipe03_U31 ( .A(DP_reg_pipe03_n20), .B(DP_sw2[15]), .S(1'b1), 
        .Z(DP_reg_pipe03_n79) );
  INV_X1 DP_reg_pipe03_U30 ( .A(DP_reg_pipe03_n103), .ZN(DP_reg_pipe03_n20) );
  MUX2_X1 DP_reg_pipe03_U29 ( .A(DP_pipe03[14]), .B(DP_sw2[14]), .S(1'b1), .Z(
        DP_reg_pipe03_n80) );
  MUX2_X1 DP_reg_pipe03_U28 ( .A(DP_reg_pipe03_n18), .B(DP_sw2[13]), .S(1'b1), 
        .Z(DP_reg_pipe03_n81) );
  INV_X1 DP_reg_pipe03_U27 ( .A(DP_reg_pipe03_n104), .ZN(DP_reg_pipe03_n18) );
  MUX2_X1 DP_reg_pipe03_U26 ( .A(DP_reg_pipe03_n17), .B(DP_sw2[12]), .S(1'b1), 
        .Z(DP_reg_pipe03_n82) );
  INV_X1 DP_reg_pipe03_U25 ( .A(DP_reg_pipe03_n105), .ZN(DP_reg_pipe03_n17) );
  MUX2_X1 DP_reg_pipe03_U24 ( .A(DP_reg_pipe03_n16), .B(DP_sw2[11]), .S(1'b1), 
        .Z(DP_reg_pipe03_n83) );
  INV_X1 DP_reg_pipe03_U23 ( .A(DP_reg_pipe03_n106), .ZN(DP_reg_pipe03_n16) );
  MUX2_X1 DP_reg_pipe03_U22 ( .A(DP_reg_pipe03_n15), .B(DP_sw2[10]), .S(1'b1), 
        .Z(DP_reg_pipe03_n84) );
  INV_X1 DP_reg_pipe03_U21 ( .A(DP_reg_pipe03_n107), .ZN(DP_reg_pipe03_n15) );
  MUX2_X1 DP_reg_pipe03_U20 ( .A(DP_pipe03[9]), .B(DP_sw2[9]), .S(1'b1), .Z(
        DP_reg_pipe03_n85) );
  MUX2_X1 DP_reg_pipe03_U19 ( .A(DP_pipe03[8]), .B(DP_sw2[8]), .S(1'b1), .Z(
        DP_reg_pipe03_n86) );
  MUX2_X1 DP_reg_pipe03_U18 ( .A(DP_reg_pipe03_n12), .B(DP_sw2[7]), .S(1'b1), 
        .Z(DP_reg_pipe03_n87) );
  INV_X1 DP_reg_pipe03_U17 ( .A(DP_reg_pipe03_n108), .ZN(DP_reg_pipe03_n12) );
  MUX2_X1 DP_reg_pipe03_U16 ( .A(DP_reg_pipe03_n11), .B(DP_sw2[6]), .S(1'b1), 
        .Z(DP_reg_pipe03_n88) );
  INV_X1 DP_reg_pipe03_U15 ( .A(DP_reg_pipe03_n109), .ZN(DP_reg_pipe03_n11) );
  MUX2_X1 DP_reg_pipe03_U14 ( .A(DP_reg_pipe03_n10), .B(DP_sw2[5]), .S(1'b1), 
        .Z(DP_reg_pipe03_n89) );
  INV_X1 DP_reg_pipe03_U13 ( .A(DP_reg_pipe03_n110), .ZN(DP_reg_pipe03_n10) );
  MUX2_X1 DP_reg_pipe03_U12 ( .A(DP_reg_pipe03_n9), .B(DP_sw2[4]), .S(1'b1), 
        .Z(DP_reg_pipe03_n90) );
  INV_X1 DP_reg_pipe03_U11 ( .A(DP_reg_pipe03_n111), .ZN(DP_reg_pipe03_n9) );
  MUX2_X1 DP_reg_pipe03_U10 ( .A(DP_reg_pipe03_n8), .B(DP_sw2[3]), .S(1'b1), 
        .Z(DP_reg_pipe03_n91) );
  INV_X1 DP_reg_pipe03_U9 ( .A(DP_reg_pipe03_n112), .ZN(DP_reg_pipe03_n8) );
  MUX2_X1 DP_reg_pipe03_U8 ( .A(DP_pipe03[2]), .B(DP_sw2[2]), .S(1'b1), .Z(
        DP_reg_pipe03_n92) );
  MUX2_X1 DP_reg_pipe03_U7 ( .A(DP_reg_pipe03_n6), .B(DP_sw2[1]), .S(1'b1), 
        .Z(DP_reg_pipe03_n93) );
  INV_X1 DP_reg_pipe03_U6 ( .A(DP_reg_pipe03_n113), .ZN(DP_reg_pipe03_n6) );
  MUX2_X1 DP_reg_pipe03_U5 ( .A(DP_reg_pipe03_n5), .B(DP_sw2[0]), .S(1'b1), 
        .Z(DP_reg_pipe03_n94) );
  BUF_X1 DP_reg_pipe03_U4 ( .A(DP_n6), .Z(DP_reg_pipe03_n3) );
  BUF_X1 DP_reg_pipe03_U3 ( .A(DP_n6), .Z(DP_reg_pipe03_n4) );
  INV_X2 DP_reg_pipe03_U2 ( .A(DP_reg_pipe03_n1), .ZN(DP_pipe03[0]) );
  DFFR_X1 DP_reg_pipe03_Q_reg_0_ ( .D(DP_reg_pipe03_n94), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_reg_pipe03_n5), .QN(DP_reg_pipe03_n1) );
  DFFR_X1 DP_reg_pipe03_Q_reg_1_ ( .D(DP_reg_pipe03_n93), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[1]), .QN(DP_reg_pipe03_n113) );
  DFFR_X1 DP_reg_pipe03_Q_reg_2_ ( .D(DP_reg_pipe03_n92), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[2]) );
  DFFR_X1 DP_reg_pipe03_Q_reg_3_ ( .D(DP_reg_pipe03_n91), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[3]), .QN(DP_reg_pipe03_n112) );
  DFFR_X1 DP_reg_pipe03_Q_reg_4_ ( .D(DP_reg_pipe03_n90), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[4]), .QN(DP_reg_pipe03_n111) );
  DFFR_X1 DP_reg_pipe03_Q_reg_5_ ( .D(DP_reg_pipe03_n89), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[5]), .QN(DP_reg_pipe03_n110) );
  DFFR_X1 DP_reg_pipe03_Q_reg_6_ ( .D(DP_reg_pipe03_n88), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[6]), .QN(DP_reg_pipe03_n109) );
  DFFR_X1 DP_reg_pipe03_Q_reg_7_ ( .D(DP_reg_pipe03_n87), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[7]), .QN(DP_reg_pipe03_n108) );
  DFFR_X1 DP_reg_pipe03_Q_reg_8_ ( .D(DP_reg_pipe03_n86), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[8]) );
  DFFR_X1 DP_reg_pipe03_Q_reg_9_ ( .D(DP_reg_pipe03_n85), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[9]) );
  DFFR_X1 DP_reg_pipe03_Q_reg_10_ ( .D(DP_reg_pipe03_n84), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[10]), .QN(DP_reg_pipe03_n107) );
  DFFR_X1 DP_reg_pipe03_Q_reg_11_ ( .D(DP_reg_pipe03_n83), .CK(clk), .RN(
        DP_reg_pipe03_n4), .Q(DP_pipe03[11]), .QN(DP_reg_pipe03_n106) );
  DFFR_X1 DP_reg_pipe03_Q_reg_12_ ( .D(DP_reg_pipe03_n82), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[12]), .QN(DP_reg_pipe03_n105) );
  DFFR_X1 DP_reg_pipe03_Q_reg_13_ ( .D(DP_reg_pipe03_n81), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[13]), .QN(DP_reg_pipe03_n104) );
  DFFR_X1 DP_reg_pipe03_Q_reg_14_ ( .D(DP_reg_pipe03_n80), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[14]) );
  DFFR_X1 DP_reg_pipe03_Q_reg_15_ ( .D(DP_reg_pipe03_n79), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[15]), .QN(DP_reg_pipe03_n103) );
  DFFR_X1 DP_reg_pipe03_Q_reg_16_ ( .D(DP_reg_pipe03_n78), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[16]), .QN(DP_reg_pipe03_n102) );
  DFFR_X1 DP_reg_pipe03_Q_reg_17_ ( .D(DP_reg_pipe03_n77), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[17]), .QN(DP_reg_pipe03_n101) );
  DFFR_X1 DP_reg_pipe03_Q_reg_18_ ( .D(DP_reg_pipe03_n76), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[18]), .QN(DP_reg_pipe03_n100) );
  DFFR_X1 DP_reg_pipe03_Q_reg_19_ ( .D(DP_reg_pipe03_n75), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[19]), .QN(DP_reg_pipe03_n99) );
  DFFR_X1 DP_reg_pipe03_Q_reg_20_ ( .D(DP_reg_pipe03_n74), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[20]), .QN(DP_reg_pipe03_n98) );
  DFFR_X1 DP_reg_pipe03_Q_reg_21_ ( .D(DP_reg_pipe03_n73), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[21]), .QN(DP_reg_pipe03_n97) );
  DFFR_X1 DP_reg_pipe03_Q_reg_22_ ( .D(DP_reg_pipe03_n72), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[22]), .QN(DP_reg_pipe03_n96) );
  DFFR_X1 DP_reg_pipe03_Q_reg_23_ ( .D(DP_reg_pipe03_n39), .CK(clk), .RN(
        DP_reg_pipe03_n3), .Q(DP_pipe03[23]), .QN(DP_reg_pipe03_n95) );
  MUX2_X1 DP_reg_pipe10_U50 ( .A(DP_pipe10[23]), .B(DP_pipe0_coeff_pipe00[23]), 
        .S(1'b1), .Z(DP_reg_pipe10_n84) );
  NAND2_X1 DP_reg_pipe10_U49 ( .A1(DP_reg_pipe10_n81), .A2(DP_reg_pipe10_n82), 
        .ZN(DP_reg_pipe10_n85) );
  NAND2_X1 DP_reg_pipe10_U48 ( .A1(DP_pipe0_coeff_pipe00[22]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n81) );
  NAND2_X1 DP_reg_pipe10_U47 ( .A1(DP_pipe10[22]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n82) );
  NAND2_X1 DP_reg_pipe10_U46 ( .A1(DP_reg_pipe10_n77), .A2(DP_reg_pipe10_n78), 
        .ZN(DP_reg_pipe10_n86) );
  NAND2_X1 DP_reg_pipe10_U45 ( .A1(DP_pipe0_coeff_pipe00[21]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n77) );
  NAND2_X1 DP_reg_pipe10_U44 ( .A1(DP_pipe10[21]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n78) );
  NAND2_X1 DP_reg_pipe10_U43 ( .A1(DP_reg_pipe10_n74), .A2(DP_reg_pipe10_n75), 
        .ZN(DP_reg_pipe10_n87) );
  NAND2_X1 DP_reg_pipe10_U42 ( .A1(DP_pipe0_coeff_pipe00[20]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n74) );
  NAND2_X1 DP_reg_pipe10_U41 ( .A1(DP_pipe10[20]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n75) );
  NAND2_X1 DP_reg_pipe10_U40 ( .A1(DP_reg_pipe10_n47), .A2(DP_reg_pipe10_n48), 
        .ZN(DP_reg_pipe10_n88) );
  NAND2_X1 DP_reg_pipe10_U39 ( .A1(DP_pipe0_coeff_pipe00[19]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n47) );
  NAND2_X1 DP_reg_pipe10_U38 ( .A1(DP_pipe10[19]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n48) );
  NAND2_X1 DP_reg_pipe10_U37 ( .A1(DP_reg_pipe10_n44), .A2(DP_reg_pipe10_n45), 
        .ZN(DP_reg_pipe10_n89) );
  NAND2_X1 DP_reg_pipe10_U36 ( .A1(DP_pipe0_coeff_pipe00[18]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n44) );
  NAND2_X1 DP_reg_pipe10_U35 ( .A1(DP_pipe10[18]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n45) );
  NAND2_X1 DP_reg_pipe10_U34 ( .A1(DP_reg_pipe10_n41), .A2(DP_reg_pipe10_n42), 
        .ZN(DP_reg_pipe10_n90) );
  NAND2_X1 DP_reg_pipe10_U33 ( .A1(DP_pipe0_coeff_pipe00[17]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n41) );
  NAND2_X1 DP_reg_pipe10_U32 ( .A1(DP_pipe10[17]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n42) );
  NAND2_X1 DP_reg_pipe10_U31 ( .A1(DP_reg_pipe10_n38), .A2(DP_reg_pipe10_n39), 
        .ZN(DP_reg_pipe10_n91) );
  NAND2_X1 DP_reg_pipe10_U30 ( .A1(DP_pipe0_coeff_pipe00[16]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n38) );
  NAND2_X1 DP_reg_pipe10_U29 ( .A1(DP_pipe10[16]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n39) );
  NAND2_X1 DP_reg_pipe10_U28 ( .A1(DP_reg_pipe10_n35), .A2(DP_reg_pipe10_n36), 
        .ZN(DP_reg_pipe10_n92) );
  NAND2_X1 DP_reg_pipe10_U27 ( .A1(DP_pipe0_coeff_pipe00[15]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n35) );
  NAND2_X1 DP_reg_pipe10_U26 ( .A1(DP_pipe10[15]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n36) );
  NAND2_X1 DP_reg_pipe10_U25 ( .A1(DP_reg_pipe10_n32), .A2(DP_reg_pipe10_n33), 
        .ZN(DP_reg_pipe10_n93) );
  NAND2_X1 DP_reg_pipe10_U24 ( .A1(DP_pipe0_coeff_pipe00[14]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n32) );
  NAND2_X1 DP_reg_pipe10_U23 ( .A1(DP_pipe10[14]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n33) );
  NAND2_X1 DP_reg_pipe10_U22 ( .A1(DP_reg_pipe10_n29), .A2(DP_reg_pipe10_n30), 
        .ZN(DP_reg_pipe10_n94) );
  NAND2_X1 DP_reg_pipe10_U21 ( .A1(DP_pipe0_coeff_pipe00[13]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n29) );
  NAND2_X1 DP_reg_pipe10_U20 ( .A1(DP_pipe10[13]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n30) );
  NAND2_X1 DP_reg_pipe10_U19 ( .A1(DP_reg_pipe10_n27), .A2(DP_reg_pipe10_n26), 
        .ZN(DP_reg_pipe10_n95) );
  NAND2_X1 DP_reg_pipe10_U18 ( .A1(DP_pipe10[12]), .A2(DP_reg_pipe10_n79), 
        .ZN(DP_reg_pipe10_n26) );
  INV_X1 DP_reg_pipe10_U17 ( .A(1'b1), .ZN(DP_reg_pipe10_n79) );
  NAND2_X1 DP_reg_pipe10_U16 ( .A1(DP_pipe0_coeff_pipe00[12]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n27) );
  MUX2_X1 DP_reg_pipe10_U15 ( .A(DP_pipe10[11]), .B(DP_pipe0_coeff_pipe00[11]), 
        .S(1'b1), .Z(DP_reg_pipe10_n96) );
  MUX2_X1 DP_reg_pipe10_U14 ( .A(DP_pipe10[10]), .B(DP_pipe0_coeff_pipe00[10]), 
        .S(1'b1), .Z(DP_reg_pipe10_n97) );
  MUX2_X1 DP_reg_pipe10_U13 ( .A(DP_pipe10[9]), .B(DP_pipe0_coeff_pipe00[9]), 
        .S(1'b1), .Z(DP_reg_pipe10_n98) );
  MUX2_X1 DP_reg_pipe10_U12 ( .A(DP_pipe10[8]), .B(DP_pipe0_coeff_pipe00[8]), 
        .S(1'b1), .Z(DP_reg_pipe10_n99) );
  MUX2_X1 DP_reg_pipe10_U11 ( .A(DP_pipe10[7]), .B(DP_pipe0_coeff_pipe00[7]), 
        .S(1'b1), .Z(DP_reg_pipe10_n100) );
  MUX2_X1 DP_reg_pipe10_U10 ( .A(DP_pipe10[6]), .B(DP_pipe0_coeff_pipe00[6]), 
        .S(1'b1), .Z(DP_reg_pipe10_n101) );
  MUX2_X1 DP_reg_pipe10_U9 ( .A(DP_pipe10[5]), .B(DP_pipe0_coeff_pipe00[5]), 
        .S(1'b1), .Z(DP_reg_pipe10_n102) );
  MUX2_X1 DP_reg_pipe10_U8 ( .A(DP_pipe10[4]), .B(DP_pipe0_coeff_pipe00[4]), 
        .S(1'b1), .Z(DP_reg_pipe10_n103) );
  MUX2_X1 DP_reg_pipe10_U7 ( .A(DP_pipe10[3]), .B(DP_pipe0_coeff_pipe00[3]), 
        .S(1'b1), .Z(DP_reg_pipe10_n104) );
  MUX2_X1 DP_reg_pipe10_U6 ( .A(DP_pipe10[2]), .B(DP_pipe0_coeff_pipe00[2]), 
        .S(1'b1), .Z(DP_reg_pipe10_n105) );
  MUX2_X1 DP_reg_pipe10_U5 ( .A(DP_pipe10[1]), .B(DP_pipe0_coeff_pipe00[1]), 
        .S(1'b1), .Z(DP_reg_pipe10_n106) );
  MUX2_X1 DP_reg_pipe10_U4 ( .A(DP_pipe10[0]), .B(DP_pipe0_coeff_pipe00[0]), 
        .S(1'b1), .Z(DP_reg_pipe10_n107) );
  BUF_X1 DP_reg_pipe10_U3 ( .A(DP_n6), .Z(DP_reg_pipe10_n12) );
  BUF_X1 DP_reg_pipe10_U2 ( .A(DP_n6), .Z(DP_reg_pipe10_n13) );
  DFFR_X1 DP_reg_pipe10_Q_reg_1_ ( .D(DP_reg_pipe10_n106), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[1]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_13_ ( .D(DP_reg_pipe10_n94), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[13]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_20_ ( .D(DP_reg_pipe10_n87), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[20]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_21_ ( .D(DP_reg_pipe10_n86), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[21]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_17_ ( .D(DP_reg_pipe10_n90), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[17]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_18_ ( .D(DP_reg_pipe10_n89), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[18]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_22_ ( .D(DP_reg_pipe10_n85), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[22]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_14_ ( .D(DP_reg_pipe10_n93), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[14]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_15_ ( .D(DP_reg_pipe10_n92), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[15]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_16_ ( .D(DP_reg_pipe10_n91), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[16]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_19_ ( .D(DP_reg_pipe10_n88), .CK(clk), .RN(DP_n6), .Q(DP_pipe10[19]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_0_ ( .D(DP_reg_pipe10_n107), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[0]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_2_ ( .D(DP_reg_pipe10_n105), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[2]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_3_ ( .D(DP_reg_pipe10_n104), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[3]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_4_ ( .D(DP_reg_pipe10_n103), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[4]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_5_ ( .D(DP_reg_pipe10_n102), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[5]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_6_ ( .D(DP_reg_pipe10_n101), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[6]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_7_ ( .D(DP_reg_pipe10_n100), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[7]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_8_ ( .D(DP_reg_pipe10_n99), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[8]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_9_ ( .D(DP_reg_pipe10_n98), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[9]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_10_ ( .D(DP_reg_pipe10_n97), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[10]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_11_ ( .D(DP_reg_pipe10_n96), .CK(clk), .RN(
        DP_reg_pipe10_n13), .Q(DP_pipe10[11]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_12_ ( .D(DP_reg_pipe10_n95), .CK(clk), .RN(
        DP_reg_pipe10_n12), .Q(DP_pipe10[12]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_23_ ( .D(DP_reg_pipe10_n84), .CK(clk), .RN(
        DP_reg_pipe10_n12), .Q(DP_pipe10[23]) );
  MUX2_X1 DP_reg_pipe11_U50 ( .A(DP_pipe11[23]), .B(DP_pipe0_coeff_pipe01[23]), 
        .S(1'b1), .Z(DP_reg_pipe11_n74) );
  NAND2_X1 DP_reg_pipe11_U49 ( .A1(DP_reg_pipe11_n48), .A2(DP_reg_pipe11_n73), 
        .ZN(DP_reg_pipe11_n75) );
  NAND2_X1 DP_reg_pipe11_U48 ( .A1(DP_pipe0_coeff_pipe01[22]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n48) );
  NAND2_X1 DP_reg_pipe11_U47 ( .A1(DP_pipe11[22]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n73) );
  NAND2_X1 DP_reg_pipe11_U46 ( .A1(DP_reg_pipe11_n45), .A2(DP_reg_pipe11_n46), 
        .ZN(DP_reg_pipe11_n76) );
  NAND2_X1 DP_reg_pipe11_U45 ( .A1(DP_pipe0_coeff_pipe01[21]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n45) );
  NAND2_X1 DP_reg_pipe11_U44 ( .A1(DP_pipe11[21]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n46) );
  NAND2_X1 DP_reg_pipe11_U43 ( .A1(DP_reg_pipe11_n43), .A2(DP_reg_pipe11_n44), 
        .ZN(DP_reg_pipe11_n77) );
  NAND2_X1 DP_reg_pipe11_U42 ( .A1(DP_pipe0_coeff_pipe01[20]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n43) );
  NAND2_X1 DP_reg_pipe11_U41 ( .A1(DP_pipe11[20]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n44) );
  NAND2_X1 DP_reg_pipe11_U40 ( .A1(DP_reg_pipe11_n41), .A2(DP_reg_pipe11_n42), 
        .ZN(DP_reg_pipe11_n78) );
  NAND2_X1 DP_reg_pipe11_U39 ( .A1(DP_pipe0_coeff_pipe01[19]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n41) );
  NAND2_X1 DP_reg_pipe11_U38 ( .A1(DP_pipe11[19]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n42) );
  NAND2_X1 DP_reg_pipe11_U37 ( .A1(DP_reg_pipe11_n39), .A2(DP_reg_pipe11_n40), 
        .ZN(DP_reg_pipe11_n79) );
  NAND2_X1 DP_reg_pipe11_U36 ( .A1(DP_pipe0_coeff_pipe01[18]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n39) );
  NAND2_X1 DP_reg_pipe11_U35 ( .A1(DP_pipe11[18]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n40) );
  NAND2_X1 DP_reg_pipe11_U34 ( .A1(DP_reg_pipe11_n37), .A2(DP_reg_pipe11_n38), 
        .ZN(DP_reg_pipe11_n80) );
  NAND2_X1 DP_reg_pipe11_U33 ( .A1(DP_pipe0_coeff_pipe01[17]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n37) );
  NAND2_X1 DP_reg_pipe11_U32 ( .A1(DP_pipe11[17]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n38) );
  NAND2_X1 DP_reg_pipe11_U31 ( .A1(DP_reg_pipe11_n35), .A2(DP_reg_pipe11_n36), 
        .ZN(DP_reg_pipe11_n81) );
  NAND2_X1 DP_reg_pipe11_U30 ( .A1(DP_pipe0_coeff_pipe01[16]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n35) );
  NAND2_X1 DP_reg_pipe11_U29 ( .A1(DP_pipe11[16]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n36) );
  NAND2_X1 DP_reg_pipe11_U28 ( .A1(DP_reg_pipe11_n33), .A2(DP_reg_pipe11_n34), 
        .ZN(DP_reg_pipe11_n82) );
  NAND2_X1 DP_reg_pipe11_U27 ( .A1(DP_pipe0_coeff_pipe01[15]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n33) );
  NAND2_X1 DP_reg_pipe11_U26 ( .A1(DP_pipe11[15]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n34) );
  NAND2_X1 DP_reg_pipe11_U25 ( .A1(DP_reg_pipe11_n31), .A2(DP_reg_pipe11_n32), 
        .ZN(DP_reg_pipe11_n83) );
  NAND2_X1 DP_reg_pipe11_U24 ( .A1(DP_pipe0_coeff_pipe01[14]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n31) );
  NAND2_X1 DP_reg_pipe11_U23 ( .A1(DP_pipe11[14]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n32) );
  NAND2_X1 DP_reg_pipe11_U22 ( .A1(DP_reg_pipe11_n29), .A2(DP_reg_pipe11_n30), 
        .ZN(DP_reg_pipe11_n84) );
  NAND2_X1 DP_reg_pipe11_U21 ( .A1(DP_pipe0_coeff_pipe01[13]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n29) );
  NAND2_X1 DP_reg_pipe11_U20 ( .A1(DP_pipe11[13]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n30) );
  NAND2_X1 DP_reg_pipe11_U19 ( .A1(DP_reg_pipe11_n28), .A2(DP_reg_pipe11_n27), 
        .ZN(DP_reg_pipe11_n85) );
  NAND2_X1 DP_reg_pipe11_U18 ( .A1(DP_pipe11[12]), .A2(DP_reg_pipe11_n47), 
        .ZN(DP_reg_pipe11_n27) );
  INV_X1 DP_reg_pipe11_U17 ( .A(1'b1), .ZN(DP_reg_pipe11_n47) );
  NAND2_X1 DP_reg_pipe11_U16 ( .A1(DP_pipe0_coeff_pipe01[12]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n28) );
  MUX2_X1 DP_reg_pipe11_U15 ( .A(DP_pipe11[4]), .B(DP_pipe0_coeff_pipe01[4]), 
        .S(1'b1), .Z(DP_reg_pipe11_n93) );
  MUX2_X1 DP_reg_pipe11_U14 ( .A(DP_pipe11[3]), .B(DP_pipe0_coeff_pipe01[3]), 
        .S(1'b1), .Z(DP_reg_pipe11_n94) );
  MUX2_X1 DP_reg_pipe11_U13 ( .A(DP_pipe11[2]), .B(DP_pipe0_coeff_pipe01[2]), 
        .S(1'b1), .Z(DP_reg_pipe11_n95) );
  MUX2_X1 DP_reg_pipe11_U12 ( .A(DP_pipe11[1]), .B(DP_pipe0_coeff_pipe01[1]), 
        .S(1'b1), .Z(DP_reg_pipe11_n96) );
  BUF_X1 DP_reg_pipe11_U11 ( .A(DP_n5), .Z(DP_reg_pipe11_n26) );
  MUX2_X1 DP_reg_pipe11_U10 ( .A(DP_pipe0_coeff_pipe01[11]), .B(DP_pipe11[11]), 
        .S(DP_reg_pipe11_n3), .Z(DP_reg_pipe11_n86) );
  MUX2_X1 DP_reg_pipe11_U9 ( .A(DP_pipe0_coeff_pipe01[10]), .B(DP_pipe11[10]), 
        .S(DP_reg_pipe11_n3), .Z(DP_reg_pipe11_n87) );
  MUX2_X1 DP_reg_pipe11_U8 ( .A(DP_pipe0_coeff_pipe01[9]), .B(DP_pipe11[9]), 
        .S(DP_reg_pipe11_n47), .Z(DP_reg_pipe11_n88) );
  MUX2_X1 DP_reg_pipe11_U7 ( .A(DP_pipe0_coeff_pipe01[8]), .B(DP_pipe11[8]), 
        .S(DP_reg_pipe11_n47), .Z(DP_reg_pipe11_n89) );
  MUX2_X1 DP_reg_pipe11_U6 ( .A(DP_pipe0_coeff_pipe01[7]), .B(DP_pipe11[7]), 
        .S(DP_reg_pipe11_n47), .Z(DP_reg_pipe11_n90) );
  MUX2_X1 DP_reg_pipe11_U5 ( .A(DP_pipe0_coeff_pipe01[6]), .B(DP_pipe11[6]), 
        .S(DP_reg_pipe11_n47), .Z(DP_reg_pipe11_n91) );
  MUX2_X1 DP_reg_pipe11_U4 ( .A(DP_pipe0_coeff_pipe01[5]), .B(DP_pipe11[5]), 
        .S(DP_reg_pipe11_n47), .Z(DP_reg_pipe11_n92) );
  MUX2_X1 DP_reg_pipe11_U3 ( .A(DP_pipe0_coeff_pipe01[0]), .B(DP_pipe11[0]), 
        .S(DP_reg_pipe11_n3), .Z(DP_reg_pipe11_n97) );
  INV_X1 DP_reg_pipe11_U2 ( .A(1'b1), .ZN(DP_reg_pipe11_n3) );
  DFFR_X1 DP_reg_pipe11_Q_reg_22_ ( .D(DP_reg_pipe11_n75), .CK(clk), .RN(
        DP_reg_pipe11_n26), .Q(DP_pipe11[22]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_17_ ( .D(DP_reg_pipe11_n80), .CK(clk), .RN(
        DP_reg_pipe11_n26), .Q(DP_pipe11[17]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_4_ ( .D(DP_reg_pipe11_n93), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[4]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_5_ ( .D(DP_reg_pipe11_n92), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[5]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_6_ ( .D(DP_reg_pipe11_n91), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[6]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_7_ ( .D(DP_reg_pipe11_n90), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[7]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_8_ ( .D(DP_reg_pipe11_n89), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[8]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_9_ ( .D(DP_reg_pipe11_n88), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[9]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_10_ ( .D(DP_reg_pipe11_n87), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[10]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_11_ ( .D(DP_reg_pipe11_n86), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[11]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_14_ ( .D(DP_reg_pipe11_n83), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[14]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_18_ ( .D(DP_reg_pipe11_n79), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[18]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_19_ ( .D(DP_reg_pipe11_n78), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[19]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_13_ ( .D(DP_reg_pipe11_n84), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[13]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_15_ ( .D(DP_reg_pipe11_n82), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[15]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_20_ ( .D(DP_reg_pipe11_n77), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[20]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_21_ ( .D(DP_reg_pipe11_n76), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[21]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_12_ ( .D(DP_reg_pipe11_n85), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[12]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_23_ ( .D(DP_reg_pipe11_n74), .CK(clk), .RN(DP_n5), .Q(DP_pipe11[23]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_3_ ( .D(DP_reg_pipe11_n94), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[3]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_0_ ( .D(DP_reg_pipe11_n97), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[0]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_2_ ( .D(DP_reg_pipe11_n95), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[2]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_1_ ( .D(DP_reg_pipe11_n96), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe11[1]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_16_ ( .D(DP_reg_pipe11_n81), .CK(clk), .RN(
        DP_reg_pipe11_n26), .Q(DP_pipe11[16]) );
  MUX2_X1 DP_reg_pipe12_U50 ( .A(DP_pipe12[23]), .B(DP_pipe0_coeff_pipe02[23]), 
        .S(1'b1), .Z(DP_reg_pipe12_n78) );
  NAND2_X1 DP_reg_pipe12_U49 ( .A1(DP_reg_pipe12_n75), .A2(DP_reg_pipe12_n76), 
        .ZN(DP_reg_pipe12_n79) );
  NAND2_X1 DP_reg_pipe12_U48 ( .A1(DP_pipe0_coeff_pipe02[22]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n75) );
  NAND2_X1 DP_reg_pipe12_U47 ( .A1(DP_pipe12[22]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n76) );
  NAND2_X1 DP_reg_pipe12_U46 ( .A1(DP_reg_pipe12_n47), .A2(DP_reg_pipe12_n48), 
        .ZN(DP_reg_pipe12_n80) );
  NAND2_X1 DP_reg_pipe12_U45 ( .A1(DP_pipe0_coeff_pipe02[21]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n47) );
  NAND2_X1 DP_reg_pipe12_U44 ( .A1(DP_pipe12[21]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n48) );
  NAND2_X1 DP_reg_pipe12_U43 ( .A1(DP_reg_pipe12_n44), .A2(DP_reg_pipe12_n45), 
        .ZN(DP_reg_pipe12_n81) );
  NAND2_X1 DP_reg_pipe12_U42 ( .A1(DP_pipe0_coeff_pipe02[20]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n44) );
  NAND2_X1 DP_reg_pipe12_U41 ( .A1(DP_pipe12[20]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n45) );
  NAND2_X1 DP_reg_pipe12_U40 ( .A1(DP_reg_pipe12_n41), .A2(DP_reg_pipe12_n42), 
        .ZN(DP_reg_pipe12_n82) );
  NAND2_X1 DP_reg_pipe12_U39 ( .A1(DP_pipe0_coeff_pipe02[19]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n41) );
  NAND2_X1 DP_reg_pipe12_U38 ( .A1(DP_pipe12[19]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n42) );
  NAND2_X1 DP_reg_pipe12_U37 ( .A1(DP_reg_pipe12_n38), .A2(DP_reg_pipe12_n39), 
        .ZN(DP_reg_pipe12_n83) );
  NAND2_X1 DP_reg_pipe12_U36 ( .A1(DP_pipe0_coeff_pipe02[18]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n38) );
  NAND2_X1 DP_reg_pipe12_U35 ( .A1(DP_pipe12[18]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n39) );
  NAND2_X1 DP_reg_pipe12_U34 ( .A1(DP_reg_pipe12_n35), .A2(DP_reg_pipe12_n36), 
        .ZN(DP_reg_pipe12_n84) );
  NAND2_X1 DP_reg_pipe12_U33 ( .A1(DP_pipe0_coeff_pipe02[17]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n35) );
  NAND2_X1 DP_reg_pipe12_U32 ( .A1(DP_pipe12[17]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n36) );
  NAND2_X1 DP_reg_pipe12_U31 ( .A1(DP_reg_pipe12_n32), .A2(DP_reg_pipe12_n33), 
        .ZN(DP_reg_pipe12_n85) );
  NAND2_X1 DP_reg_pipe12_U30 ( .A1(DP_pipe0_coeff_pipe02[16]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n32) );
  NAND2_X1 DP_reg_pipe12_U29 ( .A1(DP_pipe12[16]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n33) );
  NAND2_X1 DP_reg_pipe12_U28 ( .A1(DP_reg_pipe12_n29), .A2(DP_reg_pipe12_n30), 
        .ZN(DP_reg_pipe12_n86) );
  NAND2_X1 DP_reg_pipe12_U27 ( .A1(DP_pipe0_coeff_pipe02[15]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n29) );
  NAND2_X1 DP_reg_pipe12_U26 ( .A1(DP_pipe12[15]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n30) );
  NAND2_X1 DP_reg_pipe12_U25 ( .A1(DP_reg_pipe12_n26), .A2(DP_reg_pipe12_n27), 
        .ZN(DP_reg_pipe12_n87) );
  NAND2_X1 DP_reg_pipe12_U24 ( .A1(DP_pipe0_coeff_pipe02[14]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n26) );
  NAND2_X1 DP_reg_pipe12_U23 ( .A1(DP_pipe12[14]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n27) );
  NAND2_X1 DP_reg_pipe12_U22 ( .A1(DP_reg_pipe12_n23), .A2(DP_reg_pipe12_n24), 
        .ZN(DP_reg_pipe12_n88) );
  NAND2_X1 DP_reg_pipe12_U21 ( .A1(DP_pipe0_coeff_pipe02[13]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n23) );
  NAND2_X1 DP_reg_pipe12_U20 ( .A1(DP_pipe12[13]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n24) );
  NAND2_X1 DP_reg_pipe12_U19 ( .A1(DP_reg_pipe12_n21), .A2(DP_reg_pipe12_n20), 
        .ZN(DP_reg_pipe12_n89) );
  NAND2_X1 DP_reg_pipe12_U18 ( .A1(DP_pipe12[12]), .A2(DP_reg_pipe12_n73), 
        .ZN(DP_reg_pipe12_n20) );
  INV_X1 DP_reg_pipe12_U17 ( .A(1'b1), .ZN(DP_reg_pipe12_n73) );
  NAND2_X1 DP_reg_pipe12_U16 ( .A1(DP_pipe0_coeff_pipe02[12]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n21) );
  MUX2_X1 DP_reg_pipe12_U15 ( .A(DP_pipe12[11]), .B(DP_pipe0_coeff_pipe02[11]), 
        .S(1'b1), .Z(DP_reg_pipe12_n90) );
  MUX2_X1 DP_reg_pipe12_U14 ( .A(DP_pipe12[10]), .B(DP_pipe0_coeff_pipe02[10]), 
        .S(1'b1), .Z(DP_reg_pipe12_n91) );
  MUX2_X1 DP_reg_pipe12_U13 ( .A(DP_pipe12[9]), .B(DP_pipe0_coeff_pipe02[9]), 
        .S(1'b1), .Z(DP_reg_pipe12_n92) );
  MUX2_X1 DP_reg_pipe12_U12 ( .A(DP_pipe12[8]), .B(DP_pipe0_coeff_pipe02[8]), 
        .S(1'b1), .Z(DP_reg_pipe12_n93) );
  MUX2_X1 DP_reg_pipe12_U11 ( .A(DP_pipe12[7]), .B(DP_pipe0_coeff_pipe02[7]), 
        .S(1'b1), .Z(DP_reg_pipe12_n94) );
  MUX2_X1 DP_reg_pipe12_U10 ( .A(DP_pipe12[6]), .B(DP_pipe0_coeff_pipe02[6]), 
        .S(1'b1), .Z(DP_reg_pipe12_n95) );
  MUX2_X1 DP_reg_pipe12_U9 ( .A(DP_pipe12[5]), .B(DP_pipe0_coeff_pipe02[5]), 
        .S(1'b1), .Z(DP_reg_pipe12_n96) );
  MUX2_X1 DP_reg_pipe12_U8 ( .A(DP_pipe12[4]), .B(DP_pipe0_coeff_pipe02[4]), 
        .S(1'b1), .Z(DP_reg_pipe12_n97) );
  MUX2_X1 DP_reg_pipe12_U7 ( .A(DP_pipe12[3]), .B(DP_pipe0_coeff_pipe02[3]), 
        .S(1'b1), .Z(DP_reg_pipe12_n98) );
  MUX2_X1 DP_reg_pipe12_U6 ( .A(DP_pipe12[2]), .B(DP_pipe0_coeff_pipe02[2]), 
        .S(1'b1), .Z(DP_reg_pipe12_n99) );
  MUX2_X1 DP_reg_pipe12_U5 ( .A(DP_pipe12[1]), .B(DP_pipe0_coeff_pipe02[1]), 
        .S(1'b1), .Z(DP_reg_pipe12_n100) );
  BUF_X1 DP_reg_pipe12_U4 ( .A(DP_n5), .Z(DP_reg_pipe12_n7) );
  BUF_X1 DP_reg_pipe12_U3 ( .A(DP_n5), .Z(DP_reg_pipe12_n8) );
  MUX2_X1 DP_reg_pipe12_U2 ( .A(DP_pipe0_coeff_pipe02[0]), .B(DP_pipe12[0]), 
        .S(DP_reg_pipe12_n73), .Z(DP_reg_pipe12_n101) );
  DFFR_X1 DP_reg_pipe12_Q_reg_9_ ( .D(DP_reg_pipe12_n92), .CK(clk), .RN(DP_n5), 
        .Q(DP_pipe12[9]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_1_ ( .D(DP_reg_pipe12_n100), .CK(clk), .RN(DP_n5), .Q(DP_pipe12[1]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_16_ ( .D(DP_reg_pipe12_n85), .CK(clk), .RN(DP_n5), .Q(DP_pipe12[16]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_20_ ( .D(DP_reg_pipe12_n81), .CK(clk), .RN(DP_n5), .Q(DP_pipe12[20]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_21_ ( .D(DP_reg_pipe12_n80), .CK(clk), .RN(DP_n5), .Q(DP_pipe12[21]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_3_ ( .D(DP_reg_pipe12_n98), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[3]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_0_ ( .D(DP_reg_pipe12_n101), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[0]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_2_ ( .D(DP_reg_pipe12_n99), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[2]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_4_ ( .D(DP_reg_pipe12_n97), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[4]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_5_ ( .D(DP_reg_pipe12_n96), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[5]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_6_ ( .D(DP_reg_pipe12_n95), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[6]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_7_ ( .D(DP_reg_pipe12_n94), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[7]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_8_ ( .D(DP_reg_pipe12_n93), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[8]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_10_ ( .D(DP_reg_pipe12_n91), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[10]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_11_ ( .D(DP_reg_pipe12_n90), .CK(clk), .RN(
        DP_reg_pipe12_n8), .Q(DP_pipe12[11]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_12_ ( .D(DP_reg_pipe12_n89), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[12]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_13_ ( .D(DP_reg_pipe12_n88), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[13]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_14_ ( .D(DP_reg_pipe12_n87), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[14]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_15_ ( .D(DP_reg_pipe12_n86), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[15]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_17_ ( .D(DP_reg_pipe12_n84), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[17]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_18_ ( .D(DP_reg_pipe12_n83), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[18]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_19_ ( .D(DP_reg_pipe12_n82), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[19]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_22_ ( .D(DP_reg_pipe12_n79), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[22]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_23_ ( .D(DP_reg_pipe12_n78), .CK(clk), .RN(
        DP_reg_pipe12_n7), .Q(DP_pipe12[23]) );
  MUX2_X1 DP_reg_pipe13_U50 ( .A(DP_pipe13[23]), .B(DP_pipe0_coeff_pipe03[23]), 
        .S(1'b1), .Z(DP_reg_pipe13_n83) );
  NAND2_X1 DP_reg_pipe13_U49 ( .A1(DP_reg_pipe13_n80), .A2(DP_reg_pipe13_n81), 
        .ZN(DP_reg_pipe13_n84) );
  NAND2_X1 DP_reg_pipe13_U48 ( .A1(DP_pipe0_coeff_pipe03[22]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n80) );
  NAND2_X1 DP_reg_pipe13_U47 ( .A1(DP_pipe13[22]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n81) );
  NAND2_X1 DP_reg_pipe13_U46 ( .A1(DP_reg_pipe13_n76), .A2(DP_reg_pipe13_n77), 
        .ZN(DP_reg_pipe13_n85) );
  NAND2_X1 DP_reg_pipe13_U45 ( .A1(DP_pipe0_coeff_pipe03[21]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n76) );
  NAND2_X1 DP_reg_pipe13_U44 ( .A1(DP_pipe13[21]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n77) );
  NAND2_X1 DP_reg_pipe13_U43 ( .A1(DP_reg_pipe13_n73), .A2(DP_reg_pipe13_n74), 
        .ZN(DP_reg_pipe13_n86) );
  NAND2_X1 DP_reg_pipe13_U42 ( .A1(DP_pipe0_coeff_pipe03[20]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n73) );
  NAND2_X1 DP_reg_pipe13_U41 ( .A1(DP_pipe13[20]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n74) );
  NAND2_X1 DP_reg_pipe13_U40 ( .A1(DP_reg_pipe13_n47), .A2(DP_reg_pipe13_n46), 
        .ZN(DP_reg_pipe13_n87) );
  NAND2_X1 DP_reg_pipe13_U39 ( .A1(DP_pipe0_coeff_pipe03[19]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n46) );
  NAND2_X1 DP_reg_pipe13_U38 ( .A1(DP_pipe13[19]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n47) );
  NAND2_X1 DP_reg_pipe13_U37 ( .A1(DP_reg_pipe13_n43), .A2(DP_reg_pipe13_n44), 
        .ZN(DP_reg_pipe13_n88) );
  NAND2_X1 DP_reg_pipe13_U36 ( .A1(DP_pipe0_coeff_pipe03[18]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n43) );
  NAND2_X1 DP_reg_pipe13_U35 ( .A1(DP_pipe13[18]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n44) );
  NAND2_X1 DP_reg_pipe13_U34 ( .A1(DP_reg_pipe13_n40), .A2(DP_reg_pipe13_n41), 
        .ZN(DP_reg_pipe13_n89) );
  NAND2_X1 DP_reg_pipe13_U33 ( .A1(DP_pipe0_coeff_pipe03[17]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n40) );
  NAND2_X1 DP_reg_pipe13_U32 ( .A1(DP_pipe13[17]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n41) );
  NAND2_X1 DP_reg_pipe13_U31 ( .A1(DP_reg_pipe13_n37), .A2(DP_reg_pipe13_n38), 
        .ZN(DP_reg_pipe13_n90) );
  NAND2_X1 DP_reg_pipe13_U30 ( .A1(DP_pipe0_coeff_pipe03[16]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n37) );
  NAND2_X1 DP_reg_pipe13_U29 ( .A1(DP_pipe13[16]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n38) );
  NAND2_X1 DP_reg_pipe13_U28 ( .A1(DP_reg_pipe13_n34), .A2(DP_reg_pipe13_n35), 
        .ZN(DP_reg_pipe13_n91) );
  NAND2_X1 DP_reg_pipe13_U27 ( .A1(DP_pipe0_coeff_pipe03[15]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n34) );
  NAND2_X1 DP_reg_pipe13_U26 ( .A1(DP_pipe13[15]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n35) );
  NAND2_X1 DP_reg_pipe13_U25 ( .A1(DP_reg_pipe13_n31), .A2(DP_reg_pipe13_n32), 
        .ZN(DP_reg_pipe13_n92) );
  NAND2_X1 DP_reg_pipe13_U24 ( .A1(DP_pipe0_coeff_pipe03[14]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n31) );
  NAND2_X1 DP_reg_pipe13_U23 ( .A1(DP_pipe13[14]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n32) );
  NAND2_X1 DP_reg_pipe13_U22 ( .A1(DP_reg_pipe13_n28), .A2(DP_reg_pipe13_n29), 
        .ZN(DP_reg_pipe13_n93) );
  NAND2_X1 DP_reg_pipe13_U21 ( .A1(DP_pipe0_coeff_pipe03[13]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n28) );
  NAND2_X1 DP_reg_pipe13_U20 ( .A1(DP_pipe13[13]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n29) );
  NAND2_X1 DP_reg_pipe13_U19 ( .A1(DP_reg_pipe13_n26), .A2(DP_reg_pipe13_n25), 
        .ZN(DP_reg_pipe13_n94) );
  NAND2_X1 DP_reg_pipe13_U18 ( .A1(DP_pipe13[12]), .A2(DP_reg_pipe13_n78), 
        .ZN(DP_reg_pipe13_n25) );
  INV_X1 DP_reg_pipe13_U17 ( .A(1'b1), .ZN(DP_reg_pipe13_n78) );
  NAND2_X1 DP_reg_pipe13_U16 ( .A1(DP_pipe0_coeff_pipe03[12]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n26) );
  MUX2_X1 DP_reg_pipe13_U15 ( .A(DP_pipe13[11]), .B(DP_pipe0_coeff_pipe03[11]), 
        .S(1'b1), .Z(DP_reg_pipe13_n95) );
  MUX2_X1 DP_reg_pipe13_U14 ( .A(DP_pipe13[10]), .B(DP_pipe0_coeff_pipe03[10]), 
        .S(1'b1), .Z(DP_reg_pipe13_n96) );
  MUX2_X1 DP_reg_pipe13_U13 ( .A(DP_pipe13[9]), .B(DP_pipe0_coeff_pipe03[9]), 
        .S(1'b1), .Z(DP_reg_pipe13_n97) );
  MUX2_X1 DP_reg_pipe13_U12 ( .A(DP_pipe13[8]), .B(DP_pipe0_coeff_pipe03[8]), 
        .S(1'b1), .Z(DP_reg_pipe13_n98) );
  MUX2_X1 DP_reg_pipe13_U11 ( .A(DP_pipe13[7]), .B(DP_pipe0_coeff_pipe03[7]), 
        .S(1'b1), .Z(DP_reg_pipe13_n99) );
  MUX2_X1 DP_reg_pipe13_U10 ( .A(DP_pipe13[6]), .B(DP_pipe0_coeff_pipe03[6]), 
        .S(1'b1), .Z(DP_reg_pipe13_n100) );
  MUX2_X1 DP_reg_pipe13_U9 ( .A(DP_pipe13[5]), .B(DP_pipe0_coeff_pipe03[5]), 
        .S(1'b1), .Z(DP_reg_pipe13_n101) );
  MUX2_X1 DP_reg_pipe13_U8 ( .A(DP_pipe13[4]), .B(DP_pipe0_coeff_pipe03[4]), 
        .S(1'b1), .Z(DP_reg_pipe13_n102) );
  MUX2_X1 DP_reg_pipe13_U7 ( .A(DP_pipe13[3]), .B(DP_pipe0_coeff_pipe03[3]), 
        .S(1'b1), .Z(DP_reg_pipe13_n103) );
  MUX2_X1 DP_reg_pipe13_U6 ( .A(DP_pipe13[2]), .B(DP_pipe0_coeff_pipe03[2]), 
        .S(1'b1), .Z(DP_reg_pipe13_n104) );
  MUX2_X1 DP_reg_pipe13_U5 ( .A(DP_pipe13[1]), .B(DP_pipe0_coeff_pipe03[1]), 
        .S(1'b1), .Z(DP_reg_pipe13_n105) );
  BUF_X1 DP_reg_pipe13_U4 ( .A(DP_n4), .Z(DP_reg_pipe13_n13) );
  BUF_X1 DP_reg_pipe13_U3 ( .A(DP_n4), .Z(DP_reg_pipe13_n14) );
  MUX2_X1 DP_reg_pipe13_U2 ( .A(DP_pipe0_coeff_pipe03[0]), .B(DP_pipe13[0]), 
        .S(DP_reg_pipe13_n78), .Z(DP_reg_pipe13_n106) );
  DFFR_X1 DP_reg_pipe13_Q_reg_9_ ( .D(DP_reg_pipe13_n97), .CK(clk), .RN(DP_n4), 
        .Q(DP_pipe13[9]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_3_ ( .D(DP_reg_pipe13_n103), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[3]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_1_ ( .D(DP_reg_pipe13_n105), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[1]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_13_ ( .D(DP_reg_pipe13_n93), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[13]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_14_ ( .D(DP_reg_pipe13_n92), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[14]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_21_ ( .D(DP_reg_pipe13_n85), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[21]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_22_ ( .D(DP_reg_pipe13_n84), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[22]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_18_ ( .D(DP_reg_pipe13_n88), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[18]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_19_ ( .D(DP_reg_pipe13_n87), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[19]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_15_ ( .D(DP_reg_pipe13_n91), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[15]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_17_ ( .D(DP_reg_pipe13_n89), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[17]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_20_ ( .D(DP_reg_pipe13_n86), .CK(clk), .RN(DP_n4), .Q(DP_pipe13[20]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_0_ ( .D(DP_reg_pipe13_n106), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[0]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_2_ ( .D(DP_reg_pipe13_n104), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[2]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_4_ ( .D(DP_reg_pipe13_n102), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[4]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_5_ ( .D(DP_reg_pipe13_n101), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[5]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_6_ ( .D(DP_reg_pipe13_n100), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[6]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_7_ ( .D(DP_reg_pipe13_n99), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[7]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_8_ ( .D(DP_reg_pipe13_n98), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[8]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_10_ ( .D(DP_reg_pipe13_n96), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[10]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_11_ ( .D(DP_reg_pipe13_n95), .CK(clk), .RN(
        DP_reg_pipe13_n14), .Q(DP_pipe13[11]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_12_ ( .D(DP_reg_pipe13_n94), .CK(clk), .RN(
        DP_reg_pipe13_n13), .Q(DP_pipe13[12]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_16_ ( .D(DP_reg_pipe13_n90), .CK(clk), .RN(
        DP_reg_pipe13_n13), .Q(DP_pipe13[16]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_23_ ( .D(DP_reg_pipe13_n83), .CK(clk), .RN(
        DP_reg_pipe13_n13), .Q(DP_pipe13[23]) );
  MUX2_X1 DP_reg_out_U14 ( .A(dOut[11]), .B(DP_y_23), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n14) );
  MUX2_X1 DP_reg_out_U13 ( .A(dOut[10]), .B(DP_y_out[10]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n15) );
  MUX2_X1 DP_reg_out_U12 ( .A(dOut[9]), .B(DP_y_out[9]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n16) );
  MUX2_X1 DP_reg_out_U11 ( .A(dOut[8]), .B(DP_y_out[8]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n17) );
  MUX2_X1 DP_reg_out_U10 ( .A(dOut[7]), .B(DP_y_out[7]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n18) );
  MUX2_X1 DP_reg_out_U9 ( .A(dOut[6]), .B(DP_y_out[6]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n19) );
  MUX2_X1 DP_reg_out_U8 ( .A(dOut[5]), .B(DP_y_out[5]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n20) );
  MUX2_X1 DP_reg_out_U7 ( .A(dOut[4]), .B(DP_y_out[4]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n21) );
  MUX2_X1 DP_reg_out_U6 ( .A(dOut[3]), .B(DP_y_out[3]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n22) );
  MUX2_X1 DP_reg_out_U5 ( .A(dOut[2]), .B(DP_y_out[2]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n23) );
  MUX2_X1 DP_reg_out_U4 ( .A(dOut[1]), .B(DP_y_out[1]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n24) );
  MUX2_X1 DP_reg_out_U3 ( .A(dOut[0]), .B(DP_y_out[0]), .S(
        delayed_controls_2__0_), .Z(DP_reg_out_n26) );
  BUF_X1 DP_reg_out_U2 ( .A(DP_n4), .Z(DP_reg_out_n1) );
  DFFR_X1 DP_reg_out_Q_reg_0_ ( .D(DP_reg_out_n26), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[0]) );
  DFFR_X1 DP_reg_out_Q_reg_1_ ( .D(DP_reg_out_n24), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[1]) );
  DFFR_X1 DP_reg_out_Q_reg_2_ ( .D(DP_reg_out_n23), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[2]) );
  DFFR_X1 DP_reg_out_Q_reg_3_ ( .D(DP_reg_out_n22), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[3]) );
  DFFR_X1 DP_reg_out_Q_reg_4_ ( .D(DP_reg_out_n21), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[4]) );
  DFFR_X1 DP_reg_out_Q_reg_5_ ( .D(DP_reg_out_n20), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[5]) );
  DFFR_X1 DP_reg_out_Q_reg_6_ ( .D(DP_reg_out_n19), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[6]) );
  DFFR_X1 DP_reg_out_Q_reg_7_ ( .D(DP_reg_out_n18), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[7]) );
  DFFR_X1 DP_reg_out_Q_reg_8_ ( .D(DP_reg_out_n17), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[8]) );
  DFFR_X1 DP_reg_out_Q_reg_9_ ( .D(DP_reg_out_n16), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[9]) );
  DFFR_X1 DP_reg_out_Q_reg_10_ ( .D(DP_reg_out_n15), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[10]) );
  DFFR_X1 DP_reg_out_Q_reg_11_ ( .D(DP_reg_out_n14), .CK(clk), .RN(
        DP_reg_out_n1), .Q(dOut[11]) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U467 ( .A1(DP_pipe11[21]), .A2(
        DP_pipe13[21]), .ZN(DP_add_2_root_add_0_root_add_223_n47) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U466 ( .A1(DP_pipe11[19]), .A2(
        DP_pipe13[19]), .ZN(DP_add_2_root_add_0_root_add_223_n65) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U465 ( .A1(DP_pipe11[17]), .A2(
        DP_pipe13[17]), .ZN(DP_add_2_root_add_0_root_add_223_n83) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U464 ( .A1(DP_pipe11[7]), .A2(
        DP_pipe13[7]), .ZN(DP_add_2_root_add_0_root_add_223_n162) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U463 ( .A1(DP_pipe11[15]), .A2(
        DP_pipe13[15]), .ZN(DP_add_2_root_add_0_root_add_223_n95) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U462 ( .A1(DP_pipe11[3]), .A2(
        DP_pipe13[3]), .ZN(DP_add_2_root_add_0_root_add_223_n181) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U461 ( .A1(DP_pipe11[5]), .A2(
        DP_pipe13[5]), .ZN(DP_add_2_root_add_0_root_add_223_n170) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U460 ( .A1(DP_pipe11[13]), .A2(
        DP_pipe13[13]), .ZN(DP_add_2_root_add_0_root_add_223_n115) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U459 ( .A1(DP_pipe11[9]), .A2(
        DP_pipe13[9]), .ZN(DP_add_2_root_add_0_root_add_223_n151) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U458 ( .A1(DP_pipe11[1]), .A2(
        DP_pipe13[1]), .ZN(DP_add_2_root_add_0_root_add_223_n188) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U457 ( .A1(DP_pipe11[11]), .A2(
        DP_pipe13[11]), .ZN(DP_add_2_root_add_0_root_add_223_n133) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U456 ( .A1(DP_pipe11[22]), .A2(
        DP_pipe13[22]), .ZN(DP_add_2_root_add_0_root_add_223_n38) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U455 ( .A1(DP_pipe11[0]), .A2(
        DP_pipe13[0]), .ZN(DP_add_2_root_add_0_root_add_223_n190) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U454 ( .A1(DP_pipe11[6]), .A2(
        DP_pipe13[6]), .ZN(DP_add_2_root_add_0_root_add_223_n165) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U453 ( .A1(DP_pipe11[2]), .A2(
        DP_pipe13[2]), .ZN(DP_add_2_root_add_0_root_add_223_n184) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U452 ( .A1(DP_pipe11[8]), .A2(
        DP_pipe13[8]), .ZN(DP_add_2_root_add_0_root_add_223_n154) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U451 ( .A1(DP_pipe11[4]), .A2(
        DP_pipe13[4]), .ZN(DP_add_2_root_add_0_root_add_223_n175) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U450 ( .A1(DP_pipe11[10]), .A2(
        DP_pipe13[10]), .ZN(DP_add_2_root_add_0_root_add_223_n140) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U449 ( .A1(DP_pipe11[16]), .A2(
        DP_pipe13[16]), .ZN(DP_add_2_root_add_0_root_add_223_n86) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U448 ( .A1(DP_pipe11[14]), .A2(
        DP_pipe13[14]), .ZN(DP_add_2_root_add_0_root_add_223_n104) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U447 ( .A1(DP_pipe11[20]), .A2(
        DP_pipe13[20]), .ZN(DP_add_2_root_add_0_root_add_223_n54) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U446 ( .A1(DP_pipe11[18]), .A2(
        DP_pipe13[18]), .ZN(DP_add_2_root_add_0_root_add_223_n72) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U445 ( .A1(DP_pipe11[12]), .A2(
        DP_pipe13[12]), .ZN(DP_add_2_root_add_0_root_add_223_n122) );
  OR2_X1 DP_add_2_root_add_0_root_add_223_U444 ( .A1(DP_pipe11[23]), .A2(
        DP_pipe13[23]), .ZN(DP_add_2_root_add_0_root_add_223_n296) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U443 ( .A1(DP_pipe11[23]), .A2(
        DP_pipe13[23]), .ZN(DP_add_2_root_add_0_root_add_223_n27) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U442 ( .B1(
        DP_add_2_root_add_0_root_add_223_n1), .B2(
        DP_add_2_root_add_0_root_add_223_n295), .A(
        DP_add_2_root_add_0_root_add_223_n30), .ZN(
        DP_add_2_root_add_0_root_add_223_n28) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U441 ( .A1(
        DP_add_2_root_add_0_root_add_223_n296), .A2(
        DP_add_2_root_add_0_root_add_223_n27), .ZN(
        DP_add_2_root_add_0_root_add_223_n2) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U440 ( .A(
        DP_add_2_root_add_0_root_add_223_n28), .B(
        DP_add_2_root_add_0_root_add_223_n2), .ZN(DP_ff_23_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U439 ( .A(
        DP_add_2_root_add_0_root_add_223_n38), .ZN(
        DP_add_2_root_add_0_root_add_223_n36) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U438 ( .B1(
        DP_add_2_root_add_0_root_add_223_n45), .B2(
        DP_add_2_root_add_0_root_add_223_n35), .A(
        DP_add_2_root_add_0_root_add_223_n36), .ZN(
        DP_add_2_root_add_0_root_add_223_n34) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U437 ( .B1(
        DP_add_2_root_add_0_root_add_223_n61), .B2(
        DP_add_2_root_add_0_root_add_223_n33), .A(
        DP_add_2_root_add_0_root_add_223_n34), .ZN(
        DP_add_2_root_add_0_root_add_223_n32) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U436 ( .A(
        DP_add_2_root_add_0_root_add_223_n32), .ZN(
        DP_add_2_root_add_0_root_add_223_n30) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U435 ( .A(
        DP_add_2_root_add_0_root_add_223_n175), .ZN(
        DP_add_2_root_add_0_root_add_223_n173) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U434 ( .A(
        DP_add_2_root_add_0_root_add_223_n180), .ZN(
        DP_add_2_root_add_0_root_add_223_n211) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U433 ( .A1(
        DP_add_2_root_add_0_root_add_223_n211), .A2(
        DP_add_2_root_add_0_root_add_223_n181), .ZN(
        DP_add_2_root_add_0_root_add_223_n22) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U432 ( .B1(
        DP_add_2_root_add_0_root_add_223_n185), .B2(
        DP_add_2_root_add_0_root_add_223_n183), .A(
        DP_add_2_root_add_0_root_add_223_n184), .ZN(
        DP_add_2_root_add_0_root_add_223_n182) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U431 ( .A(
        DP_add_2_root_add_0_root_add_223_n182), .B(
        DP_add_2_root_add_0_root_add_223_n22), .ZN(DP_ff_3_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U430 ( .A(
        DP_add_2_root_add_0_root_add_223_n183), .ZN(
        DP_add_2_root_add_0_root_add_223_n212) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U429 ( .A1(
        DP_add_2_root_add_0_root_add_223_n212), .A2(
        DP_add_2_root_add_0_root_add_223_n184), .ZN(
        DP_add_2_root_add_0_root_add_223_n23) );
  XOR2_X1 DP_add_2_root_add_0_root_add_223_U428 ( .A(
        DP_add_2_root_add_0_root_add_223_n185), .B(
        DP_add_2_root_add_0_root_add_223_n23), .Z(DP_ff_2_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U427 ( .A(
        DP_add_2_root_add_0_root_add_223_n103), .ZN(
        DP_add_2_root_add_0_root_add_223_n102) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U426 ( .A(
        DP_add_2_root_add_0_root_add_223_n102), .ZN(
        DP_add_2_root_add_0_root_add_223_n101) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U425 ( .A(
        DP_add_2_root_add_0_root_add_223_n174), .ZN(
        DP_add_2_root_add_0_root_add_223_n172) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U424 ( .A(
        DP_add_2_root_add_0_root_add_223_n37), .ZN(
        DP_add_2_root_add_0_root_add_223_n35) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U423 ( .A(
        DP_add_2_root_add_0_root_add_223_n139), .ZN(
        DP_add_2_root_add_0_root_add_223_n137) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U422 ( .A(
        DP_add_2_root_add_0_root_add_223_n71), .ZN(
        DP_add_2_root_add_0_root_add_223_n69) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U421 ( .A(
        DP_add_2_root_add_0_root_add_223_n53), .ZN(
        DP_add_2_root_add_0_root_add_223_n51) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U420 ( .A(
        DP_add_2_root_add_0_root_add_223_n121), .ZN(
        DP_add_2_root_add_0_root_add_223_n119) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U419 ( .A(
        DP_add_2_root_add_0_root_add_223_n114), .ZN(
        DP_add_2_root_add_0_root_add_223_n201) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U418 ( .B1(
        DP_add_2_root_add_0_root_add_223_n155), .B2(
        DP_add_2_root_add_0_root_add_223_n117), .A(
        DP_add_2_root_add_0_root_add_223_n118), .ZN(
        DP_add_2_root_add_0_root_add_223_n116) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U417 ( .A1(
        DP_add_2_root_add_0_root_add_223_n201), .A2(
        DP_add_2_root_add_0_root_add_223_n115), .ZN(
        DP_add_2_root_add_0_root_add_223_n12) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U416 ( .A(
        DP_add_2_root_add_0_root_add_223_n116), .B(
        DP_add_2_root_add_0_root_add_223_n12), .ZN(DP_ff_13_) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U415 ( .B1(
        DP_add_2_root_add_0_root_add_223_n161), .B2(
        DP_add_2_root_add_0_root_add_223_n165), .A(
        DP_add_2_root_add_0_root_add_223_n162), .ZN(
        DP_add_2_root_add_0_root_add_223_n160) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U414 ( .A(
        DP_add_2_root_add_0_root_add_223_n72), .ZN(
        DP_add_2_root_add_0_root_add_223_n70) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U413 ( .B1(
        DP_add_2_root_add_0_root_add_223_n77), .B2(
        DP_add_2_root_add_0_root_add_223_n69), .A(
        DP_add_2_root_add_0_root_add_223_n70), .ZN(
        DP_add_2_root_add_0_root_add_223_n68) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U412 ( .A(
        DP_add_2_root_add_0_root_add_223_n54), .ZN(
        DP_add_2_root_add_0_root_add_223_n52) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U411 ( .B1(
        DP_add_2_root_add_0_root_add_223_n59), .B2(
        DP_add_2_root_add_0_root_add_223_n51), .A(
        DP_add_2_root_add_0_root_add_223_n52), .ZN(
        DP_add_2_root_add_0_root_add_223_n50) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U410 ( .A(
        DP_add_2_root_add_0_root_add_223_n140), .ZN(
        DP_add_2_root_add_0_root_add_223_n138) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U409 ( .B1(
        DP_add_2_root_add_0_root_add_223_n145), .B2(
        DP_add_2_root_add_0_root_add_223_n137), .A(
        DP_add_2_root_add_0_root_add_223_n138), .ZN(
        DP_add_2_root_add_0_root_add_223_n136) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U408 ( .A(
        DP_add_2_root_add_0_root_add_223_n122), .ZN(
        DP_add_2_root_add_0_root_add_223_n120) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U407 ( .B1(
        DP_add_2_root_add_0_root_add_223_n127), .B2(
        DP_add_2_root_add_0_root_add_223_n119), .A(
        DP_add_2_root_add_0_root_add_223_n120), .ZN(
        DP_add_2_root_add_0_root_add_223_n118) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U406 ( .B1(
        DP_add_2_root_add_0_root_add_223_n111), .B2(
        DP_add_2_root_add_0_root_add_223_n101), .A(
        DP_add_2_root_add_0_root_add_223_n104), .ZN(
        DP_add_2_root_add_0_root_add_223_n100) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U405 ( .B1(
        DP_add_2_root_add_0_root_add_223_n99), .B2(
        DP_add_2_root_add_0_root_add_223_n127), .A(
        DP_add_2_root_add_0_root_add_223_n100), .ZN(
        DP_add_2_root_add_0_root_add_223_n98) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U404 ( .B1(
        DP_add_2_root_add_0_root_add_223_n94), .B2(
        DP_add_2_root_add_0_root_add_223_n104), .A(
        DP_add_2_root_add_0_root_add_223_n95), .ZN(
        DP_add_2_root_add_0_root_add_223_n93) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U403 ( .B1(
        DP_add_2_root_add_0_root_add_223_n92), .B2(
        DP_add_2_root_add_0_root_add_223_n113), .A(
        DP_add_2_root_add_0_root_add_223_n93), .ZN(
        DP_add_2_root_add_0_root_add_223_n91) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U402 ( .A1(
        DP_add_2_root_add_0_root_add_223_n153), .A2(
        DP_add_2_root_add_0_root_add_223_n150), .ZN(
        DP_add_2_root_add_0_root_add_223_n148) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U401 ( .A1(
        DP_add_2_root_add_0_root_add_223_n53), .A2(
        DP_add_2_root_add_0_root_add_223_n46), .ZN(
        DP_add_2_root_add_0_root_add_223_n44) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U400 ( .A1(
        DP_add_2_root_add_0_root_add_223_n121), .A2(
        DP_add_2_root_add_0_root_add_223_n114), .ZN(
        DP_add_2_root_add_0_root_add_223_n112) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U399 ( .A1(
        DP_add_2_root_add_0_root_add_223_n85), .A2(
        DP_add_2_root_add_0_root_add_223_n82), .ZN(
        DP_add_2_root_add_0_root_add_223_n80) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U398 ( .A1(
        DP_add_2_root_add_0_root_add_223_n139), .A2(
        DP_add_2_root_add_0_root_add_223_n132), .ZN(
        DP_add_2_root_add_0_root_add_223_n130) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U397 ( .A1(
        DP_add_2_root_add_0_root_add_223_n103), .A2(
        DP_add_2_root_add_0_root_add_223_n94), .ZN(
        DP_add_2_root_add_0_root_add_223_n92) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U396 ( .A1(
        DP_add_2_root_add_0_root_add_223_n71), .A2(
        DP_add_2_root_add_0_root_add_223_n64), .ZN(
        DP_add_2_root_add_0_root_add_223_n62) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U395 ( .A1(
        DP_add_2_root_add_0_root_add_223_n174), .A2(
        DP_add_2_root_add_0_root_add_223_n169), .ZN(
        DP_add_2_root_add_0_root_add_223_n167) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U394 ( .A1(
        DP_add_2_root_add_0_root_add_223_n164), .A2(
        DP_add_2_root_add_0_root_add_223_n161), .ZN(
        DP_add_2_root_add_0_root_add_223_n159) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U393 ( .B1(
        DP_add_2_root_add_0_root_add_223_n159), .B2(
        DP_add_2_root_add_0_root_add_223_n168), .A(
        DP_add_2_root_add_0_root_add_223_n160), .ZN(
        DP_add_2_root_add_0_root_add_223_n158) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U392 ( .A1(
        DP_add_2_root_add_0_root_add_223_n167), .A2(
        DP_add_2_root_add_0_root_add_223_n159), .ZN(
        DP_add_2_root_add_0_root_add_223_n157) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U391 ( .B1(
        DP_add_2_root_add_0_root_add_223_n177), .B2(
        DP_add_2_root_add_0_root_add_223_n157), .A(
        DP_add_2_root_add_0_root_add_223_n158), .ZN(
        DP_add_2_root_add_0_root_add_223_n156) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U390 ( .B1(
        DP_add_2_root_add_0_root_add_223_n46), .B2(
        DP_add_2_root_add_0_root_add_223_n54), .A(
        DP_add_2_root_add_0_root_add_223_n47), .ZN(
        DP_add_2_root_add_0_root_add_223_n45) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U389 ( .B1(
        DP_add_2_root_add_0_root_add_223_n169), .B2(
        DP_add_2_root_add_0_root_add_223_n175), .A(
        DP_add_2_root_add_0_root_add_223_n170), .ZN(
        DP_add_2_root_add_0_root_add_223_n168) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U388 ( .B1(
        DP_add_2_root_add_0_root_add_223_n187), .B2(
        DP_add_2_root_add_0_root_add_223_n190), .A(
        DP_add_2_root_add_0_root_add_223_n188), .ZN(
        DP_add_2_root_add_0_root_add_223_n186) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U387 ( .B1(
        DP_add_2_root_add_0_root_add_223_n150), .B2(
        DP_add_2_root_add_0_root_add_223_n154), .A(
        DP_add_2_root_add_0_root_add_223_n151), .ZN(
        DP_add_2_root_add_0_root_add_223_n149) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U386 ( .B1(
        DP_add_2_root_add_0_root_add_223_n82), .B2(
        DP_add_2_root_add_0_root_add_223_n86), .A(
        DP_add_2_root_add_0_root_add_223_n83), .ZN(
        DP_add_2_root_add_0_root_add_223_n81) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U385 ( .B1(
        DP_add_2_root_add_0_root_add_223_n114), .B2(
        DP_add_2_root_add_0_root_add_223_n122), .A(
        DP_add_2_root_add_0_root_add_223_n115), .ZN(
        DP_add_2_root_add_0_root_add_223_n113) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U384 ( .B1(
        DP_add_2_root_add_0_root_add_223_n180), .B2(
        DP_add_2_root_add_0_root_add_223_n184), .A(
        DP_add_2_root_add_0_root_add_223_n181), .ZN(
        DP_add_2_root_add_0_root_add_223_n179) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U383 ( .A1(
        DP_add_2_root_add_0_root_add_223_n183), .A2(
        DP_add_2_root_add_0_root_add_223_n180), .ZN(
        DP_add_2_root_add_0_root_add_223_n178) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U382 ( .B1(
        DP_add_2_root_add_0_root_add_223_n178), .B2(
        DP_add_2_root_add_0_root_add_223_n186), .A(
        DP_add_2_root_add_0_root_add_223_n179), .ZN(
        DP_add_2_root_add_0_root_add_223_n177) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U381 ( .B1(
        DP_add_2_root_add_0_root_add_223_n64), .B2(
        DP_add_2_root_add_0_root_add_223_n72), .A(
        DP_add_2_root_add_0_root_add_223_n65), .ZN(
        DP_add_2_root_add_0_root_add_223_n63) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U380 ( .B1(
        DP_add_2_root_add_0_root_add_223_n62), .B2(
        DP_add_2_root_add_0_root_add_223_n81), .A(
        DP_add_2_root_add_0_root_add_223_n63), .ZN(
        DP_add_2_root_add_0_root_add_223_n61) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U379 ( .B1(
        DP_add_2_root_add_0_root_add_223_n132), .B2(
        DP_add_2_root_add_0_root_add_223_n140), .A(
        DP_add_2_root_add_0_root_add_223_n133), .ZN(
        DP_add_2_root_add_0_root_add_223_n131) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U378 ( .B1(
        DP_add_2_root_add_0_root_add_223_n130), .B2(
        DP_add_2_root_add_0_root_add_223_n149), .A(
        DP_add_2_root_add_0_root_add_223_n131), .ZN(
        DP_add_2_root_add_0_root_add_223_n129) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U377 ( .A(
        DP_add_2_root_add_0_root_add_223_n82), .ZN(
        DP_add_2_root_add_0_root_add_223_n197) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U376 ( .B1(
        DP_add_2_root_add_0_root_add_223_n1), .B2(
        DP_add_2_root_add_0_root_add_223_n85), .A(
        DP_add_2_root_add_0_root_add_223_n86), .ZN(
        DP_add_2_root_add_0_root_add_223_n84) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U375 ( .A1(
        DP_add_2_root_add_0_root_add_223_n197), .A2(
        DP_add_2_root_add_0_root_add_223_n83), .ZN(
        DP_add_2_root_add_0_root_add_223_n8) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U374 ( .A(
        DP_add_2_root_add_0_root_add_223_n84), .B(
        DP_add_2_root_add_0_root_add_223_n8), .ZN(DP_ff_17_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U373 ( .A(
        DP_add_2_root_add_0_root_add_223_n64), .ZN(
        DP_add_2_root_add_0_root_add_223_n195) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U372 ( .B1(
        DP_add_2_root_add_0_root_add_223_n1), .B2(
        DP_add_2_root_add_0_root_add_223_n67), .A(
        DP_add_2_root_add_0_root_add_223_n68), .ZN(
        DP_add_2_root_add_0_root_add_223_n66) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U371 ( .A1(
        DP_add_2_root_add_0_root_add_223_n195), .A2(
        DP_add_2_root_add_0_root_add_223_n65), .ZN(
        DP_add_2_root_add_0_root_add_223_n6) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U370 ( .A(
        DP_add_2_root_add_0_root_add_223_n66), .B(
        DP_add_2_root_add_0_root_add_223_n6), .ZN(DP_ff_19_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U369 ( .A(
        DP_add_2_root_add_0_root_add_223_n46), .ZN(
        DP_add_2_root_add_0_root_add_223_n193) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U368 ( .B1(
        DP_add_2_root_add_0_root_add_223_n1), .B2(
        DP_add_2_root_add_0_root_add_223_n49), .A(
        DP_add_2_root_add_0_root_add_223_n50), .ZN(
        DP_add_2_root_add_0_root_add_223_n48) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U367 ( .A1(
        DP_add_2_root_add_0_root_add_223_n193), .A2(
        DP_add_2_root_add_0_root_add_223_n47), .ZN(
        DP_add_2_root_add_0_root_add_223_n4) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U366 ( .A(
        DP_add_2_root_add_0_root_add_223_n48), .B(
        DP_add_2_root_add_0_root_add_223_n4), .ZN(DP_ff_21_) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U365 ( .B1(
        DP_add_2_root_add_0_root_add_223_n1), .B2(
        DP_add_2_root_add_0_root_add_223_n74), .A(
        DP_add_2_root_add_0_root_add_223_n75), .ZN(
        DP_add_2_root_add_0_root_add_223_n73) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U364 ( .A1(
        DP_add_2_root_add_0_root_add_223_n69), .A2(
        DP_add_2_root_add_0_root_add_223_n72), .ZN(
        DP_add_2_root_add_0_root_add_223_n7) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U363 ( .A(
        DP_add_2_root_add_0_root_add_223_n73), .B(
        DP_add_2_root_add_0_root_add_223_n7), .ZN(DP_ff_18_) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U362 ( .B1(
        DP_add_2_root_add_0_root_add_223_n1), .B2(
        DP_add_2_root_add_0_root_add_223_n56), .A(
        DP_add_2_root_add_0_root_add_223_n57), .ZN(
        DP_add_2_root_add_0_root_add_223_n55) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U361 ( .A1(
        DP_add_2_root_add_0_root_add_223_n51), .A2(
        DP_add_2_root_add_0_root_add_223_n54), .ZN(
        DP_add_2_root_add_0_root_add_223_n5) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U360 ( .A(
        DP_add_2_root_add_0_root_add_223_n55), .B(
        DP_add_2_root_add_0_root_add_223_n5), .ZN(DP_ff_20_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U359 ( .A(
        DP_add_2_root_add_0_root_add_223_n37), .ZN(
        DP_add_2_root_add_0_root_add_223_n192) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U358 ( .B1(
        DP_add_2_root_add_0_root_add_223_n1), .B2(
        DP_add_2_root_add_0_root_add_223_n40), .A(
        DP_add_2_root_add_0_root_add_223_n41), .ZN(
        DP_add_2_root_add_0_root_add_223_n39) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U357 ( .A1(
        DP_add_2_root_add_0_root_add_223_n192), .A2(
        DP_add_2_root_add_0_root_add_223_n38), .ZN(
        DP_add_2_root_add_0_root_add_223_n3) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U356 ( .A(
        DP_add_2_root_add_0_root_add_223_n39), .B(
        DP_add_2_root_add_0_root_add_223_n3), .ZN(DP_ff_22_) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U355 ( .A1(
        DP_add_2_root_add_0_root_add_223_n172), .A2(
        DP_add_2_root_add_0_root_add_223_n175), .ZN(
        DP_add_2_root_add_0_root_add_223_n21) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U354 ( .A(
        DP_add_2_root_add_0_root_add_223_n176), .B(
        DP_add_2_root_add_0_root_add_223_n21), .ZN(DP_ff_4_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U353 ( .A(
        DP_add_2_root_add_0_root_add_223_n94), .ZN(
        DP_add_2_root_add_0_root_add_223_n199) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U352 ( .B1(
        DP_add_2_root_add_0_root_add_223_n155), .B2(
        DP_add_2_root_add_0_root_add_223_n97), .A(
        DP_add_2_root_add_0_root_add_223_n98), .ZN(
        DP_add_2_root_add_0_root_add_223_n96) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U351 ( .A1(
        DP_add_2_root_add_0_root_add_223_n199), .A2(
        DP_add_2_root_add_0_root_add_223_n95), .ZN(
        DP_add_2_root_add_0_root_add_223_n10) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U350 ( .A(
        DP_add_2_root_add_0_root_add_223_n96), .B(
        DP_add_2_root_add_0_root_add_223_n10), .ZN(DP_ff_15_) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U349 ( .B1(
        DP_add_2_root_add_0_root_add_223_n155), .B2(
        DP_add_2_root_add_0_root_add_223_n142), .A(
        DP_add_2_root_add_0_root_add_223_n143), .ZN(
        DP_add_2_root_add_0_root_add_223_n141) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U348 ( .A1(
        DP_add_2_root_add_0_root_add_223_n137), .A2(
        DP_add_2_root_add_0_root_add_223_n140), .ZN(
        DP_add_2_root_add_0_root_add_223_n15) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U347 ( .A(
        DP_add_2_root_add_0_root_add_223_n141), .B(
        DP_add_2_root_add_0_root_add_223_n15), .ZN(DP_ff_10_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U346 ( .A(
        DP_add_2_root_add_0_root_add_223_n132), .ZN(
        DP_add_2_root_add_0_root_add_223_n203) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U345 ( .B1(
        DP_add_2_root_add_0_root_add_223_n155), .B2(
        DP_add_2_root_add_0_root_add_223_n135), .A(
        DP_add_2_root_add_0_root_add_223_n136), .ZN(
        DP_add_2_root_add_0_root_add_223_n134) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U344 ( .A1(
        DP_add_2_root_add_0_root_add_223_n203), .A2(
        DP_add_2_root_add_0_root_add_223_n133), .ZN(
        DP_add_2_root_add_0_root_add_223_n14) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U343 ( .A(
        DP_add_2_root_add_0_root_add_223_n134), .B(
        DP_add_2_root_add_0_root_add_223_n14), .ZN(DP_ff_11_) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U342 ( .B1(
        DP_add_2_root_add_0_root_add_223_n155), .B2(
        DP_add_2_root_add_0_root_add_223_n124), .A(
        DP_add_2_root_add_0_root_add_223_n125), .ZN(
        DP_add_2_root_add_0_root_add_223_n123) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U341 ( .A1(
        DP_add_2_root_add_0_root_add_223_n119), .A2(
        DP_add_2_root_add_0_root_add_223_n122), .ZN(
        DP_add_2_root_add_0_root_add_223_n13) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U340 ( .A(
        DP_add_2_root_add_0_root_add_223_n123), .B(
        DP_add_2_root_add_0_root_add_223_n13), .ZN(DP_ff_12_) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U339 ( .B1(
        DP_add_2_root_add_0_root_add_223_n155), .B2(
        DP_add_2_root_add_0_root_add_223_n106), .A(
        DP_add_2_root_add_0_root_add_223_n107), .ZN(
        DP_add_2_root_add_0_root_add_223_n105) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U338 ( .A1(
        DP_add_2_root_add_0_root_add_223_n102), .A2(
        DP_add_2_root_add_0_root_add_223_n104), .ZN(
        DP_add_2_root_add_0_root_add_223_n11) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U337 ( .A(
        DP_add_2_root_add_0_root_add_223_n105), .B(
        DP_add_2_root_add_0_root_add_223_n11), .ZN(DP_ff_14_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U336 ( .A(
        DP_add_2_root_add_0_root_add_223_n161), .ZN(
        DP_add_2_root_add_0_root_add_223_n207) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U335 ( .B1(
        DP_add_2_root_add_0_root_add_223_n166), .B2(
        DP_add_2_root_add_0_root_add_223_n164), .A(
        DP_add_2_root_add_0_root_add_223_n165), .ZN(
        DP_add_2_root_add_0_root_add_223_n163) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U334 ( .A1(
        DP_add_2_root_add_0_root_add_223_n207), .A2(
        DP_add_2_root_add_0_root_add_223_n162), .ZN(
        DP_add_2_root_add_0_root_add_223_n18) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U333 ( .A(
        DP_add_2_root_add_0_root_add_223_n163), .B(
        DP_add_2_root_add_0_root_add_223_n18), .ZN(DP_ff_7_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U332 ( .A(
        DP_add_2_root_add_0_root_add_223_n150), .ZN(
        DP_add_2_root_add_0_root_add_223_n205) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U331 ( .B1(
        DP_add_2_root_add_0_root_add_223_n155), .B2(
        DP_add_2_root_add_0_root_add_223_n153), .A(
        DP_add_2_root_add_0_root_add_223_n154), .ZN(
        DP_add_2_root_add_0_root_add_223_n152) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U330 ( .A1(
        DP_add_2_root_add_0_root_add_223_n205), .A2(
        DP_add_2_root_add_0_root_add_223_n151), .ZN(
        DP_add_2_root_add_0_root_add_223_n16) );
  XNOR2_X1 DP_add_2_root_add_0_root_add_223_U329 ( .A(
        DP_add_2_root_add_0_root_add_223_n152), .B(
        DP_add_2_root_add_0_root_add_223_n16), .ZN(DP_ff_9_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U328 ( .A(
        DP_add_2_root_add_0_root_add_223_n187), .ZN(
        DP_add_2_root_add_0_root_add_223_n213) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U327 ( .A1(
        DP_add_2_root_add_0_root_add_223_n213), .A2(
        DP_add_2_root_add_0_root_add_223_n188), .ZN(
        DP_add_2_root_add_0_root_add_223_n24) );
  XOR2_X1 DP_add_2_root_add_0_root_add_223_U326 ( .A(
        DP_add_2_root_add_0_root_add_223_n24), .B(
        DP_add_2_root_add_0_root_add_223_n190), .Z(DP_ff_1_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U325 ( .A(
        DP_add_2_root_add_0_root_add_223_n169), .ZN(
        DP_add_2_root_add_0_root_add_223_n209) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U324 ( .B1(
        DP_add_2_root_add_0_root_add_223_n176), .B2(
        DP_add_2_root_add_0_root_add_223_n172), .A(
        DP_add_2_root_add_0_root_add_223_n173), .ZN(
        DP_add_2_root_add_0_root_add_223_n171) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U323 ( .A1(
        DP_add_2_root_add_0_root_add_223_n209), .A2(
        DP_add_2_root_add_0_root_add_223_n170), .ZN(
        DP_add_2_root_add_0_root_add_223_n20) );
  XOR2_X1 DP_add_2_root_add_0_root_add_223_U322 ( .A(
        DP_add_2_root_add_0_root_add_223_n171), .B(
        DP_add_2_root_add_0_root_add_223_n20), .Z(DP_ff_5_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U321 ( .A(
        DP_add_2_root_add_0_root_add_223_n164), .ZN(
        DP_add_2_root_add_0_root_add_223_n208) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U320 ( .A1(
        DP_add_2_root_add_0_root_add_223_n208), .A2(
        DP_add_2_root_add_0_root_add_223_n165), .ZN(
        DP_add_2_root_add_0_root_add_223_n19) );
  XOR2_X1 DP_add_2_root_add_0_root_add_223_U319 ( .A(
        DP_add_2_root_add_0_root_add_223_n166), .B(
        DP_add_2_root_add_0_root_add_223_n19), .Z(DP_ff_6_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U318 ( .A(
        DP_add_2_root_add_0_root_add_223_n153), .ZN(
        DP_add_2_root_add_0_root_add_223_n206) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U317 ( .A1(
        DP_add_2_root_add_0_root_add_223_n206), .A2(
        DP_add_2_root_add_0_root_add_223_n154), .ZN(
        DP_add_2_root_add_0_root_add_223_n17) );
  XOR2_X1 DP_add_2_root_add_0_root_add_223_U316 ( .A(
        DP_add_2_root_add_0_root_add_223_n155), .B(
        DP_add_2_root_add_0_root_add_223_n17), .Z(DP_ff_8_) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U315 ( .A(
        DP_add_2_root_add_0_root_add_223_n85), .ZN(
        DP_add_2_root_add_0_root_add_223_n198) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U314 ( .A1(
        DP_add_2_root_add_0_root_add_223_n198), .A2(
        DP_add_2_root_add_0_root_add_223_n86), .ZN(
        DP_add_2_root_add_0_root_add_223_n9) );
  XOR2_X1 DP_add_2_root_add_0_root_add_223_U313 ( .A(
        DP_add_2_root_add_0_root_add_223_n1), .B(
        DP_add_2_root_add_0_root_add_223_n9), .Z(DP_ff_16_) );
  OAI21_X1 DP_add_2_root_add_0_root_add_223_U312 ( .B1(
        DP_add_2_root_add_0_root_add_223_n129), .B2(
        DP_add_2_root_add_0_root_add_223_n90), .A(
        DP_add_2_root_add_0_root_add_223_n91), .ZN(
        DP_add_2_root_add_0_root_add_223_n89) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U311 ( .A1(
        DP_add_2_root_add_0_root_add_223_n128), .A2(
        DP_add_2_root_add_0_root_add_223_n90), .ZN(
        DP_add_2_root_add_0_root_add_223_n88) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U310 ( .B1(
        DP_add_2_root_add_0_root_add_223_n156), .B2(
        DP_add_2_root_add_0_root_add_223_n88), .A(
        DP_add_2_root_add_0_root_add_223_n89), .ZN(
        DP_add_2_root_add_0_root_add_223_n87) );
  BUF_X1 DP_add_2_root_add_0_root_add_223_U309 ( .A(
        DP_add_2_root_add_0_root_add_223_n87), .Z(
        DP_add_2_root_add_0_root_add_223_n1) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U308 ( .A1(
        DP_add_2_root_add_0_root_add_223_n76), .A2(
        DP_add_2_root_add_0_root_add_223_n69), .ZN(
        DP_add_2_root_add_0_root_add_223_n67) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U307 ( .A1(
        DP_add_2_root_add_0_root_add_223_n58), .A2(
        DP_add_2_root_add_0_root_add_223_n51), .ZN(
        DP_add_2_root_add_0_root_add_223_n49) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U306 ( .A1(
        DP_add_2_root_add_0_root_add_223_n148), .A2(
        DP_add_2_root_add_0_root_add_223_n137), .ZN(
        DP_add_2_root_add_0_root_add_223_n135) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U305 ( .A1(
        DP_add_2_root_add_0_root_add_223_n126), .A2(
        DP_add_2_root_add_0_root_add_223_n119), .ZN(
        DP_add_2_root_add_0_root_add_223_n117) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U304 ( .A(
        DP_add_2_root_add_0_root_add_223_n80), .ZN(
        DP_add_2_root_add_0_root_add_223_n78) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U303 ( .A(
        DP_add_2_root_add_0_root_add_223_n78), .ZN(
        DP_add_2_root_add_0_root_add_223_n76) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U302 ( .A(
        DP_add_2_root_add_0_root_add_223_n149), .ZN(
        DP_add_2_root_add_0_root_add_223_n147) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U301 ( .A(
        DP_add_2_root_add_0_root_add_223_n147), .ZN(
        DP_add_2_root_add_0_root_add_223_n145) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U300 ( .A(
        DP_add_2_root_add_0_root_add_223_n81), .ZN(
        DP_add_2_root_add_0_root_add_223_n79) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U299 ( .A(
        DP_add_2_root_add_0_root_add_223_n79), .ZN(
        DP_add_2_root_add_0_root_add_223_n77) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U298 ( .A(
        DP_add_2_root_add_0_root_add_223_n44), .ZN(
        DP_add_2_root_add_0_root_add_223_n43) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U297 ( .A(
        DP_add_2_root_add_0_root_add_223_n43), .ZN(
        DP_add_2_root_add_0_root_add_223_n42) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U296 ( .A(
        DP_add_2_root_add_0_root_add_223_n186), .ZN(
        DP_add_2_root_add_0_root_add_223_n185) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U295 ( .A(
        DP_add_2_root_add_0_root_add_223_n112), .ZN(
        DP_add_2_root_add_0_root_add_223_n110) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U294 ( .A(
        DP_add_2_root_add_0_root_add_223_n113), .ZN(
        DP_add_2_root_add_0_root_add_223_n111) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U293 ( .A(
        DP_add_2_root_add_0_root_add_223_n177), .ZN(
        DP_add_2_root_add_0_root_add_223_n176) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U292 ( .A1(
        DP_add_2_root_add_0_root_add_223_n44), .A2(
        DP_add_2_root_add_0_root_add_223_n35), .ZN(
        DP_add_2_root_add_0_root_add_223_n33) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U291 ( .A1(
        DP_add_2_root_add_0_root_add_223_n80), .A2(
        DP_add_2_root_add_0_root_add_223_n62), .ZN(
        DP_add_2_root_add_0_root_add_223_n60) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U290 ( .A1(
        DP_add_2_root_add_0_root_add_223_n148), .A2(
        DP_add_2_root_add_0_root_add_223_n130), .ZN(
        DP_add_2_root_add_0_root_add_223_n128) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U289 ( .A1(
        DP_add_2_root_add_0_root_add_223_n112), .A2(
        DP_add_2_root_add_0_root_add_223_n92), .ZN(
        DP_add_2_root_add_0_root_add_223_n90) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U288 ( .A(
        DP_add_2_root_add_0_root_add_223_n61), .ZN(
        DP_add_2_root_add_0_root_add_223_n59) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U287 ( .A(
        DP_add_2_root_add_0_root_add_223_n129), .ZN(
        DP_add_2_root_add_0_root_add_223_n127) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U286 ( .B1(
        DP_add_2_root_add_0_root_add_223_n59), .B2(
        DP_add_2_root_add_0_root_add_223_n42), .A(
        DP_add_2_root_add_0_root_add_223_n45), .ZN(
        DP_add_2_root_add_0_root_add_223_n41) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U285 ( .A1(
        DP_add_2_root_add_0_root_add_223_n110), .A2(
        DP_add_2_root_add_0_root_add_223_n101), .ZN(
        DP_add_2_root_add_0_root_add_223_n99) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U284 ( .B1(
        DP_add_2_root_add_0_root_add_223_n176), .B2(
        DP_add_2_root_add_0_root_add_223_n167), .A(
        DP_add_2_root_add_0_root_add_223_n168), .ZN(
        DP_add_2_root_add_0_root_add_223_n166) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U283 ( .A(
        DP_add_2_root_add_0_root_add_223_n77), .ZN(
        DP_add_2_root_add_0_root_add_223_n75) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U282 ( .A(
        DP_add_2_root_add_0_root_add_223_n145), .ZN(
        DP_add_2_root_add_0_root_add_223_n143) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U281 ( .A(
        DP_add_2_root_add_0_root_add_223_n76), .ZN(
        DP_add_2_root_add_0_root_add_223_n74) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U280 ( .A(
        DP_add_2_root_add_0_root_add_223_n148), .ZN(
        DP_add_2_root_add_0_root_add_223_n142) );
  OR2_X1 DP_add_2_root_add_0_root_add_223_U279 ( .A1(
        DP_add_2_root_add_0_root_add_223_n60), .A2(
        DP_add_2_root_add_0_root_add_223_n33), .ZN(
        DP_add_2_root_add_0_root_add_223_n295) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U278 ( .A(
        DP_add_2_root_add_0_root_add_223_n59), .ZN(
        DP_add_2_root_add_0_root_add_223_n57) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U277 ( .A(
        DP_add_2_root_add_0_root_add_223_n127), .ZN(
        DP_add_2_root_add_0_root_add_223_n125) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U276 ( .A1(
        DP_add_2_root_add_0_root_add_223_n58), .A2(
        DP_add_2_root_add_0_root_add_223_n42), .ZN(
        DP_add_2_root_add_0_root_add_223_n40) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U275 ( .A1(
        DP_add_2_root_add_0_root_add_223_n99), .A2(
        DP_add_2_root_add_0_root_add_223_n126), .ZN(
        DP_add_2_root_add_0_root_add_223_n97) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U274 ( .A(
        DP_add_2_root_add_0_root_add_223_n110), .ZN(
        DP_add_2_root_add_0_root_add_223_n108) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U273 ( .A(
        DP_add_2_root_add_0_root_add_223_n60), .ZN(
        DP_add_2_root_add_0_root_add_223_n58) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U272 ( .A(
        DP_add_2_root_add_0_root_add_223_n128), .ZN(
        DP_add_2_root_add_0_root_add_223_n126) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U271 ( .A(
        DP_add_2_root_add_0_root_add_223_n111), .ZN(
        DP_add_2_root_add_0_root_add_223_n109) );
  AOI21_X1 DP_add_2_root_add_0_root_add_223_U270 ( .B1(
        DP_add_2_root_add_0_root_add_223_n127), .B2(
        DP_add_2_root_add_0_root_add_223_n108), .A(
        DP_add_2_root_add_0_root_add_223_n109), .ZN(
        DP_add_2_root_add_0_root_add_223_n107) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U269 ( .A(
        DP_add_2_root_add_0_root_add_223_n58), .ZN(
        DP_add_2_root_add_0_root_add_223_n56) );
  INV_X1 DP_add_2_root_add_0_root_add_223_U268 ( .A(
        DP_add_2_root_add_0_root_add_223_n126), .ZN(
        DP_add_2_root_add_0_root_add_223_n124) );
  NAND2_X1 DP_add_2_root_add_0_root_add_223_U267 ( .A1(
        DP_add_2_root_add_0_root_add_223_n126), .A2(
        DP_add_2_root_add_0_root_add_223_n108), .ZN(
        DP_add_2_root_add_0_root_add_223_n106) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U266 ( .A1(DP_pipe11[22]), .A2(
        DP_pipe13[22]), .ZN(DP_add_2_root_add_0_root_add_223_n37) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U265 ( .A1(DP_pipe11[1]), .A2(
        DP_pipe13[1]), .ZN(DP_add_2_root_add_0_root_add_223_n187) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U264 ( .A1(DP_pipe11[8]), .A2(
        DP_pipe13[8]), .ZN(DP_add_2_root_add_0_root_add_223_n153) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U263 ( .A1(DP_pipe11[6]), .A2(
        DP_pipe13[6]), .ZN(DP_add_2_root_add_0_root_add_223_n164) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U262 ( .A1(DP_pipe11[16]), .A2(
        DP_pipe13[16]), .ZN(DP_add_2_root_add_0_root_add_223_n85) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U261 ( .A1(DP_pipe11[2]), .A2(
        DP_pipe13[2]), .ZN(DP_add_2_root_add_0_root_add_223_n183) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U260 ( .A1(DP_pipe11[9]), .A2(
        DP_pipe13[9]), .ZN(DP_add_2_root_add_0_root_add_223_n150) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U259 ( .A1(DP_pipe11[21]), .A2(
        DP_pipe13[21]), .ZN(DP_add_2_root_add_0_root_add_223_n46) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U258 ( .A1(DP_pipe11[3]), .A2(
        DP_pipe13[3]), .ZN(DP_add_2_root_add_0_root_add_223_n180) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U257 ( .A1(DP_pipe11[5]), .A2(
        DP_pipe13[5]), .ZN(DP_add_2_root_add_0_root_add_223_n169) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U256 ( .A1(DP_pipe11[7]), .A2(
        DP_pipe13[7]), .ZN(DP_add_2_root_add_0_root_add_223_n161) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U255 ( .A1(DP_pipe11[11]), .A2(
        DP_pipe13[11]), .ZN(DP_add_2_root_add_0_root_add_223_n132) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U254 ( .A1(DP_pipe11[13]), .A2(
        DP_pipe13[13]), .ZN(DP_add_2_root_add_0_root_add_223_n114) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U253 ( .A1(DP_pipe11[15]), .A2(
        DP_pipe13[15]), .ZN(DP_add_2_root_add_0_root_add_223_n94) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U252 ( .A1(DP_pipe11[17]), .A2(
        DP_pipe13[17]), .ZN(DP_add_2_root_add_0_root_add_223_n82) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U251 ( .A1(DP_pipe11[19]), .A2(
        DP_pipe13[19]), .ZN(DP_add_2_root_add_0_root_add_223_n64) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U250 ( .A1(DP_pipe11[20]), .A2(
        DP_pipe13[20]), .ZN(DP_add_2_root_add_0_root_add_223_n53) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U249 ( .A1(DP_pipe11[18]), .A2(
        DP_pipe13[18]), .ZN(DP_add_2_root_add_0_root_add_223_n71) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U248 ( .A1(DP_pipe11[12]), .A2(
        DP_pipe13[12]), .ZN(DP_add_2_root_add_0_root_add_223_n121) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U247 ( .A1(DP_pipe11[4]), .A2(
        DP_pipe13[4]), .ZN(DP_add_2_root_add_0_root_add_223_n174) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U246 ( .A1(DP_pipe11[14]), .A2(
        DP_pipe13[14]), .ZN(DP_add_2_root_add_0_root_add_223_n103) );
  NOR2_X1 DP_add_2_root_add_0_root_add_223_U245 ( .A1(DP_pipe11[10]), .A2(
        DP_pipe13[10]), .ZN(DP_add_2_root_add_0_root_add_223_n139) );
  OR2_X1 DP_add_2_root_add_0_root_add_223_U244 ( .A1(DP_pipe11[0]), .A2(
        DP_pipe13[0]), .ZN(DP_add_2_root_add_0_root_add_223_n294) );
  AND2_X1 DP_add_2_root_add_0_root_add_223_U243 ( .A1(
        DP_add_2_root_add_0_root_add_223_n294), .A2(
        DP_add_2_root_add_0_root_add_223_n190), .ZN(DP_ff_0_) );
  INV_X2 DP_add_2_root_add_0_root_add_223_U242 ( .A(
        DP_add_2_root_add_0_root_add_223_n156), .ZN(
        DP_add_2_root_add_0_root_add_223_n155) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U465 ( .B1(
        DP_add_1_root_add_0_root_add_223_n180), .B2(
        DP_add_1_root_add_0_root_add_223_n184), .A(
        DP_add_1_root_add_0_root_add_223_n181), .ZN(
        DP_add_1_root_add_0_root_add_223_n179) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U464 ( .A1(
        DP_add_1_root_add_0_root_add_223_n183), .A2(
        DP_add_1_root_add_0_root_add_223_n180), .ZN(
        DP_add_1_root_add_0_root_add_223_n178) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U463 ( .A1(DP_pipe10[3]), .A2(
        DP_pipe12[3]), .ZN(DP_add_1_root_add_0_root_add_223_n181) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U462 ( .A1(DP_pipe10[1]), .A2(
        DP_pipe12[1]), .ZN(DP_add_1_root_add_0_root_add_223_n188) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U461 ( .A1(DP_pipe10[7]), .A2(
        DP_pipe12[7]), .ZN(DP_add_1_root_add_0_root_add_223_n162) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U460 ( .A1(DP_pipe10[5]), .A2(
        DP_pipe12[5]), .ZN(DP_add_1_root_add_0_root_add_223_n170) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U459 ( .A1(DP_pipe10[9]), .A2(
        DP_pipe12[9]), .ZN(DP_add_1_root_add_0_root_add_223_n151) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U458 ( .A1(DP_pipe10[11]), .A2(
        DP_pipe12[11]), .ZN(DP_add_1_root_add_0_root_add_223_n133) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U457 ( .A1(DP_pipe10[21]), .A2(
        DP_pipe12[21]), .ZN(DP_add_1_root_add_0_root_add_223_n47) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U456 ( .A1(DP_pipe10[19]), .A2(
        DP_pipe12[19]), .ZN(DP_add_1_root_add_0_root_add_223_n65) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U455 ( .A1(DP_pipe10[17]), .A2(
        DP_pipe12[17]), .ZN(DP_add_1_root_add_0_root_add_223_n83) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U454 ( .A1(DP_pipe10[15]), .A2(
        DP_pipe12[15]), .ZN(DP_add_1_root_add_0_root_add_223_n95) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U453 ( .A1(DP_pipe10[13]), .A2(
        DP_pipe12[13]), .ZN(DP_add_1_root_add_0_root_add_223_n115) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U452 ( .A1(DP_pipe10[22]), .A2(
        DP_pipe12[22]), .ZN(DP_add_1_root_add_0_root_add_223_n38) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U451 ( .A1(DP_pipe10[2]), .A2(
        DP_pipe12[2]), .ZN(DP_add_1_root_add_0_root_add_223_n184) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U450 ( .A1(DP_pipe10[0]), .A2(
        DP_pipe12[0]), .ZN(DP_add_1_root_add_0_root_add_223_n190) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U449 ( .A1(DP_pipe10[6]), .A2(
        DP_pipe12[6]), .ZN(DP_add_1_root_add_0_root_add_223_n165) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U448 ( .A1(DP_pipe10[8]), .A2(
        DP_pipe12[8]), .ZN(DP_add_1_root_add_0_root_add_223_n154) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U447 ( .A1(DP_pipe10[4]), .A2(
        DP_pipe12[4]), .ZN(DP_add_1_root_add_0_root_add_223_n175) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U446 ( .A1(DP_pipe10[10]), .A2(
        DP_pipe12[10]), .ZN(DP_add_1_root_add_0_root_add_223_n140) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U445 ( .A1(DP_pipe10[16]), .A2(
        DP_pipe12[16]), .ZN(DP_add_1_root_add_0_root_add_223_n86) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U444 ( .A1(DP_pipe10[14]), .A2(
        DP_pipe12[14]), .ZN(DP_add_1_root_add_0_root_add_223_n104) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U443 ( .A1(DP_pipe10[20]), .A2(
        DP_pipe12[20]), .ZN(DP_add_1_root_add_0_root_add_223_n54) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U442 ( .A1(DP_pipe10[18]), .A2(
        DP_pipe12[18]), .ZN(DP_add_1_root_add_0_root_add_223_n72) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U441 ( .A1(DP_pipe10[12]), .A2(
        DP_pipe12[12]), .ZN(DP_add_1_root_add_0_root_add_223_n122) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U440 ( .A1(DP_pipe10[3]), .A2(
        DP_pipe12[3]), .ZN(DP_add_1_root_add_0_root_add_223_n180) );
  OR2_X1 DP_add_1_root_add_0_root_add_223_U439 ( .A1(DP_pipe10[23]), .A2(
        DP_pipe12[23]), .ZN(DP_add_1_root_add_0_root_add_223_n296) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U438 ( .A1(DP_pipe10[23]), .A2(
        DP_pipe12[23]), .ZN(DP_add_1_root_add_0_root_add_223_n27) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U437 ( .B1(
        DP_add_1_root_add_0_root_add_223_n1), .B2(
        DP_add_1_root_add_0_root_add_223_n295), .A(
        DP_add_1_root_add_0_root_add_223_n30), .ZN(
        DP_add_1_root_add_0_root_add_223_n28) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U436 ( .A1(
        DP_add_1_root_add_0_root_add_223_n296), .A2(
        DP_add_1_root_add_0_root_add_223_n27), .ZN(
        DP_add_1_root_add_0_root_add_223_n2) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U435 ( .A(
        DP_add_1_root_add_0_root_add_223_n28), .B(
        DP_add_1_root_add_0_root_add_223_n2), .ZN(DP_ff_part_23_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U434 ( .A(
        DP_add_1_root_add_0_root_add_223_n38), .ZN(
        DP_add_1_root_add_0_root_add_223_n36) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U433 ( .B1(
        DP_add_1_root_add_0_root_add_223_n45), .B2(
        DP_add_1_root_add_0_root_add_223_n35), .A(
        DP_add_1_root_add_0_root_add_223_n36), .ZN(
        DP_add_1_root_add_0_root_add_223_n34) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U432 ( .B1(
        DP_add_1_root_add_0_root_add_223_n61), .B2(
        DP_add_1_root_add_0_root_add_223_n33), .A(
        DP_add_1_root_add_0_root_add_223_n34), .ZN(
        DP_add_1_root_add_0_root_add_223_n32) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U431 ( .A(
        DP_add_1_root_add_0_root_add_223_n32), .ZN(
        DP_add_1_root_add_0_root_add_223_n30) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U430 ( .A(
        DP_add_1_root_add_0_root_add_223_n175), .ZN(
        DP_add_1_root_add_0_root_add_223_n173) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U429 ( .A(
        DP_add_1_root_add_0_root_add_223_n187), .ZN(
        DP_add_1_root_add_0_root_add_223_n213) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U428 ( .A1(
        DP_add_1_root_add_0_root_add_223_n213), .A2(
        DP_add_1_root_add_0_root_add_223_n188), .ZN(
        DP_add_1_root_add_0_root_add_223_n24) );
  XOR2_X1 DP_add_1_root_add_0_root_add_223_U427 ( .A(
        DP_add_1_root_add_0_root_add_223_n24), .B(
        DP_add_1_root_add_0_root_add_223_n190), .Z(DP_ff_part_1_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U426 ( .A(
        DP_add_1_root_add_0_root_add_223_n183), .ZN(
        DP_add_1_root_add_0_root_add_223_n212) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U425 ( .A1(
        DP_add_1_root_add_0_root_add_223_n212), .A2(
        DP_add_1_root_add_0_root_add_223_n184), .ZN(
        DP_add_1_root_add_0_root_add_223_n23) );
  XOR2_X1 DP_add_1_root_add_0_root_add_223_U424 ( .A(
        DP_add_1_root_add_0_root_add_223_n185), .B(
        DP_add_1_root_add_0_root_add_223_n23), .Z(DP_ff_part_2_) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U423 ( .A1(
        DP_add_1_root_add_0_root_add_223_n172), .A2(
        DP_add_1_root_add_0_root_add_223_n175), .ZN(
        DP_add_1_root_add_0_root_add_223_n21) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U422 ( .A(
        DP_add_1_root_add_0_root_add_223_n176), .B(
        DP_add_1_root_add_0_root_add_223_n21), .ZN(DP_ff_part_4_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U421 ( .A(
        DP_add_1_root_add_0_root_add_223_n103), .ZN(
        DP_add_1_root_add_0_root_add_223_n102) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U420 ( .A(
        DP_add_1_root_add_0_root_add_223_n102), .ZN(
        DP_add_1_root_add_0_root_add_223_n101) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U419 ( .A(
        DP_add_1_root_add_0_root_add_223_n174), .ZN(
        DP_add_1_root_add_0_root_add_223_n172) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U418 ( .A(
        DP_add_1_root_add_0_root_add_223_n37), .ZN(
        DP_add_1_root_add_0_root_add_223_n35) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U417 ( .A(
        DP_add_1_root_add_0_root_add_223_n139), .ZN(
        DP_add_1_root_add_0_root_add_223_n137) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U416 ( .A(
        DP_add_1_root_add_0_root_add_223_n53), .ZN(
        DP_add_1_root_add_0_root_add_223_n51) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U415 ( .A(
        DP_add_1_root_add_0_root_add_223_n71), .ZN(
        DP_add_1_root_add_0_root_add_223_n69) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U414 ( .A(
        DP_add_1_root_add_0_root_add_223_n121), .ZN(
        DP_add_1_root_add_0_root_add_223_n119) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U413 ( .B1(
        DP_add_1_root_add_0_root_add_223_n161), .B2(
        DP_add_1_root_add_0_root_add_223_n165), .A(
        DP_add_1_root_add_0_root_add_223_n162), .ZN(
        DP_add_1_root_add_0_root_add_223_n160) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U412 ( .A(
        DP_add_1_root_add_0_root_add_223_n72), .ZN(
        DP_add_1_root_add_0_root_add_223_n70) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U411 ( .B1(
        DP_add_1_root_add_0_root_add_223_n77), .B2(
        DP_add_1_root_add_0_root_add_223_n69), .A(
        DP_add_1_root_add_0_root_add_223_n70), .ZN(
        DP_add_1_root_add_0_root_add_223_n68) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U410 ( .A(
        DP_add_1_root_add_0_root_add_223_n54), .ZN(
        DP_add_1_root_add_0_root_add_223_n52) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U409 ( .B1(
        DP_add_1_root_add_0_root_add_223_n59), .B2(
        DP_add_1_root_add_0_root_add_223_n51), .A(
        DP_add_1_root_add_0_root_add_223_n52), .ZN(
        DP_add_1_root_add_0_root_add_223_n50) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U408 ( .A(
        DP_add_1_root_add_0_root_add_223_n140), .ZN(
        DP_add_1_root_add_0_root_add_223_n138) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U407 ( .B1(
        DP_add_1_root_add_0_root_add_223_n145), .B2(
        DP_add_1_root_add_0_root_add_223_n137), .A(
        DP_add_1_root_add_0_root_add_223_n138), .ZN(
        DP_add_1_root_add_0_root_add_223_n136) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U406 ( .A(
        DP_add_1_root_add_0_root_add_223_n122), .ZN(
        DP_add_1_root_add_0_root_add_223_n120) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U405 ( .B1(
        DP_add_1_root_add_0_root_add_223_n127), .B2(
        DP_add_1_root_add_0_root_add_223_n119), .A(
        DP_add_1_root_add_0_root_add_223_n120), .ZN(
        DP_add_1_root_add_0_root_add_223_n118) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U404 ( .B1(
        DP_add_1_root_add_0_root_add_223_n111), .B2(
        DP_add_1_root_add_0_root_add_223_n101), .A(
        DP_add_1_root_add_0_root_add_223_n104), .ZN(
        DP_add_1_root_add_0_root_add_223_n100) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U403 ( .B1(
        DP_add_1_root_add_0_root_add_223_n99), .B2(
        DP_add_1_root_add_0_root_add_223_n127), .A(
        DP_add_1_root_add_0_root_add_223_n100), .ZN(
        DP_add_1_root_add_0_root_add_223_n98) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U402 ( .B1(
        DP_add_1_root_add_0_root_add_223_n94), .B2(
        DP_add_1_root_add_0_root_add_223_n104), .A(
        DP_add_1_root_add_0_root_add_223_n95), .ZN(
        DP_add_1_root_add_0_root_add_223_n93) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U401 ( .B1(
        DP_add_1_root_add_0_root_add_223_n92), .B2(
        DP_add_1_root_add_0_root_add_223_n113), .A(
        DP_add_1_root_add_0_root_add_223_n93), .ZN(
        DP_add_1_root_add_0_root_add_223_n91) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U400 ( .A1(
        DP_add_1_root_add_0_root_add_223_n153), .A2(
        DP_add_1_root_add_0_root_add_223_n150), .ZN(
        DP_add_1_root_add_0_root_add_223_n148) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U399 ( .A1(
        DP_add_1_root_add_0_root_add_223_n53), .A2(
        DP_add_1_root_add_0_root_add_223_n46), .ZN(
        DP_add_1_root_add_0_root_add_223_n44) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U398 ( .A1(
        DP_add_1_root_add_0_root_add_223_n121), .A2(
        DP_add_1_root_add_0_root_add_223_n114), .ZN(
        DP_add_1_root_add_0_root_add_223_n112) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U397 ( .A1(
        DP_add_1_root_add_0_root_add_223_n85), .A2(
        DP_add_1_root_add_0_root_add_223_n82), .ZN(
        DP_add_1_root_add_0_root_add_223_n80) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U396 ( .A1(
        DP_add_1_root_add_0_root_add_223_n139), .A2(
        DP_add_1_root_add_0_root_add_223_n132), .ZN(
        DP_add_1_root_add_0_root_add_223_n130) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U395 ( .A1(
        DP_add_1_root_add_0_root_add_223_n103), .A2(
        DP_add_1_root_add_0_root_add_223_n94), .ZN(
        DP_add_1_root_add_0_root_add_223_n92) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U394 ( .A1(
        DP_add_1_root_add_0_root_add_223_n71), .A2(
        DP_add_1_root_add_0_root_add_223_n64), .ZN(
        DP_add_1_root_add_0_root_add_223_n62) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U393 ( .A1(
        DP_add_1_root_add_0_root_add_223_n174), .A2(
        DP_add_1_root_add_0_root_add_223_n169), .ZN(
        DP_add_1_root_add_0_root_add_223_n167) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U392 ( .A1(
        DP_add_1_root_add_0_root_add_223_n164), .A2(
        DP_add_1_root_add_0_root_add_223_n161), .ZN(
        DP_add_1_root_add_0_root_add_223_n159) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U391 ( .B1(
        DP_add_1_root_add_0_root_add_223_n159), .B2(
        DP_add_1_root_add_0_root_add_223_n168), .A(
        DP_add_1_root_add_0_root_add_223_n160), .ZN(
        DP_add_1_root_add_0_root_add_223_n158) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U390 ( .A1(
        DP_add_1_root_add_0_root_add_223_n167), .A2(
        DP_add_1_root_add_0_root_add_223_n159), .ZN(
        DP_add_1_root_add_0_root_add_223_n157) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U389 ( .B1(
        DP_add_1_root_add_0_root_add_223_n177), .B2(
        DP_add_1_root_add_0_root_add_223_n157), .A(
        DP_add_1_root_add_0_root_add_223_n158), .ZN(
        DP_add_1_root_add_0_root_add_223_n156) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U388 ( .B1(
        DP_add_1_root_add_0_root_add_223_n46), .B2(
        DP_add_1_root_add_0_root_add_223_n54), .A(
        DP_add_1_root_add_0_root_add_223_n47), .ZN(
        DP_add_1_root_add_0_root_add_223_n45) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U387 ( .B1(
        DP_add_1_root_add_0_root_add_223_n169), .B2(
        DP_add_1_root_add_0_root_add_223_n175), .A(
        DP_add_1_root_add_0_root_add_223_n170), .ZN(
        DP_add_1_root_add_0_root_add_223_n168) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U386 ( .B1(
        DP_add_1_root_add_0_root_add_223_n187), .B2(
        DP_add_1_root_add_0_root_add_223_n190), .A(
        DP_add_1_root_add_0_root_add_223_n188), .ZN(
        DP_add_1_root_add_0_root_add_223_n186) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U385 ( .B1(
        DP_add_1_root_add_0_root_add_223_n150), .B2(
        DP_add_1_root_add_0_root_add_223_n154), .A(
        DP_add_1_root_add_0_root_add_223_n151), .ZN(
        DP_add_1_root_add_0_root_add_223_n149) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U384 ( .B1(
        DP_add_1_root_add_0_root_add_223_n82), .B2(
        DP_add_1_root_add_0_root_add_223_n86), .A(
        DP_add_1_root_add_0_root_add_223_n83), .ZN(
        DP_add_1_root_add_0_root_add_223_n81) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U383 ( .B1(
        DP_add_1_root_add_0_root_add_223_n114), .B2(
        DP_add_1_root_add_0_root_add_223_n122), .A(
        DP_add_1_root_add_0_root_add_223_n115), .ZN(
        DP_add_1_root_add_0_root_add_223_n113) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U382 ( .B1(
        DP_add_1_root_add_0_root_add_223_n178), .B2(
        DP_add_1_root_add_0_root_add_223_n186), .A(
        DP_add_1_root_add_0_root_add_223_n179), .ZN(
        DP_add_1_root_add_0_root_add_223_n177) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U381 ( .B1(
        DP_add_1_root_add_0_root_add_223_n64), .B2(
        DP_add_1_root_add_0_root_add_223_n72), .A(
        DP_add_1_root_add_0_root_add_223_n65), .ZN(
        DP_add_1_root_add_0_root_add_223_n63) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U380 ( .B1(
        DP_add_1_root_add_0_root_add_223_n62), .B2(
        DP_add_1_root_add_0_root_add_223_n81), .A(
        DP_add_1_root_add_0_root_add_223_n63), .ZN(
        DP_add_1_root_add_0_root_add_223_n61) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U379 ( .B1(
        DP_add_1_root_add_0_root_add_223_n132), .B2(
        DP_add_1_root_add_0_root_add_223_n140), .A(
        DP_add_1_root_add_0_root_add_223_n133), .ZN(
        DP_add_1_root_add_0_root_add_223_n131) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U378 ( .B1(
        DP_add_1_root_add_0_root_add_223_n130), .B2(
        DP_add_1_root_add_0_root_add_223_n149), .A(
        DP_add_1_root_add_0_root_add_223_n131), .ZN(
        DP_add_1_root_add_0_root_add_223_n129) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U377 ( .A(
        DP_add_1_root_add_0_root_add_223_n82), .ZN(
        DP_add_1_root_add_0_root_add_223_n197) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U376 ( .B1(
        DP_add_1_root_add_0_root_add_223_n1), .B2(
        DP_add_1_root_add_0_root_add_223_n85), .A(
        DP_add_1_root_add_0_root_add_223_n86), .ZN(
        DP_add_1_root_add_0_root_add_223_n84) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U375 ( .A1(
        DP_add_1_root_add_0_root_add_223_n197), .A2(
        DP_add_1_root_add_0_root_add_223_n83), .ZN(
        DP_add_1_root_add_0_root_add_223_n8) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U374 ( .A(
        DP_add_1_root_add_0_root_add_223_n84), .B(
        DP_add_1_root_add_0_root_add_223_n8), .ZN(DP_ff_part_17_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U373 ( .A(
        DP_add_1_root_add_0_root_add_223_n64), .ZN(
        DP_add_1_root_add_0_root_add_223_n195) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U372 ( .B1(
        DP_add_1_root_add_0_root_add_223_n1), .B2(
        DP_add_1_root_add_0_root_add_223_n67), .A(
        DP_add_1_root_add_0_root_add_223_n68), .ZN(
        DP_add_1_root_add_0_root_add_223_n66) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U371 ( .A1(
        DP_add_1_root_add_0_root_add_223_n195), .A2(
        DP_add_1_root_add_0_root_add_223_n65), .ZN(
        DP_add_1_root_add_0_root_add_223_n6) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U370 ( .A(
        DP_add_1_root_add_0_root_add_223_n66), .B(
        DP_add_1_root_add_0_root_add_223_n6), .ZN(DP_ff_part_19_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U369 ( .A(
        DP_add_1_root_add_0_root_add_223_n46), .ZN(
        DP_add_1_root_add_0_root_add_223_n193) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U368 ( .B1(
        DP_add_1_root_add_0_root_add_223_n1), .B2(
        DP_add_1_root_add_0_root_add_223_n49), .A(
        DP_add_1_root_add_0_root_add_223_n50), .ZN(
        DP_add_1_root_add_0_root_add_223_n48) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U367 ( .A1(
        DP_add_1_root_add_0_root_add_223_n193), .A2(
        DP_add_1_root_add_0_root_add_223_n47), .ZN(
        DP_add_1_root_add_0_root_add_223_n4) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U366 ( .A(
        DP_add_1_root_add_0_root_add_223_n48), .B(
        DP_add_1_root_add_0_root_add_223_n4), .ZN(DP_ff_part_21_) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U365 ( .B1(
        DP_add_1_root_add_0_root_add_223_n1), .B2(
        DP_add_1_root_add_0_root_add_223_n74), .A(
        DP_add_1_root_add_0_root_add_223_n75), .ZN(
        DP_add_1_root_add_0_root_add_223_n73) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U364 ( .A1(
        DP_add_1_root_add_0_root_add_223_n69), .A2(
        DP_add_1_root_add_0_root_add_223_n72), .ZN(
        DP_add_1_root_add_0_root_add_223_n7) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U363 ( .A(
        DP_add_1_root_add_0_root_add_223_n73), .B(
        DP_add_1_root_add_0_root_add_223_n7), .ZN(DP_ff_part_18_) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U362 ( .B1(
        DP_add_1_root_add_0_root_add_223_n1), .B2(
        DP_add_1_root_add_0_root_add_223_n56), .A(
        DP_add_1_root_add_0_root_add_223_n57), .ZN(
        DP_add_1_root_add_0_root_add_223_n55) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U361 ( .A1(
        DP_add_1_root_add_0_root_add_223_n51), .A2(
        DP_add_1_root_add_0_root_add_223_n54), .ZN(
        DP_add_1_root_add_0_root_add_223_n5) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U360 ( .A(
        DP_add_1_root_add_0_root_add_223_n55), .B(
        DP_add_1_root_add_0_root_add_223_n5), .ZN(DP_ff_part_20_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U359 ( .A(
        DP_add_1_root_add_0_root_add_223_n37), .ZN(
        DP_add_1_root_add_0_root_add_223_n192) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U358 ( .B1(
        DP_add_1_root_add_0_root_add_223_n1), .B2(
        DP_add_1_root_add_0_root_add_223_n40), .A(
        DP_add_1_root_add_0_root_add_223_n41), .ZN(
        DP_add_1_root_add_0_root_add_223_n39) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U357 ( .A1(
        DP_add_1_root_add_0_root_add_223_n192), .A2(
        DP_add_1_root_add_0_root_add_223_n38), .ZN(
        DP_add_1_root_add_0_root_add_223_n3) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U356 ( .A(
        DP_add_1_root_add_0_root_add_223_n39), .B(
        DP_add_1_root_add_0_root_add_223_n3), .ZN(DP_ff_part_22_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U355 ( .A(
        DP_add_1_root_add_0_root_add_223_n94), .ZN(
        DP_add_1_root_add_0_root_add_223_n199) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U354 ( .B1(
        DP_add_1_root_add_0_root_add_223_n155), .B2(
        DP_add_1_root_add_0_root_add_223_n97), .A(
        DP_add_1_root_add_0_root_add_223_n98), .ZN(
        DP_add_1_root_add_0_root_add_223_n96) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U353 ( .A1(
        DP_add_1_root_add_0_root_add_223_n199), .A2(
        DP_add_1_root_add_0_root_add_223_n95), .ZN(
        DP_add_1_root_add_0_root_add_223_n10) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U352 ( .A(
        DP_add_1_root_add_0_root_add_223_n96), .B(
        DP_add_1_root_add_0_root_add_223_n10), .ZN(DP_ff_part_15_) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U351 ( .B1(
        DP_add_1_root_add_0_root_add_223_n155), .B2(
        DP_add_1_root_add_0_root_add_223_n142), .A(
        DP_add_1_root_add_0_root_add_223_n143), .ZN(
        DP_add_1_root_add_0_root_add_223_n141) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U350 ( .A1(
        DP_add_1_root_add_0_root_add_223_n137), .A2(
        DP_add_1_root_add_0_root_add_223_n140), .ZN(
        DP_add_1_root_add_0_root_add_223_n15) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U349 ( .A(
        DP_add_1_root_add_0_root_add_223_n141), .B(
        DP_add_1_root_add_0_root_add_223_n15), .ZN(DP_ff_part_10_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U348 ( .A(
        DP_add_1_root_add_0_root_add_223_n114), .ZN(
        DP_add_1_root_add_0_root_add_223_n201) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U347 ( .B1(
        DP_add_1_root_add_0_root_add_223_n155), .B2(
        DP_add_1_root_add_0_root_add_223_n117), .A(
        DP_add_1_root_add_0_root_add_223_n118), .ZN(
        DP_add_1_root_add_0_root_add_223_n116) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U346 ( .A1(
        DP_add_1_root_add_0_root_add_223_n201), .A2(
        DP_add_1_root_add_0_root_add_223_n115), .ZN(
        DP_add_1_root_add_0_root_add_223_n12) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U345 ( .A(
        DP_add_1_root_add_0_root_add_223_n116), .B(
        DP_add_1_root_add_0_root_add_223_n12), .ZN(DP_ff_part_13_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U344 ( .A(
        DP_add_1_root_add_0_root_add_223_n132), .ZN(
        DP_add_1_root_add_0_root_add_223_n203) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U343 ( .B1(
        DP_add_1_root_add_0_root_add_223_n155), .B2(
        DP_add_1_root_add_0_root_add_223_n135), .A(
        DP_add_1_root_add_0_root_add_223_n136), .ZN(
        DP_add_1_root_add_0_root_add_223_n134) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U342 ( .A1(
        DP_add_1_root_add_0_root_add_223_n203), .A2(
        DP_add_1_root_add_0_root_add_223_n133), .ZN(
        DP_add_1_root_add_0_root_add_223_n14) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U341 ( .A(
        DP_add_1_root_add_0_root_add_223_n134), .B(
        DP_add_1_root_add_0_root_add_223_n14), .ZN(DP_ff_part_11_) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U340 ( .B1(
        DP_add_1_root_add_0_root_add_223_n155), .B2(
        DP_add_1_root_add_0_root_add_223_n124), .A(
        DP_add_1_root_add_0_root_add_223_n125), .ZN(
        DP_add_1_root_add_0_root_add_223_n123) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U339 ( .A1(
        DP_add_1_root_add_0_root_add_223_n119), .A2(
        DP_add_1_root_add_0_root_add_223_n122), .ZN(
        DP_add_1_root_add_0_root_add_223_n13) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U338 ( .A(
        DP_add_1_root_add_0_root_add_223_n123), .B(
        DP_add_1_root_add_0_root_add_223_n13), .ZN(DP_ff_part_12_) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U337 ( .B1(
        DP_add_1_root_add_0_root_add_223_n155), .B2(
        DP_add_1_root_add_0_root_add_223_n106), .A(
        DP_add_1_root_add_0_root_add_223_n107), .ZN(
        DP_add_1_root_add_0_root_add_223_n105) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U336 ( .A1(
        DP_add_1_root_add_0_root_add_223_n102), .A2(
        DP_add_1_root_add_0_root_add_223_n104), .ZN(
        DP_add_1_root_add_0_root_add_223_n11) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U335 ( .A(
        DP_add_1_root_add_0_root_add_223_n105), .B(
        DP_add_1_root_add_0_root_add_223_n11), .ZN(DP_ff_part_14_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U334 ( .A(
        DP_add_1_root_add_0_root_add_223_n180), .ZN(
        DP_add_1_root_add_0_root_add_223_n211) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U333 ( .B1(
        DP_add_1_root_add_0_root_add_223_n185), .B2(
        DP_add_1_root_add_0_root_add_223_n183), .A(
        DP_add_1_root_add_0_root_add_223_n184), .ZN(
        DP_add_1_root_add_0_root_add_223_n182) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U332 ( .A1(
        DP_add_1_root_add_0_root_add_223_n211), .A2(
        DP_add_1_root_add_0_root_add_223_n181), .ZN(
        DP_add_1_root_add_0_root_add_223_n22) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U331 ( .A(
        DP_add_1_root_add_0_root_add_223_n182), .B(
        DP_add_1_root_add_0_root_add_223_n22), .ZN(DP_ff_part_3_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U330 ( .A(
        DP_add_1_root_add_0_root_add_223_n161), .ZN(
        DP_add_1_root_add_0_root_add_223_n207) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U329 ( .B1(
        DP_add_1_root_add_0_root_add_223_n166), .B2(
        DP_add_1_root_add_0_root_add_223_n164), .A(
        DP_add_1_root_add_0_root_add_223_n165), .ZN(
        DP_add_1_root_add_0_root_add_223_n163) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U328 ( .A1(
        DP_add_1_root_add_0_root_add_223_n207), .A2(
        DP_add_1_root_add_0_root_add_223_n162), .ZN(
        DP_add_1_root_add_0_root_add_223_n18) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U327 ( .A(
        DP_add_1_root_add_0_root_add_223_n163), .B(
        DP_add_1_root_add_0_root_add_223_n18), .ZN(DP_ff_part_7_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U326 ( .A(
        DP_add_1_root_add_0_root_add_223_n150), .ZN(
        DP_add_1_root_add_0_root_add_223_n205) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U325 ( .B1(
        DP_add_1_root_add_0_root_add_223_n155), .B2(
        DP_add_1_root_add_0_root_add_223_n153), .A(
        DP_add_1_root_add_0_root_add_223_n154), .ZN(
        DP_add_1_root_add_0_root_add_223_n152) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U324 ( .A1(
        DP_add_1_root_add_0_root_add_223_n205), .A2(
        DP_add_1_root_add_0_root_add_223_n151), .ZN(
        DP_add_1_root_add_0_root_add_223_n16) );
  XNOR2_X1 DP_add_1_root_add_0_root_add_223_U323 ( .A(
        DP_add_1_root_add_0_root_add_223_n152), .B(
        DP_add_1_root_add_0_root_add_223_n16), .ZN(DP_ff_part_9_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U322 ( .A(
        DP_add_1_root_add_0_root_add_223_n169), .ZN(
        DP_add_1_root_add_0_root_add_223_n209) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U321 ( .B1(
        DP_add_1_root_add_0_root_add_223_n176), .B2(
        DP_add_1_root_add_0_root_add_223_n172), .A(
        DP_add_1_root_add_0_root_add_223_n173), .ZN(
        DP_add_1_root_add_0_root_add_223_n171) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U320 ( .A1(
        DP_add_1_root_add_0_root_add_223_n209), .A2(
        DP_add_1_root_add_0_root_add_223_n170), .ZN(
        DP_add_1_root_add_0_root_add_223_n20) );
  XOR2_X1 DP_add_1_root_add_0_root_add_223_U319 ( .A(
        DP_add_1_root_add_0_root_add_223_n171), .B(
        DP_add_1_root_add_0_root_add_223_n20), .Z(DP_ff_part_5_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U318 ( .A(
        DP_add_1_root_add_0_root_add_223_n164), .ZN(
        DP_add_1_root_add_0_root_add_223_n208) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U317 ( .A1(
        DP_add_1_root_add_0_root_add_223_n208), .A2(
        DP_add_1_root_add_0_root_add_223_n165), .ZN(
        DP_add_1_root_add_0_root_add_223_n19) );
  XOR2_X1 DP_add_1_root_add_0_root_add_223_U316 ( .A(
        DP_add_1_root_add_0_root_add_223_n166), .B(
        DP_add_1_root_add_0_root_add_223_n19), .Z(DP_ff_part_6_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U315 ( .A(
        DP_add_1_root_add_0_root_add_223_n153), .ZN(
        DP_add_1_root_add_0_root_add_223_n206) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U314 ( .A1(
        DP_add_1_root_add_0_root_add_223_n206), .A2(
        DP_add_1_root_add_0_root_add_223_n154), .ZN(
        DP_add_1_root_add_0_root_add_223_n17) );
  XOR2_X1 DP_add_1_root_add_0_root_add_223_U313 ( .A(
        DP_add_1_root_add_0_root_add_223_n155), .B(
        DP_add_1_root_add_0_root_add_223_n17), .Z(DP_ff_part_8_) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U312 ( .A(
        DP_add_1_root_add_0_root_add_223_n85), .ZN(
        DP_add_1_root_add_0_root_add_223_n198) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U311 ( .A1(
        DP_add_1_root_add_0_root_add_223_n198), .A2(
        DP_add_1_root_add_0_root_add_223_n86), .ZN(
        DP_add_1_root_add_0_root_add_223_n9) );
  XOR2_X1 DP_add_1_root_add_0_root_add_223_U310 ( .A(
        DP_add_1_root_add_0_root_add_223_n1), .B(
        DP_add_1_root_add_0_root_add_223_n9), .Z(DP_ff_part_16_) );
  OAI21_X1 DP_add_1_root_add_0_root_add_223_U309 ( .B1(
        DP_add_1_root_add_0_root_add_223_n129), .B2(
        DP_add_1_root_add_0_root_add_223_n90), .A(
        DP_add_1_root_add_0_root_add_223_n91), .ZN(
        DP_add_1_root_add_0_root_add_223_n89) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U308 ( .A1(
        DP_add_1_root_add_0_root_add_223_n128), .A2(
        DP_add_1_root_add_0_root_add_223_n90), .ZN(
        DP_add_1_root_add_0_root_add_223_n88) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U307 ( .B1(
        DP_add_1_root_add_0_root_add_223_n156), .B2(
        DP_add_1_root_add_0_root_add_223_n88), .A(
        DP_add_1_root_add_0_root_add_223_n89), .ZN(
        DP_add_1_root_add_0_root_add_223_n87) );
  BUF_X1 DP_add_1_root_add_0_root_add_223_U306 ( .A(
        DP_add_1_root_add_0_root_add_223_n87), .Z(
        DP_add_1_root_add_0_root_add_223_n1) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U305 ( .A1(
        DP_add_1_root_add_0_root_add_223_n80), .A2(
        DP_add_1_root_add_0_root_add_223_n69), .ZN(
        DP_add_1_root_add_0_root_add_223_n67) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U304 ( .A1(
        DP_add_1_root_add_0_root_add_223_n148), .A2(
        DP_add_1_root_add_0_root_add_223_n137), .ZN(
        DP_add_1_root_add_0_root_add_223_n135) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U303 ( .A1(
        DP_add_1_root_add_0_root_add_223_n58), .A2(
        DP_add_1_root_add_0_root_add_223_n51), .ZN(
        DP_add_1_root_add_0_root_add_223_n49) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U302 ( .A1(
        DP_add_1_root_add_0_root_add_223_n126), .A2(
        DP_add_1_root_add_0_root_add_223_n119), .ZN(
        DP_add_1_root_add_0_root_add_223_n117) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U301 ( .A(
        DP_add_1_root_add_0_root_add_223_n149), .ZN(
        DP_add_1_root_add_0_root_add_223_n147) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U300 ( .A(
        DP_add_1_root_add_0_root_add_223_n147), .ZN(
        DP_add_1_root_add_0_root_add_223_n145) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U299 ( .A(
        DP_add_1_root_add_0_root_add_223_n81), .ZN(
        DP_add_1_root_add_0_root_add_223_n79) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U298 ( .A(
        DP_add_1_root_add_0_root_add_223_n79), .ZN(
        DP_add_1_root_add_0_root_add_223_n77) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U297 ( .A(
        DP_add_1_root_add_0_root_add_223_n44), .ZN(
        DP_add_1_root_add_0_root_add_223_n43) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U296 ( .A(
        DP_add_1_root_add_0_root_add_223_n43), .ZN(
        DP_add_1_root_add_0_root_add_223_n42) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U295 ( .A(
        DP_add_1_root_add_0_root_add_223_n186), .ZN(
        DP_add_1_root_add_0_root_add_223_n185) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U294 ( .A(
        DP_add_1_root_add_0_root_add_223_n112), .ZN(
        DP_add_1_root_add_0_root_add_223_n110) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U293 ( .A(
        DP_add_1_root_add_0_root_add_223_n113), .ZN(
        DP_add_1_root_add_0_root_add_223_n111) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U292 ( .A1(
        DP_add_1_root_add_0_root_add_223_n44), .A2(
        DP_add_1_root_add_0_root_add_223_n35), .ZN(
        DP_add_1_root_add_0_root_add_223_n33) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U291 ( .A1(
        DP_add_1_root_add_0_root_add_223_n80), .A2(
        DP_add_1_root_add_0_root_add_223_n62), .ZN(
        DP_add_1_root_add_0_root_add_223_n60) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U290 ( .A1(
        DP_add_1_root_add_0_root_add_223_n148), .A2(
        DP_add_1_root_add_0_root_add_223_n130), .ZN(
        DP_add_1_root_add_0_root_add_223_n128) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U289 ( .A(
        DP_add_1_root_add_0_root_add_223_n177), .ZN(
        DP_add_1_root_add_0_root_add_223_n176) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U288 ( .A1(
        DP_add_1_root_add_0_root_add_223_n112), .A2(
        DP_add_1_root_add_0_root_add_223_n92), .ZN(
        DP_add_1_root_add_0_root_add_223_n90) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U287 ( .A(
        DP_add_1_root_add_0_root_add_223_n61), .ZN(
        DP_add_1_root_add_0_root_add_223_n59) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U286 ( .A(
        DP_add_1_root_add_0_root_add_223_n129), .ZN(
        DP_add_1_root_add_0_root_add_223_n127) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U285 ( .B1(
        DP_add_1_root_add_0_root_add_223_n59), .B2(
        DP_add_1_root_add_0_root_add_223_n42), .A(
        DP_add_1_root_add_0_root_add_223_n45), .ZN(
        DP_add_1_root_add_0_root_add_223_n41) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U284 ( .A1(
        DP_add_1_root_add_0_root_add_223_n110), .A2(
        DP_add_1_root_add_0_root_add_223_n101), .ZN(
        DP_add_1_root_add_0_root_add_223_n99) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U283 ( .B1(
        DP_add_1_root_add_0_root_add_223_n176), .B2(
        DP_add_1_root_add_0_root_add_223_n167), .A(
        DP_add_1_root_add_0_root_add_223_n168), .ZN(
        DP_add_1_root_add_0_root_add_223_n166) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U282 ( .A(
        DP_add_1_root_add_0_root_add_223_n77), .ZN(
        DP_add_1_root_add_0_root_add_223_n75) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U281 ( .A(
        DP_add_1_root_add_0_root_add_223_n145), .ZN(
        DP_add_1_root_add_0_root_add_223_n143) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U280 ( .A(
        DP_add_1_root_add_0_root_add_223_n80), .ZN(
        DP_add_1_root_add_0_root_add_223_n74) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U279 ( .A(
        DP_add_1_root_add_0_root_add_223_n148), .ZN(
        DP_add_1_root_add_0_root_add_223_n142) );
  OR2_X1 DP_add_1_root_add_0_root_add_223_U278 ( .A1(
        DP_add_1_root_add_0_root_add_223_n60), .A2(
        DP_add_1_root_add_0_root_add_223_n33), .ZN(
        DP_add_1_root_add_0_root_add_223_n295) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U277 ( .A(
        DP_add_1_root_add_0_root_add_223_n59), .ZN(
        DP_add_1_root_add_0_root_add_223_n57) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U276 ( .A(
        DP_add_1_root_add_0_root_add_223_n127), .ZN(
        DP_add_1_root_add_0_root_add_223_n125) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U275 ( .A1(
        DP_add_1_root_add_0_root_add_223_n58), .A2(
        DP_add_1_root_add_0_root_add_223_n42), .ZN(
        DP_add_1_root_add_0_root_add_223_n40) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U274 ( .A1(
        DP_add_1_root_add_0_root_add_223_n99), .A2(
        DP_add_1_root_add_0_root_add_223_n126), .ZN(
        DP_add_1_root_add_0_root_add_223_n97) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U273 ( .A(
        DP_add_1_root_add_0_root_add_223_n110), .ZN(
        DP_add_1_root_add_0_root_add_223_n108) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U272 ( .A(
        DP_add_1_root_add_0_root_add_223_n60), .ZN(
        DP_add_1_root_add_0_root_add_223_n58) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U271 ( .A(
        DP_add_1_root_add_0_root_add_223_n128), .ZN(
        DP_add_1_root_add_0_root_add_223_n126) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U270 ( .A(
        DP_add_1_root_add_0_root_add_223_n111), .ZN(
        DP_add_1_root_add_0_root_add_223_n109) );
  AOI21_X1 DP_add_1_root_add_0_root_add_223_U269 ( .B1(
        DP_add_1_root_add_0_root_add_223_n127), .B2(
        DP_add_1_root_add_0_root_add_223_n108), .A(
        DP_add_1_root_add_0_root_add_223_n109), .ZN(
        DP_add_1_root_add_0_root_add_223_n107) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U268 ( .A(
        DP_add_1_root_add_0_root_add_223_n58), .ZN(
        DP_add_1_root_add_0_root_add_223_n56) );
  INV_X1 DP_add_1_root_add_0_root_add_223_U267 ( .A(
        DP_add_1_root_add_0_root_add_223_n126), .ZN(
        DP_add_1_root_add_0_root_add_223_n124) );
  NAND2_X1 DP_add_1_root_add_0_root_add_223_U266 ( .A1(
        DP_add_1_root_add_0_root_add_223_n126), .A2(
        DP_add_1_root_add_0_root_add_223_n108), .ZN(
        DP_add_1_root_add_0_root_add_223_n106) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U265 ( .A1(DP_pipe10[22]), .A2(
        DP_pipe12[22]), .ZN(DP_add_1_root_add_0_root_add_223_n37) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U264 ( .A1(DP_pipe10[1]), .A2(
        DP_pipe12[1]), .ZN(DP_add_1_root_add_0_root_add_223_n187) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U263 ( .A1(DP_pipe10[8]), .A2(
        DP_pipe12[8]), .ZN(DP_add_1_root_add_0_root_add_223_n153) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U262 ( .A1(DP_pipe10[2]), .A2(
        DP_pipe12[2]), .ZN(DP_add_1_root_add_0_root_add_223_n183) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U261 ( .A1(DP_pipe10[6]), .A2(
        DP_pipe12[6]), .ZN(DP_add_1_root_add_0_root_add_223_n164) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U260 ( .A1(DP_pipe10[16]), .A2(
        DP_pipe12[16]), .ZN(DP_add_1_root_add_0_root_add_223_n85) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U259 ( .A1(DP_pipe10[9]), .A2(
        DP_pipe12[9]), .ZN(DP_add_1_root_add_0_root_add_223_n150) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U258 ( .A1(DP_pipe10[5]), .A2(
        DP_pipe12[5]), .ZN(DP_add_1_root_add_0_root_add_223_n169) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U257 ( .A1(DP_pipe10[7]), .A2(
        DP_pipe12[7]), .ZN(DP_add_1_root_add_0_root_add_223_n161) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U256 ( .A1(DP_pipe10[11]), .A2(
        DP_pipe12[11]), .ZN(DP_add_1_root_add_0_root_add_223_n132) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U255 ( .A1(DP_pipe10[21]), .A2(
        DP_pipe12[21]), .ZN(DP_add_1_root_add_0_root_add_223_n46) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U254 ( .A1(DP_pipe10[13]), .A2(
        DP_pipe12[13]), .ZN(DP_add_1_root_add_0_root_add_223_n114) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U253 ( .A1(DP_pipe10[15]), .A2(
        DP_pipe12[15]), .ZN(DP_add_1_root_add_0_root_add_223_n94) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U252 ( .A1(DP_pipe10[17]), .A2(
        DP_pipe12[17]), .ZN(DP_add_1_root_add_0_root_add_223_n82) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U251 ( .A1(DP_pipe10[19]), .A2(
        DP_pipe12[19]), .ZN(DP_add_1_root_add_0_root_add_223_n64) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U250 ( .A1(DP_pipe10[4]), .A2(
        DP_pipe12[4]), .ZN(DP_add_1_root_add_0_root_add_223_n174) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U249 ( .A1(DP_pipe10[10]), .A2(
        DP_pipe12[10]), .ZN(DP_add_1_root_add_0_root_add_223_n139) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U248 ( .A1(DP_pipe10[20]), .A2(
        DP_pipe12[20]), .ZN(DP_add_1_root_add_0_root_add_223_n53) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U247 ( .A1(DP_pipe10[18]), .A2(
        DP_pipe12[18]), .ZN(DP_add_1_root_add_0_root_add_223_n71) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U246 ( .A1(DP_pipe10[12]), .A2(
        DP_pipe12[12]), .ZN(DP_add_1_root_add_0_root_add_223_n121) );
  NOR2_X1 DP_add_1_root_add_0_root_add_223_U245 ( .A1(DP_pipe10[14]), .A2(
        DP_pipe12[14]), .ZN(DP_add_1_root_add_0_root_add_223_n103) );
  OR2_X1 DP_add_1_root_add_0_root_add_223_U244 ( .A1(DP_pipe10[0]), .A2(
        DP_pipe12[0]), .ZN(DP_add_1_root_add_0_root_add_223_n294) );
  AND2_X1 DP_add_1_root_add_0_root_add_223_U243 ( .A1(
        DP_add_1_root_add_0_root_add_223_n294), .A2(
        DP_add_1_root_add_0_root_add_223_n190), .ZN(DP_ff_part_0_) );
  INV_X2 DP_add_1_root_add_0_root_add_223_U242 ( .A(
        DP_add_1_root_add_0_root_add_223_n156), .ZN(
        DP_add_1_root_add_0_root_add_223_n155) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U465 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n153), .A2(
        DP_add_1_root_sub_0_root_sub_217_n150), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n148) );
  XOR2_X1 DP_add_1_root_sub_0_root_sub_217_U464 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n1), .B(
        DP_add_1_root_sub_0_root_sub_217_n9), .Z(DP_fb_16_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U463 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n177), .B2(
        DP_add_1_root_sub_0_root_sub_217_n157), .A(
        DP_add_1_root_sub_0_root_sub_217_n158), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n156) );
  OR2_X1 DP_add_1_root_sub_0_root_sub_217_U462 ( .A1(DP_ret0[23]), .A2(
        DP_ret1[23]), .ZN(DP_add_1_root_sub_0_root_sub_217_n297) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U461 ( .A1(DP_ret0[9]), .A2(
        DP_ret1[9]), .ZN(DP_add_1_root_sub_0_root_sub_217_n151) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U460 ( .A1(DP_ret0[3]), .A2(
        DP_ret1[3]), .ZN(DP_add_1_root_sub_0_root_sub_217_n181) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U459 ( .A1(DP_ret0[1]), .A2(
        DP_ret1[1]), .ZN(DP_add_1_root_sub_0_root_sub_217_n188) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U458 ( .A1(DP_ret0[7]), .A2(
        DP_ret1[7]), .ZN(DP_add_1_root_sub_0_root_sub_217_n162) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U457 ( .A1(DP_ret0[5]), .A2(
        DP_ret1[5]), .ZN(DP_add_1_root_sub_0_root_sub_217_n170) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U456 ( .A1(DP_ret0[11]), .A2(
        DP_ret1[11]), .ZN(DP_add_1_root_sub_0_root_sub_217_n133) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U455 ( .A1(DP_ret0[21]), .A2(
        DP_ret1[21]), .ZN(DP_add_1_root_sub_0_root_sub_217_n47) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U454 ( .A1(DP_ret0[19]), .A2(
        DP_ret1[19]), .ZN(DP_add_1_root_sub_0_root_sub_217_n65) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U453 ( .A1(DP_ret0[13]), .A2(
        DP_ret1[13]), .ZN(DP_add_1_root_sub_0_root_sub_217_n115) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U452 ( .A1(DP_ret0[17]), .A2(
        DP_ret1[17]), .ZN(DP_add_1_root_sub_0_root_sub_217_n83) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U451 ( .A1(DP_ret0[15]), .A2(
        DP_ret1[15]), .ZN(DP_add_1_root_sub_0_root_sub_217_n95) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U450 ( .A1(DP_ret0[22]), .A2(
        DP_ret1[22]), .ZN(DP_add_1_root_sub_0_root_sub_217_n38) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U449 ( .A1(DP_ret0[0]), .A2(
        DP_ret1[0]), .ZN(DP_add_1_root_sub_0_root_sub_217_n190) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U448 ( .A1(DP_ret0[8]), .A2(
        DP_ret1[8]), .ZN(DP_add_1_root_sub_0_root_sub_217_n154) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U447 ( .A1(DP_ret0[6]), .A2(
        DP_ret1[6]), .ZN(DP_add_1_root_sub_0_root_sub_217_n165) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U446 ( .A1(DP_ret0[2]), .A2(
        DP_ret1[2]), .ZN(DP_add_1_root_sub_0_root_sub_217_n184) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U445 ( .A1(DP_ret0[4]), .A2(
        DP_ret1[4]), .ZN(DP_add_1_root_sub_0_root_sub_217_n175) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U444 ( .A1(DP_ret0[10]), .A2(
        DP_ret1[10]), .ZN(DP_add_1_root_sub_0_root_sub_217_n140) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U443 ( .A1(DP_ret0[14]), .A2(
        DP_ret1[14]), .ZN(DP_add_1_root_sub_0_root_sub_217_n104) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U442 ( .A1(DP_ret0[16]), .A2(
        DP_ret1[16]), .ZN(DP_add_1_root_sub_0_root_sub_217_n86) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U441 ( .A1(DP_ret0[20]), .A2(
        DP_ret1[20]), .ZN(DP_add_1_root_sub_0_root_sub_217_n54) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U440 ( .A1(DP_ret0[18]), .A2(
        DP_ret1[18]), .ZN(DP_add_1_root_sub_0_root_sub_217_n72) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U439 ( .A1(DP_ret0[12]), .A2(
        DP_ret1[12]), .ZN(DP_add_1_root_sub_0_root_sub_217_n122) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U438 ( .A1(DP_ret0[9]), .A2(
        DP_ret1[9]), .ZN(DP_add_1_root_sub_0_root_sub_217_n150) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U437 ( .A1(DP_ret0[23]), .A2(
        DP_ret1[23]), .ZN(DP_add_1_root_sub_0_root_sub_217_n27) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U436 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n1), .B2(
        DP_add_1_root_sub_0_root_sub_217_n296), .A(
        DP_add_1_root_sub_0_root_sub_217_n30), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n28) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U435 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n297), .A2(
        DP_add_1_root_sub_0_root_sub_217_n27), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n2) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U434 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n28), .B(
        DP_add_1_root_sub_0_root_sub_217_n2), .ZN(DP_fb_23_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U433 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n38), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n36) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U432 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n45), .B2(
        DP_add_1_root_sub_0_root_sub_217_n293), .A(
        DP_add_1_root_sub_0_root_sub_217_n36), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n34) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U431 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n61), .B2(
        DP_add_1_root_sub_0_root_sub_217_n33), .A(
        DP_add_1_root_sub_0_root_sub_217_n34), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n32) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U430 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n32), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n30) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U429 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n175), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n173) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U428 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n187), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n213) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U427 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n213), .A2(
        DP_add_1_root_sub_0_root_sub_217_n188), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n24) );
  XOR2_X1 DP_add_1_root_sub_0_root_sub_217_U426 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n24), .B(
        DP_add_1_root_sub_0_root_sub_217_n190), .Z(DP_fb_1_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U425 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n183), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n212) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U424 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n212), .A2(
        DP_add_1_root_sub_0_root_sub_217_n184), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n23) );
  XOR2_X1 DP_add_1_root_sub_0_root_sub_217_U423 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n185), .B(
        DP_add_1_root_sub_0_root_sub_217_n23), .Z(DP_fb_2_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U422 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n132), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n203) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U421 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n46), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n193) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U420 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n114), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n201) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U419 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n64), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n195) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U418 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n94), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n199) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U417 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n82), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n197) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U416 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n1), .B2(
        DP_add_1_root_sub_0_root_sub_217_n74), .A(
        DP_add_1_root_sub_0_root_sub_217_n75), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n73) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U415 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n69), .A2(
        DP_add_1_root_sub_0_root_sub_217_n72), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n7) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U414 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n73), .B(
        DP_add_1_root_sub_0_root_sub_217_n7), .ZN(DP_fb_18_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U413 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n103), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n102) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U412 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n102), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n101) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U411 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n174), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n172) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U410 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n1), .B2(
        DP_add_1_root_sub_0_root_sub_217_n40), .A(
        DP_add_1_root_sub_0_root_sub_217_n41), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n39) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U409 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n293), .A2(
        DP_add_1_root_sub_0_root_sub_217_n38), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n3) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U408 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n39), .B(
        DP_add_1_root_sub_0_root_sub_217_n3), .ZN(DP_fb_22_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U407 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n1), .B2(
        DP_add_1_root_sub_0_root_sub_217_n56), .A(
        DP_add_1_root_sub_0_root_sub_217_n57), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n55) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U406 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n51), .A2(
        DP_add_1_root_sub_0_root_sub_217_n54), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n5) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U405 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n55), .B(
        DP_add_1_root_sub_0_root_sub_217_n5), .ZN(DP_fb_20_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U404 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n1), .B2(
        DP_add_1_root_sub_0_root_sub_217_n49), .A(
        DP_add_1_root_sub_0_root_sub_217_n50), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n48) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U403 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n193), .A2(
        DP_add_1_root_sub_0_root_sub_217_n47), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n4) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U402 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n48), .B(
        DP_add_1_root_sub_0_root_sub_217_n4), .ZN(DP_fb_21_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U401 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n155), .B2(
        DP_add_1_root_sub_0_root_sub_217_n106), .A(
        DP_add_1_root_sub_0_root_sub_217_n107), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n105) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U400 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n102), .A2(
        DP_add_1_root_sub_0_root_sub_217_n104), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n11) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U399 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n105), .B(
        DP_add_1_root_sub_0_root_sub_217_n11), .ZN(DP_fb_14_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U398 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n155), .B2(
        DP_add_1_root_sub_0_root_sub_217_n117), .A(
        DP_add_1_root_sub_0_root_sub_217_n118), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n116) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U397 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n201), .A2(
        DP_add_1_root_sub_0_root_sub_217_n115), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n12) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U396 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n116), .B(
        DP_add_1_root_sub_0_root_sub_217_n12), .ZN(DP_fb_13_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U395 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n1), .B2(
        DP_add_1_root_sub_0_root_sub_217_n67), .A(
        DP_add_1_root_sub_0_root_sub_217_n68), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n66) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U394 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n195), .A2(
        DP_add_1_root_sub_0_root_sub_217_n65), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n6) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U393 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n66), .B(
        DP_add_1_root_sub_0_root_sub_217_n6), .ZN(DP_fb_19_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U392 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n155), .B2(
        DP_add_1_root_sub_0_root_sub_217_n97), .A(
        DP_add_1_root_sub_0_root_sub_217_n98), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n96) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U391 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n199), .A2(
        DP_add_1_root_sub_0_root_sub_217_n95), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n10) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U390 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n96), .B(
        DP_add_1_root_sub_0_root_sub_217_n10), .ZN(DP_fb_15_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U389 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n1), .B2(
        DP_add_1_root_sub_0_root_sub_217_n85), .A(
        DP_add_1_root_sub_0_root_sub_217_n86), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n84) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U388 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n197), .A2(
        DP_add_1_root_sub_0_root_sub_217_n83), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n8) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U387 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n84), .B(
        DP_add_1_root_sub_0_root_sub_217_n8), .ZN(DP_fb_17_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U386 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n139), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n137) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U385 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n53), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n51) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U384 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n121), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n119) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U383 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n71), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n69) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U382 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n155), .B2(
        DP_add_1_root_sub_0_root_sub_217_n135), .A(
        DP_add_1_root_sub_0_root_sub_217_n136), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n134) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U381 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n203), .A2(
        DP_add_1_root_sub_0_root_sub_217_n133), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n14) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U380 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n134), .B(
        DP_add_1_root_sub_0_root_sub_217_n14), .ZN(DP_fb_11_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U379 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n161), .B2(
        DP_add_1_root_sub_0_root_sub_217_n165), .A(
        DP_add_1_root_sub_0_root_sub_217_n162), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n160) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U378 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n132), .B2(
        DP_add_1_root_sub_0_root_sub_217_n140), .A(
        DP_add_1_root_sub_0_root_sub_217_n133), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n131) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U377 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n130), .B2(
        DP_add_1_root_sub_0_root_sub_217_n149), .A(
        DP_add_1_root_sub_0_root_sub_217_n131), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n129) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U376 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n54), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n52) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U375 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n59), .B2(
        DP_add_1_root_sub_0_root_sub_217_n51), .A(
        DP_add_1_root_sub_0_root_sub_217_n52), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n50) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U374 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n72), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n70) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U373 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n77), .B2(
        DP_add_1_root_sub_0_root_sub_217_n69), .A(
        DP_add_1_root_sub_0_root_sub_217_n70), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n68) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U372 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n122), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n120) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U371 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n127), .B2(
        DP_add_1_root_sub_0_root_sub_217_n119), .A(
        DP_add_1_root_sub_0_root_sub_217_n120), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n118) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U370 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n140), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n138) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U369 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n145), .B2(
        DP_add_1_root_sub_0_root_sub_217_n137), .A(
        DP_add_1_root_sub_0_root_sub_217_n138), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n136) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U368 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n111), .B2(
        DP_add_1_root_sub_0_root_sub_217_n101), .A(
        DP_add_1_root_sub_0_root_sub_217_n104), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n100) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U367 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n99), .B2(
        DP_add_1_root_sub_0_root_sub_217_n127), .A(
        DP_add_1_root_sub_0_root_sub_217_n100), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n98) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U366 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n94), .B2(
        DP_add_1_root_sub_0_root_sub_217_n104), .A(
        DP_add_1_root_sub_0_root_sub_217_n95), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n93) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U365 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n92), .B2(
        DP_add_1_root_sub_0_root_sub_217_n113), .A(
        DP_add_1_root_sub_0_root_sub_217_n93), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n91) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U364 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n85), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n198) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U363 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n198), .A2(
        DP_add_1_root_sub_0_root_sub_217_n86), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n9) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U362 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n53), .A2(
        DP_add_1_root_sub_0_root_sub_217_n46), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n44) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U361 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n121), .A2(
        DP_add_1_root_sub_0_root_sub_217_n114), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n112) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U360 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n85), .A2(
        DP_add_1_root_sub_0_root_sub_217_n82), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n80) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U359 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n139), .A2(
        DP_add_1_root_sub_0_root_sub_217_n132), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n130) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U358 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n103), .A2(
        DP_add_1_root_sub_0_root_sub_217_n94), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n92) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U357 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n71), .A2(
        DP_add_1_root_sub_0_root_sub_217_n64), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n62) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U356 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n174), .A2(
        DP_add_1_root_sub_0_root_sub_217_n169), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n167) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U355 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n180), .B2(
        DP_add_1_root_sub_0_root_sub_217_n184), .A(
        DP_add_1_root_sub_0_root_sub_217_n181), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n179) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U354 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n183), .A2(
        DP_add_1_root_sub_0_root_sub_217_n180), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n178) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U353 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n178), .B2(
        DP_add_1_root_sub_0_root_sub_217_n186), .A(
        DP_add_1_root_sub_0_root_sub_217_n179), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n177) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U352 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n46), .B2(
        DP_add_1_root_sub_0_root_sub_217_n54), .A(
        DP_add_1_root_sub_0_root_sub_217_n47), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n45) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U351 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n169), .B2(
        DP_add_1_root_sub_0_root_sub_217_n175), .A(
        DP_add_1_root_sub_0_root_sub_217_n170), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n168) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U350 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n187), .B2(
        DP_add_1_root_sub_0_root_sub_217_n190), .A(
        DP_add_1_root_sub_0_root_sub_217_n188), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n186) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U349 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n82), .B2(
        DP_add_1_root_sub_0_root_sub_217_n86), .A(
        DP_add_1_root_sub_0_root_sub_217_n83), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n81) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U348 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n114), .B2(
        DP_add_1_root_sub_0_root_sub_217_n122), .A(
        DP_add_1_root_sub_0_root_sub_217_n115), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n113) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U347 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n64), .B2(
        DP_add_1_root_sub_0_root_sub_217_n72), .A(
        DP_add_1_root_sub_0_root_sub_217_n65), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n63) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U346 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n62), .B2(
        DP_add_1_root_sub_0_root_sub_217_n81), .A(
        DP_add_1_root_sub_0_root_sub_217_n63), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n61) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U345 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n155), .B2(
        DP_add_1_root_sub_0_root_sub_217_n124), .A(
        DP_add_1_root_sub_0_root_sub_217_n125), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n123) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U344 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n119), .A2(
        DP_add_1_root_sub_0_root_sub_217_n122), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n13) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U343 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n123), .B(
        DP_add_1_root_sub_0_root_sub_217_n13), .ZN(DP_fb_12_) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U342 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n172), .A2(
        DP_add_1_root_sub_0_root_sub_217_n175), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n21) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U341 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n176), .B(
        DP_add_1_root_sub_0_root_sub_217_n21), .ZN(DP_fb_4_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U340 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n180), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n211) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U339 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n211), .A2(
        DP_add_1_root_sub_0_root_sub_217_n181), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n22) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U338 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n185), .B2(
        DP_add_1_root_sub_0_root_sub_217_n183), .A(
        DP_add_1_root_sub_0_root_sub_217_n184), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n182) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U337 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n182), .B(
        DP_add_1_root_sub_0_root_sub_217_n22), .ZN(DP_fb_3_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U336 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n150), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n205) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U335 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n155), .B2(
        DP_add_1_root_sub_0_root_sub_217_n153), .A(
        DP_add_1_root_sub_0_root_sub_217_n154), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n152) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U334 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n205), .A2(
        DP_add_1_root_sub_0_root_sub_217_n151), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n16) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U333 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n152), .B(
        DP_add_1_root_sub_0_root_sub_217_n16), .ZN(DP_fb_9_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U332 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n161), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n207) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U331 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n166), .B2(
        DP_add_1_root_sub_0_root_sub_217_n164), .A(
        DP_add_1_root_sub_0_root_sub_217_n165), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n163) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U330 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n207), .A2(
        DP_add_1_root_sub_0_root_sub_217_n162), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n18) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U329 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n163), .B(
        DP_add_1_root_sub_0_root_sub_217_n18), .ZN(DP_fb_7_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U328 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n155), .B2(
        DP_add_1_root_sub_0_root_sub_217_n142), .A(
        DP_add_1_root_sub_0_root_sub_217_n143), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n141) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U327 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n137), .A2(
        DP_add_1_root_sub_0_root_sub_217_n140), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n15) );
  XNOR2_X1 DP_add_1_root_sub_0_root_sub_217_U326 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n141), .B(
        DP_add_1_root_sub_0_root_sub_217_n15), .ZN(DP_fb_10_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U325 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n169), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n209) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U324 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n176), .B2(
        DP_add_1_root_sub_0_root_sub_217_n172), .A(
        DP_add_1_root_sub_0_root_sub_217_n173), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n171) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U323 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n209), .A2(
        DP_add_1_root_sub_0_root_sub_217_n170), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n20) );
  XOR2_X1 DP_add_1_root_sub_0_root_sub_217_U322 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n171), .B(
        DP_add_1_root_sub_0_root_sub_217_n20), .Z(DP_fb_5_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U321 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n153), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n206) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U320 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n206), .A2(
        DP_add_1_root_sub_0_root_sub_217_n154), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n17) );
  XOR2_X1 DP_add_1_root_sub_0_root_sub_217_U319 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n155), .B(
        DP_add_1_root_sub_0_root_sub_217_n17), .Z(DP_fb_8_) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U318 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n164), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n208) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U317 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n208), .A2(
        DP_add_1_root_sub_0_root_sub_217_n165), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n19) );
  XOR2_X1 DP_add_1_root_sub_0_root_sub_217_U316 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n166), .B(
        DP_add_1_root_sub_0_root_sub_217_n19), .Z(DP_fb_6_) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U315 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n150), .B2(
        DP_add_1_root_sub_0_root_sub_217_n154), .A(
        DP_add_1_root_sub_0_root_sub_217_n151), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n149) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U314 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n164), .A2(
        DP_add_1_root_sub_0_root_sub_217_n161), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n159) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U313 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n159), .B2(
        DP_add_1_root_sub_0_root_sub_217_n168), .A(
        DP_add_1_root_sub_0_root_sub_217_n160), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n158) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U312 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n167), .A2(
        DP_add_1_root_sub_0_root_sub_217_n159), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n157) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U311 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n44), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n43) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U310 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n43), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n42) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U309 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n76), .A2(
        DP_add_1_root_sub_0_root_sub_217_n69), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n67) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U308 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n58), .A2(
        DP_add_1_root_sub_0_root_sub_217_n51), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n49) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U307 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n126), .A2(
        DP_add_1_root_sub_0_root_sub_217_n119), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n117) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U306 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n148), .A2(
        DP_add_1_root_sub_0_root_sub_217_n137), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n135) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U305 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n80), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n78) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U304 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n78), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n76) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U303 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n81), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n79) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U302 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n79), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n77) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U301 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n149), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n147) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U300 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n147), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n145) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U299 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n186), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n185) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U298 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n112), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n110) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U297 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n113), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n111) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U296 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n177), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n176) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U295 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n44), .A2(
        DP_add_1_root_sub_0_root_sub_217_n293), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n33) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U294 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n80), .A2(
        DP_add_1_root_sub_0_root_sub_217_n62), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n60) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U293 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n112), .A2(
        DP_add_1_root_sub_0_root_sub_217_n92), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n90) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U292 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n61), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n59) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U291 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n129), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n127) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U290 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n148), .A2(
        DP_add_1_root_sub_0_root_sub_217_n130), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n128) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U289 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n59), .B2(
        DP_add_1_root_sub_0_root_sub_217_n42), .A(
        DP_add_1_root_sub_0_root_sub_217_n45), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n41) );
  OAI21_X1 DP_add_1_root_sub_0_root_sub_217_U288 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n129), .B2(
        DP_add_1_root_sub_0_root_sub_217_n90), .A(
        DP_add_1_root_sub_0_root_sub_217_n91), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n89) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U287 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n128), .A2(
        DP_add_1_root_sub_0_root_sub_217_n90), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n88) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U286 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n156), .B2(
        DP_add_1_root_sub_0_root_sub_217_n88), .A(
        DP_add_1_root_sub_0_root_sub_217_n89), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n87) );
  BUF_X1 DP_add_1_root_sub_0_root_sub_217_U285 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n87), .Z(
        DP_add_1_root_sub_0_root_sub_217_n1) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U284 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n110), .A2(
        DP_add_1_root_sub_0_root_sub_217_n101), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n99) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U283 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n176), .B2(
        DP_add_1_root_sub_0_root_sub_217_n167), .A(
        DP_add_1_root_sub_0_root_sub_217_n168), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n166) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U282 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n156), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n155) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U281 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n145), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n143) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U280 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n77), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n75) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U279 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n76), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n74) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U278 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n148), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n142) );
  OR2_X1 DP_add_1_root_sub_0_root_sub_217_U277 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n60), .A2(
        DP_add_1_root_sub_0_root_sub_217_n33), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n296) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U276 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n59), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n57) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U275 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n127), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n125) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U274 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n58), .A2(
        DP_add_1_root_sub_0_root_sub_217_n42), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n40) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U273 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n99), .A2(
        DP_add_1_root_sub_0_root_sub_217_n126), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n97) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U272 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n110), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n108) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U271 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n60), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n58) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U270 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n128), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n126) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U269 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n111), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n109) );
  AOI21_X1 DP_add_1_root_sub_0_root_sub_217_U268 ( .B1(
        DP_add_1_root_sub_0_root_sub_217_n127), .B2(
        DP_add_1_root_sub_0_root_sub_217_n108), .A(
        DP_add_1_root_sub_0_root_sub_217_n109), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n107) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U267 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n58), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n56) );
  INV_X1 DP_add_1_root_sub_0_root_sub_217_U266 ( .A(
        DP_add_1_root_sub_0_root_sub_217_n126), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n124) );
  NAND2_X1 DP_add_1_root_sub_0_root_sub_217_U265 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n126), .A2(
        DP_add_1_root_sub_0_root_sub_217_n108), .ZN(
        DP_add_1_root_sub_0_root_sub_217_n106) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U264 ( .A1(DP_ret0[16]), .A2(
        DP_ret1[16]), .ZN(DP_add_1_root_sub_0_root_sub_217_n85) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U263 ( .A1(DP_ret0[21]), .A2(
        DP_ret1[21]), .ZN(DP_add_1_root_sub_0_root_sub_217_n46) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U262 ( .A1(DP_ret0[17]), .A2(
        DP_ret1[17]), .ZN(DP_add_1_root_sub_0_root_sub_217_n82) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U261 ( .A1(DP_ret0[19]), .A2(
        DP_ret1[19]), .ZN(DP_add_1_root_sub_0_root_sub_217_n64) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U260 ( .A1(DP_ret0[20]), .A2(
        DP_ret1[20]), .ZN(DP_add_1_root_sub_0_root_sub_217_n53) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U259 ( .A1(DP_ret0[18]), .A2(
        DP_ret1[18]), .ZN(DP_add_1_root_sub_0_root_sub_217_n71) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U258 ( .A1(DP_ret0[1]), .A2(
        DP_ret1[1]), .ZN(DP_add_1_root_sub_0_root_sub_217_n187) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U257 ( .A1(DP_ret0[6]), .A2(
        DP_ret1[6]), .ZN(DP_add_1_root_sub_0_root_sub_217_n164) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U256 ( .A1(DP_ret0[8]), .A2(
        DP_ret1[8]), .ZN(DP_add_1_root_sub_0_root_sub_217_n153) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U255 ( .A1(DP_ret0[2]), .A2(
        DP_ret1[2]), .ZN(DP_add_1_root_sub_0_root_sub_217_n183) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U254 ( .A1(DP_ret0[3]), .A2(
        DP_ret1[3]), .ZN(DP_add_1_root_sub_0_root_sub_217_n180) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U253 ( .A1(DP_ret0[11]), .A2(
        DP_ret1[11]), .ZN(DP_add_1_root_sub_0_root_sub_217_n132) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U252 ( .A1(DP_ret0[7]), .A2(
        DP_ret1[7]), .ZN(DP_add_1_root_sub_0_root_sub_217_n161) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U251 ( .A1(DP_ret0[5]), .A2(
        DP_ret1[5]), .ZN(DP_add_1_root_sub_0_root_sub_217_n169) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U250 ( .A1(DP_ret0[15]), .A2(
        DP_ret1[15]), .ZN(DP_add_1_root_sub_0_root_sub_217_n94) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U249 ( .A1(DP_ret0[13]), .A2(
        DP_ret1[13]), .ZN(DP_add_1_root_sub_0_root_sub_217_n114) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U248 ( .A1(DP_ret0[10]), .A2(
        DP_ret1[10]), .ZN(DP_add_1_root_sub_0_root_sub_217_n139) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U247 ( .A1(DP_ret0[4]), .A2(
        DP_ret1[4]), .ZN(DP_add_1_root_sub_0_root_sub_217_n174) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U246 ( .A1(DP_ret0[12]), .A2(
        DP_ret1[12]), .ZN(DP_add_1_root_sub_0_root_sub_217_n121) );
  NOR2_X1 DP_add_1_root_sub_0_root_sub_217_U245 ( .A1(DP_ret0[14]), .A2(
        DP_ret1[14]), .ZN(DP_add_1_root_sub_0_root_sub_217_n103) );
  OR2_X1 DP_add_1_root_sub_0_root_sub_217_U244 ( .A1(DP_ret0[0]), .A2(
        DP_ret1[0]), .ZN(DP_add_1_root_sub_0_root_sub_217_n295) );
  AND2_X1 DP_add_1_root_sub_0_root_sub_217_U243 ( .A1(
        DP_add_1_root_sub_0_root_sub_217_n295), .A2(
        DP_add_1_root_sub_0_root_sub_217_n190), .ZN(DP_w_0_) );
  OR2_X1 DP_add_1_root_sub_0_root_sub_217_U242 ( .A1(DP_ret0[22]), .A2(
        DP_ret1[22]), .ZN(DP_add_1_root_sub_0_root_sub_217_n293) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U364 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n60), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n53), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n51) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U363 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n1), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n25), .A(
        DP_sub_0_root_sub_0_root_sub_217_n26), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n24) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U362 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n1), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n238), .A(
        DP_sub_0_root_sub_0_root_sub_217_n19), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n17) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U361 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n1), .B(
        DP_sub_0_root_sub_0_root_sub_217_n4), .Z(DP_w_21_) );
  AOI21_X1 DP_sub_0_root_sub_0_root_sub_217_U360 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n38), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n66), .A(
        DP_sub_0_root_sub_0_root_sub_217_n39), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n37) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U359 ( .A(DP_fb_12_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n159) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U358 ( .A(DP_x_11_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n161) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U357 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n153), .A2(DP_x_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n54) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U356 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n157), .A2(DP_x_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n90) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U355 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n151), .A2(DP_x_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n34) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U354 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n155), .A2(DP_x_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n72) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U353 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n159), .A2(DP_x_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n101) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U352 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n150), .A2(DP_x_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n26) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U351 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n154), .A2(DP_x_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n61) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U350 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n158), .A2(DP_x_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n93) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U349 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n152), .A2(DP_x_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n43) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U348 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n160), .A2(DP_x_0_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n104) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U347 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n156), .A2(DP_x_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n79) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U346 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n149), .A2(DP_x_11_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n23) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U345 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n153), .A2(DP_x_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n53) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U344 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n22), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n26), .A(
        DP_sub_0_root_sub_0_root_sub_217_n23), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n21) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U343 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n21), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n19) );
  OR2_X1 DP_sub_0_root_sub_0_root_sub_217_U342 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n161), .A2(DP_fb_23_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n239) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U341 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n103), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n148) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U340 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n148), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n104), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n14) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U339 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n105), .B(
        DP_sub_0_root_sub_0_root_sub_217_n14), .Z(DP_w_11_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U338 ( .A(DP_w_0_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n135) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U337 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n42), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n41) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U336 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n41), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n40) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U335 ( .A(DP_fb_18_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n153) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U334 ( .A(DP_fb_22_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n149) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U333 ( .A(DP_fb_20_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n151) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U332 ( .A(DP_fb_21_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n150) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U331 ( .A(DP_fb_14_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n157) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U330 ( .A(DP_fb_13_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n158) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U329 ( .A(DP_fb_19_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n152) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U328 ( .A(DP_fb_15_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n156) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U327 ( .A(DP_fb_17_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n154) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U326 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n60), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n58) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U325 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n78), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n76) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U324 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n94), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n45), .A(
        DP_sub_0_root_sub_0_root_sub_217_n46), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n44) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U323 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n41), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n43), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n6) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U322 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n44), .B(
        DP_sub_0_root_sub_0_root_sub_217_n6), .ZN(DP_w_19_) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U321 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n94), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n63), .A(
        DP_sub_0_root_sub_0_root_sub_217_n64), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n62) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U320 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n58), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n61), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n8) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U319 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n62), .B(
        DP_sub_0_root_sub_0_root_sub_217_n8), .ZN(DP_w_17_) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U318 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n94), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n81), .A(
        DP_sub_0_root_sub_0_root_sub_217_n82), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n80) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U317 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n76), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n79), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n10) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U316 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n80), .B(
        DP_sub_0_root_sub_0_root_sub_217_n10), .ZN(DP_w_15_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U315 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n53), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n141) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U314 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n94), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n56), .A(
        DP_sub_0_root_sub_0_root_sub_217_n57), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n55) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U313 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n141), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n54), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n7) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U312 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n55), .B(
        DP_sub_0_root_sub_0_root_sub_217_n7), .ZN(DP_w_18_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U311 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n71), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n143) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U310 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n94), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n74), .A(
        DP_sub_0_root_sub_0_root_sub_217_n75), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n73) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U309 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n143), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n72), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n9) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U308 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n73), .B(
        DP_sub_0_root_sub_0_root_sub_217_n9), .ZN(DP_w_16_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U307 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n33), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n139) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U306 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n36), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n94), .A(
        DP_sub_0_root_sub_0_root_sub_217_n37), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n35) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U305 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n139), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n34), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n5) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U304 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n35), .B(
        DP_sub_0_root_sub_0_root_sub_217_n5), .ZN(DP_w_20_) );
  OR2_X1 DP_sub_0_root_sub_0_root_sub_217_U303 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n25), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n22), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n238) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U302 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n161), .A2(DP_fb_23_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n16) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U301 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n239), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n16), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n2) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U300 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n17), .B(
        DP_sub_0_root_sub_0_root_sub_217_n2), .ZN(DP_w_23_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U299 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n100), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n147) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U298 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n105), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n103), .A(
        DP_sub_0_root_sub_0_root_sub_217_n104), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n102) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U297 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n147), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n101), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n13) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U296 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n102), .B(
        DP_sub_0_root_sub_0_root_sub_217_n13), .ZN(DP_w_12_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U295 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n89), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n145) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U294 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n94), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n92), .A(
        DP_sub_0_root_sub_0_root_sub_217_n93), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n91) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U293 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n145), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n90), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n11) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U292 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n91), .B(
        DP_sub_0_root_sub_0_root_sub_217_n11), .ZN(DP_w_14_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U291 ( .A(DP_fb_11_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n160) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U290 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n92), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n146) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U289 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n146), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n93), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n12) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U288 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n94), .B(
        DP_sub_0_root_sub_0_root_sub_217_n12), .Z(DP_w_13_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U287 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n79), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n77) );
  AOI21_X1 DP_sub_0_root_sub_0_root_sub_217_U286 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n84), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n76), .A(
        DP_sub_0_root_sub_0_root_sub_217_n77), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n75) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U285 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n61), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n59) );
  AOI21_X1 DP_sub_0_root_sub_0_root_sub_217_U284 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n66), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n58), .A(
        DP_sub_0_root_sub_0_root_sub_217_n59), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n57) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U283 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n33), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n43), .A(
        DP_sub_0_root_sub_0_root_sub_217_n34), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n32) );
  AOI21_X1 DP_sub_0_root_sub_0_root_sub_217_U282 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n31), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n52), .A(
        DP_sub_0_root_sub_0_root_sub_217_n32), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n30) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U281 ( .A(DP_fb_16_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n155) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U280 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n92), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n89), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n87) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U279 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n42), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n33), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n31) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U278 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n78), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n71), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n69) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U277 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n25), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n138) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U276 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n138), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n26), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n4) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U275 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n71), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n79), .A(
        DP_sub_0_root_sub_0_root_sub_217_n72), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n70) );
  AOI21_X1 DP_sub_0_root_sub_0_root_sub_217_U274 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n69), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n88), .A(
        DP_sub_0_root_sub_0_root_sub_217_n70), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n68) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U273 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n103), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n100), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n98) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U272 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n99), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n97) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U271 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n98), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n106), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n96) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U270 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n96), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n114), .A(
        DP_sub_0_root_sub_0_root_sub_217_n97), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n95) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U269 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n89), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n93), .A(
        DP_sub_0_root_sub_0_root_sub_217_n90), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n88) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U268 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n22), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n137) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U267 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n137), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n23), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n3) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U266 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n24), .B(
        DP_sub_0_root_sub_0_root_sub_217_n3), .ZN(DP_w_22_) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U265 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n100), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n104), .A(
        DP_sub_0_root_sub_0_root_sub_217_n101), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n99) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U264 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n53), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n61), .A(
        DP_sub_0_root_sub_0_root_sub_217_n54), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n52) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U263 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n50), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n40), .A(
        DP_sub_0_root_sub_0_root_sub_217_n43), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n39) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U262 ( .A(DP_fb_1_), .B(
        DP_sub_0_root_sub_0_root_sub_217_n135), .ZN(DP_w_1_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U261 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n65), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n58), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n56) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U260 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n87), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n76), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n74) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U259 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n88), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n86) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U258 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n86), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n84) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U257 ( .A(DP_fb_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n125) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U256 ( .A(DP_fb_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n131) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U255 ( .A(DP_fb_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n112) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U254 ( .A(DP_fb_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n119) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U253 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n52), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n50) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U252 ( .A(DP_fb_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n117) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U251 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n119), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n117), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n116) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U250 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n121), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n116), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n115) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U249 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n115), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n127), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n114) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U248 ( .A(DP_fb_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n134) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U247 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n134), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n135), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n133) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U246 ( .A(DP_fb_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n110) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U245 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n112), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n110), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n109) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U244 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n87), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n69), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n67) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U243 ( .A(DP_fb_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n122) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U242 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n125), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n122), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n121) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U241 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n51), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n49) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U240 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n125), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n124) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U239 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n126), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n124), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n123) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U238 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n123), .B(DP_fb_5_), .ZN(DP_w_5_) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U237 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n120), .B(DP_fb_6_), .ZN(DP_w_6_) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U236 ( .A(DP_fb_2_), .B(
        DP_sub_0_root_sub_0_root_sub_217_n132), .ZN(DP_w_2_) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U235 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n113), .B(DP_fb_8_), .ZN(DP_w_8_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U234 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n109), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n108) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U233 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n113), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n108), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n107) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U232 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n107), .B(DP_fb_10_), .Z(DP_w_10_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U231 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n132), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n131), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n130) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U230 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n130), .B(DP_fb_3_), .Z(DP_w_3_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U229 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n120), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n119), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n118) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U228 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n118), .B(DP_fb_7_), .Z(DP_w_7_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U227 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n113), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n112), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n111) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U226 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n111), .B(DP_fb_9_), .Z(DP_w_9_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U225 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n126), .B(DP_fb_4_), .Z(DP_w_4_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U224 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n51), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n31), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n29) );
  OAI21_X1 DP_sub_0_root_sub_0_root_sub_217_U223 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n68), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n29), .A(
        DP_sub_0_root_sub_0_root_sub_217_n30), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n28) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U222 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n67), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n29), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n27) );
  AOI21_X1 DP_sub_0_root_sub_0_root_sub_217_U221 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n27), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n95), .A(
        DP_sub_0_root_sub_0_root_sub_217_n28), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n1) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U220 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n109), .A2(DP_fb_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n106) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U219 ( .A(DP_fb_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n129) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U218 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n131), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n129), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n128) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U217 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n128), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n133), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n127) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U216 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n49), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n40), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n38) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U215 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n68), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n66) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U214 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n95), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n94) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U213 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n84), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n82) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U212 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n87), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n81) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U211 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n66), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n64) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U210 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n133), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n132) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U209 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n38), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n65), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n36) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U208 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n49), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n47) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U207 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n113), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n106), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n105) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U206 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n127), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n126) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U205 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n114), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n113) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U204 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n67), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n65) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U203 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n126), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n121), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n120) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U202 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n50), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n48) );
  AOI21_X1 DP_sub_0_root_sub_0_root_sub_217_U201 ( .B1(
        DP_sub_0_root_sub_0_root_sub_217_n66), .B2(
        DP_sub_0_root_sub_0_root_sub_217_n47), .A(
        DP_sub_0_root_sub_0_root_sub_217_n48), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n46) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_217_U200 ( .A(
        DP_sub_0_root_sub_0_root_sub_217_n65), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n63) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_217_U199 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n65), .A2(
        DP_sub_0_root_sub_0_root_sub_217_n47), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n45) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U198 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n150), .A2(DP_x_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n25) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U197 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n149), .A2(DP_x_11_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n22) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U196 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n158), .A2(DP_x_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n92) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U195 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n160), .A2(DP_x_0_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n103) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U194 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n151), .A2(DP_x_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n33) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U193 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n157), .A2(DP_x_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n89) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U192 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n159), .A2(DP_x_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n100) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U191 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n155), .A2(DP_x_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n71) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U190 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n152), .A2(DP_x_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n42) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U189 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n154), .A2(DP_x_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n60) );
  NOR2_X1 DP_sub_0_root_sub_0_root_sub_217_U188 ( .A1(
        DP_sub_0_root_sub_0_root_sub_217_n156), .A2(DP_x_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_217_n78) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U369 ( .B1(
        DP_add_0_root_add_0_root_add_223_n1), .B2(
        DP_add_0_root_add_0_root_add_223_n29), .A(
        DP_add_0_root_add_0_root_add_223_n30), .ZN(
        DP_add_0_root_add_0_root_add_223_n28) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U368 ( .A(
        DP_add_0_root_add_0_root_add_223_n28), .B(
        DP_add_0_root_add_0_root_add_223_n3), .ZN(DP_y_11_) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U367 ( .B1(
        DP_add_0_root_add_0_root_add_223_n121), .B2(
        DP_add_0_root_add_0_root_add_223_n129), .A(
        DP_add_0_root_add_0_root_add_223_n122), .ZN(
        DP_add_0_root_add_0_root_add_223_n120) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U366 ( .A1(
        DP_add_0_root_add_0_root_add_223_n128), .A2(
        DP_add_0_root_add_0_root_add_223_n121), .ZN(
        DP_add_0_root_add_0_root_add_223_n119) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U365 ( .A(
        DP_add_0_root_add_0_root_add_223_n71), .ZN(
        DP_add_0_root_add_0_root_add_223_n169) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U364 ( .B1(
        DP_add_0_root_add_0_root_add_223_n50), .B2(
        DP_add_0_root_add_0_root_add_223_n22), .A(
        DP_add_0_root_add_0_root_add_223_n23), .ZN(
        DP_add_0_root_add_0_root_add_223_n21) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U363 ( .A(
        DP_add_0_root_add_0_root_add_223_n50), .ZN(
        DP_add_0_root_add_0_root_add_223_n48) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U362 ( .A(
        DP_add_0_root_add_0_root_add_223_n37), .B(
        DP_add_0_root_add_0_root_add_223_n4), .ZN(DP_y_10_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U361 ( .A(
        DP_add_0_root_add_0_root_add_223_n44), .B(
        DP_add_0_root_add_0_root_add_223_n5), .ZN(DP_y_9_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U360 ( .A(
        DP_add_0_root_add_0_root_add_223_n55), .B(
        DP_add_0_root_add_0_root_add_223_n6), .ZN(DP_y_8_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U359 ( .A(
        DP_add_0_root_add_0_root_add_223_n62), .B(
        DP_add_0_root_add_0_root_add_223_n7), .ZN(DP_y_7_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U358 ( .A(
        DP_add_0_root_add_0_root_add_223_n73), .B(
        DP_add_0_root_add_0_root_add_223_n8), .ZN(DP_y_6_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_223_U357 ( .A(
        DP_add_0_root_add_0_root_add_223_n1), .B(
        DP_add_0_root_add_0_root_add_223_n9), .Z(DP_y_5_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U356 ( .A(
        DP_add_0_root_add_0_root_add_223_n85), .B(
        DP_add_0_root_add_0_root_add_223_n10), .ZN(DP_y_4_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U355 ( .A(
        DP_add_0_root_add_0_root_add_223_n94), .B(
        DP_add_0_root_add_0_root_add_223_n11), .ZN(DP_y_3_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U354 ( .A(
        DP_add_0_root_add_0_root_add_223_n105), .B(
        DP_add_0_root_add_0_root_add_223_n12), .ZN(DP_y_2_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U353 ( .A(
        DP_add_0_root_add_0_root_add_223_n112), .B(
        DP_add_0_root_add_0_root_add_223_n13), .ZN(DP_y_1_) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U352 ( .A(
        DP_add_0_root_add_0_root_add_223_n123), .B(
        DP_add_0_root_add_0_root_add_223_n14), .ZN(DP_y_0_) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U351 ( .A1(DP_ff_0_), .A2(
        DP_ff_part_0_), .ZN(DP_add_0_root_add_0_root_add_223_n162) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U350 ( .A1(DP_ff_1_), .A2(
        DP_ff_part_1_), .ZN(DP_add_0_root_add_0_root_add_223_n160) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U349 ( .A1(DP_ff_1_), .A2(
        DP_ff_part_1_), .ZN(DP_add_0_root_add_0_root_add_223_n161) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U348 ( .B1(
        DP_add_0_root_add_0_root_add_223_n160), .B2(
        DP_add_0_root_add_0_root_add_223_n162), .A(
        DP_add_0_root_add_0_root_add_223_n161), .ZN(
        DP_add_0_root_add_0_root_add_223_n159) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U347 ( .A1(DP_ff_23_), .A2(
        DP_ff_part_23_), .ZN(DP_add_0_root_add_0_root_add_223_n16) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U346 ( .B1(
        DP_add_0_root_add_0_root_add_223_n1), .B2(
        DP_add_0_root_add_0_root_add_223_n244), .A(
        DP_add_0_root_add_0_root_add_223_n19), .ZN(
        DP_add_0_root_add_0_root_add_223_n17) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U345 ( .A1(
        DP_add_0_root_add_0_root_add_223_n245), .A2(
        DP_add_0_root_add_0_root_add_223_n16), .ZN(
        DP_add_0_root_add_0_root_add_223_n2) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_223_U344 ( .A(
        DP_add_0_root_add_0_root_add_223_n17), .B(
        DP_add_0_root_add_0_root_add_223_n2), .ZN(DP_y_23) );
  OR2_X1 DP_add_0_root_add_0_root_add_223_U343 ( .A1(DP_ff_23_), .A2(
        DP_ff_part_23_), .ZN(DP_add_0_root_add_0_root_add_223_n245) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U342 ( .A1(DP_ff_17_), .A2(
        DP_ff_part_17_), .ZN(DP_add_0_root_add_0_root_add_223_n72) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U341 ( .A1(DP_ff_10_), .A2(
        DP_ff_part_10_), .ZN(DP_add_0_root_add_0_root_add_223_n129) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U340 ( .A1(DP_ff_11_), .A2(
        DP_ff_part_11_), .ZN(DP_add_0_root_add_0_root_add_223_n122) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U339 ( .A1(DP_ff_4_), .A2(
        DP_ff_part_4_), .ZN(DP_add_0_root_add_0_root_add_223_n150) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U338 ( .A1(
        DP_add_0_root_add_0_root_add_223_n150), .A2(
        DP_add_0_root_add_0_root_add_223_n148), .ZN(
        DP_add_0_root_add_0_root_add_223_n146) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U337 ( .A1(DP_ff_2_), .A2(
        DP_ff_part_2_), .ZN(DP_add_0_root_add_0_root_add_223_n157) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U336 ( .A1(
        DP_add_0_root_add_0_root_add_223_n157), .A2(
        DP_add_0_root_add_0_root_add_223_n155), .ZN(
        DP_add_0_root_add_0_root_add_223_n153) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U335 ( .A1(DP_ff_21_), .A2(
        DP_ff_part_21_), .ZN(DP_add_0_root_add_0_root_add_223_n36) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U334 ( .A1(DP_ff_19_), .A2(
        DP_ff_part_19_), .ZN(DP_add_0_root_add_0_root_add_223_n54) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U333 ( .A1(DP_ff_15_), .A2(
        DP_ff_part_15_), .ZN(DP_add_0_root_add_0_root_add_223_n84) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U332 ( .A1(DP_ff_13_), .A2(
        DP_ff_part_13_), .ZN(DP_add_0_root_add_0_root_add_223_n104) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U331 ( .A1(DP_ff_22_), .A2(
        DP_ff_part_22_), .ZN(DP_add_0_root_add_0_root_add_223_n27) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U330 ( .A1(DP_ff_10_), .A2(
        DP_ff_part_10_), .ZN(DP_add_0_root_add_0_root_add_223_n128) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U329 ( .A1(DP_ff_2_), .A2(
        DP_ff_part_2_), .ZN(DP_add_0_root_add_0_root_add_223_n158) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U328 ( .A1(DP_ff_3_), .A2(
        DP_ff_part_3_), .ZN(DP_add_0_root_add_0_root_add_223_n156) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U327 ( .B1(
        DP_add_0_root_add_0_root_add_223_n155), .B2(
        DP_add_0_root_add_0_root_add_223_n158), .A(
        DP_add_0_root_add_0_root_add_223_n156), .ZN(
        DP_add_0_root_add_0_root_add_223_n154) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U326 ( .A1(DP_ff_7_), .A2(
        DP_ff_part_7_), .ZN(DP_add_0_root_add_0_root_add_223_n143) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U325 ( .A1(DP_ff_6_), .A2(
        DP_ff_part_6_), .ZN(DP_add_0_root_add_0_root_add_223_n145) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U324 ( .B1(
        DP_add_0_root_add_0_root_add_223_n142), .B2(
        DP_add_0_root_add_0_root_add_223_n145), .A(
        DP_add_0_root_add_0_root_add_223_n143), .ZN(
        DP_add_0_root_add_0_root_add_223_n141) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U323 ( .A1(DP_ff_16_), .A2(
        DP_ff_part_16_), .ZN(DP_add_0_root_add_0_root_add_223_n75) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U322 ( .A1(DP_ff_14_), .A2(
        DP_ff_part_14_), .ZN(DP_add_0_root_add_0_root_add_223_n93) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U321 ( .A1(DP_ff_20_), .A2(
        DP_ff_part_20_), .ZN(DP_add_0_root_add_0_root_add_223_n43) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U320 ( .A1(DP_ff_18_), .A2(
        DP_ff_part_18_), .ZN(DP_add_0_root_add_0_root_add_223_n61) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U319 ( .A1(DP_ff_12_), .A2(
        DP_ff_part_12_), .ZN(DP_add_0_root_add_0_root_add_223_n111) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U318 ( .A1(DP_ff_5_), .A2(
        DP_ff_part_5_), .ZN(DP_add_0_root_add_0_root_add_223_n149) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U317 ( .A1(DP_ff_4_), .A2(
        DP_ff_part_4_), .ZN(DP_add_0_root_add_0_root_add_223_n151) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U316 ( .B1(
        DP_add_0_root_add_0_root_add_223_n148), .B2(
        DP_add_0_root_add_0_root_add_223_n151), .A(
        DP_add_0_root_add_0_root_add_223_n149), .ZN(
        DP_add_0_root_add_0_root_add_223_n147) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U315 ( .A1(DP_ff_11_), .A2(
        DP_ff_part_11_), .ZN(DP_add_0_root_add_0_root_add_223_n121) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U314 ( .A1(DP_ff_8_), .A2(
        DP_ff_part_8_), .ZN(DP_add_0_root_add_0_root_add_223_n134) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U313 ( .A1(
        DP_add_0_root_add_0_root_add_223_n134), .A2(
        DP_add_0_root_add_0_root_add_223_n132), .ZN(
        DP_add_0_root_add_0_root_add_223_n130) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U312 ( .A1(DP_ff_6_), .A2(
        DP_ff_part_6_), .ZN(DP_add_0_root_add_0_root_add_223_n144) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U311 ( .A1(
        DP_add_0_root_add_0_root_add_223_n144), .A2(
        DP_add_0_root_add_0_root_add_223_n142), .ZN(
        DP_add_0_root_add_0_root_add_223_n140) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U310 ( .A1(DP_ff_5_), .A2(
        DP_ff_part_5_), .ZN(DP_add_0_root_add_0_root_add_223_n148) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U309 ( .A1(DP_ff_3_), .A2(
        DP_ff_part_3_), .ZN(DP_add_0_root_add_0_root_add_223_n155) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U308 ( .A1(DP_ff_7_), .A2(
        DP_ff_part_7_), .ZN(DP_add_0_root_add_0_root_add_223_n142) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U307 ( .A1(DP_ff_9_), .A2(
        DP_ff_part_9_), .ZN(DP_add_0_root_add_0_root_add_223_n132) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U306 ( .A1(
        DP_add_0_root_add_0_root_add_223_n146), .A2(
        DP_add_0_root_add_0_root_add_223_n140), .ZN(
        DP_add_0_root_add_0_root_add_223_n138) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U305 ( .B1(
        DP_add_0_root_add_0_root_add_223_n140), .B2(
        DP_add_0_root_add_0_root_add_223_n147), .A(
        DP_add_0_root_add_0_root_add_223_n141), .ZN(
        DP_add_0_root_add_0_root_add_223_n139) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U304 ( .B1(
        DP_add_0_root_add_0_root_add_223_n153), .B2(
        DP_add_0_root_add_0_root_add_223_n159), .A(
        DP_add_0_root_add_0_root_add_223_n154), .ZN(
        DP_add_0_root_add_0_root_add_223_n152) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U303 ( .B1(
        DP_add_0_root_add_0_root_add_223_n152), .B2(
        DP_add_0_root_add_0_root_add_223_n138), .A(
        DP_add_0_root_add_0_root_add_223_n139), .ZN(
        DP_add_0_root_add_0_root_add_223_n137) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U302 ( .A1(DP_ff_9_), .A2(
        DP_ff_part_9_), .ZN(DP_add_0_root_add_0_root_add_223_n133) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U301 ( .A1(DP_ff_8_), .A2(
        DP_ff_part_8_), .ZN(DP_add_0_root_add_0_root_add_223_n135) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U300 ( .B1(
        DP_add_0_root_add_0_root_add_223_n132), .B2(
        DP_add_0_root_add_0_root_add_223_n135), .A(
        DP_add_0_root_add_0_root_add_223_n133), .ZN(
        DP_add_0_root_add_0_root_add_223_n131) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U299 ( .A1(DP_ff_17_), .A2(
        DP_ff_part_17_), .ZN(DP_add_0_root_add_0_root_add_223_n71) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U298 ( .A(
        DP_add_0_root_add_0_root_add_223_n129), .ZN(
        DP_add_0_root_add_0_root_add_223_n127) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U297 ( .A(
        DP_add_0_root_add_0_root_add_223_n111), .ZN(
        DP_add_0_root_add_0_root_add_223_n109) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U296 ( .A(
        DP_add_0_root_add_0_root_add_223_n61), .ZN(
        DP_add_0_root_add_0_root_add_223_n59) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U295 ( .A(
        DP_add_0_root_add_0_root_add_223_n43), .ZN(
        DP_add_0_root_add_0_root_add_223_n41) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U294 ( .A(
        DP_add_0_root_add_0_root_add_223_n121), .ZN(
        DP_add_0_root_add_0_root_add_223_n175) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U293 ( .A1(
        DP_add_0_root_add_0_root_add_223_n175), .A2(
        DP_add_0_root_add_0_root_add_223_n122), .ZN(
        DP_add_0_root_add_0_root_add_223_n14) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U292 ( .A(
        DP_add_0_root_add_0_root_add_223_n83), .ZN(
        DP_add_0_root_add_0_root_add_223_n171) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U291 ( .A1(
        DP_add_0_root_add_0_root_add_223_n171), .A2(
        DP_add_0_root_add_0_root_add_223_n84), .ZN(
        DP_add_0_root_add_0_root_add_223_n10) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U290 ( .A(
        DP_add_0_root_add_0_root_add_223_n103), .ZN(
        DP_add_0_root_add_0_root_add_223_n173) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U289 ( .A1(
        DP_add_0_root_add_0_root_add_223_n173), .A2(
        DP_add_0_root_add_0_root_add_223_n104), .ZN(
        DP_add_0_root_add_0_root_add_223_n12) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U288 ( .A(
        DP_add_0_root_add_0_root_add_223_n74), .ZN(
        DP_add_0_root_add_0_root_add_223_n170) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U287 ( .A1(
        DP_add_0_root_add_0_root_add_223_n170), .A2(
        DP_add_0_root_add_0_root_add_223_n75), .ZN(
        DP_add_0_root_add_0_root_add_223_n9) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U286 ( .A1(
        DP_add_0_root_add_0_root_add_223_n91), .A2(
        DP_add_0_root_add_0_root_add_223_n93), .ZN(
        DP_add_0_root_add_0_root_add_223_n11) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U285 ( .A1(
        DP_add_0_root_add_0_root_add_223_n108), .A2(
        DP_add_0_root_add_0_root_add_223_n111), .ZN(
        DP_add_0_root_add_0_root_add_223_n13) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U284 ( .A1(
        DP_add_0_root_add_0_root_add_223_n58), .A2(
        DP_add_0_root_add_0_root_add_223_n61), .ZN(
        DP_add_0_root_add_0_root_add_223_n7) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U283 ( .A(
        DP_add_0_root_add_0_root_add_223_n42), .ZN(
        DP_add_0_root_add_0_root_add_223_n166) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U282 ( .A1(
        DP_add_0_root_add_0_root_add_223_n166), .A2(
        DP_add_0_root_add_0_root_add_223_n43), .ZN(
        DP_add_0_root_add_0_root_add_223_n5) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U281 ( .A(
        DP_add_0_root_add_0_root_add_223_n35), .ZN(
        DP_add_0_root_add_0_root_add_223_n165) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U280 ( .A1(
        DP_add_0_root_add_0_root_add_223_n165), .A2(
        DP_add_0_root_add_0_root_add_223_n36), .ZN(
        DP_add_0_root_add_0_root_add_223_n4) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U279 ( .A(
        DP_add_0_root_add_0_root_add_223_n53), .ZN(
        DP_add_0_root_add_0_root_add_223_n167) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U278 ( .A1(
        DP_add_0_root_add_0_root_add_223_n167), .A2(
        DP_add_0_root_add_0_root_add_223_n54), .ZN(
        DP_add_0_root_add_0_root_add_223_n6) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U277 ( .A(
        DP_add_0_root_add_0_root_add_223_n27), .ZN(
        DP_add_0_root_add_0_root_add_223_n25) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U276 ( .B1(
        DP_add_0_root_add_0_root_add_223_n34), .B2(
        DP_add_0_root_add_0_root_add_223_n243), .A(
        DP_add_0_root_add_0_root_add_223_n25), .ZN(
        DP_add_0_root_add_0_root_add_223_n23) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U275 ( .A(
        DP_add_0_root_add_0_root_add_223_n21), .ZN(
        DP_add_0_root_add_0_root_add_223_n19) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U274 ( .A(
        DP_add_0_root_add_0_root_add_223_n92), .ZN(
        DP_add_0_root_add_0_root_add_223_n91) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U273 ( .A(
        DP_add_0_root_add_0_root_add_223_n91), .ZN(
        DP_add_0_root_add_0_root_add_223_n90) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U272 ( .B1(
        DP_add_0_root_add_0_root_add_223_n53), .B2(
        DP_add_0_root_add_0_root_add_223_n61), .A(
        DP_add_0_root_add_0_root_add_223_n54), .ZN(
        DP_add_0_root_add_0_root_add_223_n52) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U271 ( .B1(
        DP_add_0_root_add_0_root_add_223_n51), .B2(
        DP_add_0_root_add_0_root_add_223_n70), .A(
        DP_add_0_root_add_0_root_add_223_n52), .ZN(
        DP_add_0_root_add_0_root_add_223_n50) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U270 ( .A(
        DP_add_0_root_add_0_root_add_223_n128), .ZN(
        DP_add_0_root_add_0_root_add_223_n126) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U269 ( .B1(
        DP_add_0_root_add_0_root_add_223_n131), .B2(
        DP_add_0_root_add_0_root_add_223_n126), .A(
        DP_add_0_root_add_0_root_add_223_n127), .ZN(
        DP_add_0_root_add_0_root_add_223_n125) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U268 ( .A1(
        DP_add_0_root_add_0_root_add_223_n130), .A2(
        DP_add_0_root_add_0_root_add_223_n126), .ZN(
        DP_add_0_root_add_0_root_add_223_n124) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U267 ( .B1(
        DP_add_0_root_add_0_root_add_223_n136), .B2(
        DP_add_0_root_add_0_root_add_223_n124), .A(
        DP_add_0_root_add_0_root_add_223_n125), .ZN(
        DP_add_0_root_add_0_root_add_223_n123) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U266 ( .A(
        DP_add_0_root_add_0_root_add_223_n110), .ZN(
        DP_add_0_root_add_0_root_add_223_n108) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U265 ( .B1(
        DP_add_0_root_add_0_root_add_223_n116), .B2(
        DP_add_0_root_add_0_root_add_223_n108), .A(
        DP_add_0_root_add_0_root_add_223_n109), .ZN(
        DP_add_0_root_add_0_root_add_223_n107) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U264 ( .A1(
        DP_add_0_root_add_0_root_add_223_n115), .A2(
        DP_add_0_root_add_0_root_add_223_n108), .ZN(
        DP_add_0_root_add_0_root_add_223_n106) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U263 ( .B1(
        DP_add_0_root_add_0_root_add_223_n136), .B2(
        DP_add_0_root_add_0_root_add_223_n106), .A(
        DP_add_0_root_add_0_root_add_223_n107), .ZN(
        DP_add_0_root_add_0_root_add_223_n105) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U262 ( .A(
        DP_add_0_root_add_0_root_add_223_n60), .ZN(
        DP_add_0_root_add_0_root_add_223_n58) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U261 ( .B1(
        DP_add_0_root_add_0_root_add_223_n66), .B2(
        DP_add_0_root_add_0_root_add_223_n58), .A(
        DP_add_0_root_add_0_root_add_223_n59), .ZN(
        DP_add_0_root_add_0_root_add_223_n57) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U260 ( .A1(
        DP_add_0_root_add_0_root_add_223_n69), .A2(
        DP_add_0_root_add_0_root_add_223_n58), .ZN(
        DP_add_0_root_add_0_root_add_223_n56) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U259 ( .B1(
        DP_add_0_root_add_0_root_add_223_n1), .B2(
        DP_add_0_root_add_0_root_add_223_n56), .A(
        DP_add_0_root_add_0_root_add_223_n57), .ZN(
        DP_add_0_root_add_0_root_add_223_n55) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U258 ( .B1(
        DP_add_0_root_add_0_root_add_223_n48), .B2(
        DP_add_0_root_add_0_root_add_223_n166), .A(
        DP_add_0_root_add_0_root_add_223_n41), .ZN(
        DP_add_0_root_add_0_root_add_223_n39) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U257 ( .A1(
        DP_add_0_root_add_0_root_add_223_n47), .A2(
        DP_add_0_root_add_0_root_add_223_n166), .ZN(
        DP_add_0_root_add_0_root_add_223_n38) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U256 ( .B1(
        DP_add_0_root_add_0_root_add_223_n1), .B2(
        DP_add_0_root_add_0_root_add_223_n38), .A(
        DP_add_0_root_add_0_root_add_223_n39), .ZN(
        DP_add_0_root_add_0_root_add_223_n37) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U255 ( .B1(
        DP_add_0_root_add_0_root_add_223_n1), .B2(
        DP_add_0_root_add_0_root_add_223_n74), .A(
        DP_add_0_root_add_0_root_add_223_n75), .ZN(
        DP_add_0_root_add_0_root_add_223_n73) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U254 ( .A1(
        DP_add_0_root_add_0_root_add_223_n130), .A2(
        DP_add_0_root_add_0_root_add_223_n119), .ZN(
        DP_add_0_root_add_0_root_add_223_n117) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U253 ( .A1(
        DP_add_0_root_add_0_root_add_223_n169), .A2(
        DP_add_0_root_add_0_root_add_223_n72), .ZN(
        DP_add_0_root_add_0_root_add_223_n8) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U252 ( .B1(
        DP_add_0_root_add_0_root_add_223_n100), .B2(
        DP_add_0_root_add_0_root_add_223_n90), .A(
        DP_add_0_root_add_0_root_add_223_n93), .ZN(
        DP_add_0_root_add_0_root_add_223_n89) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U251 ( .A1(
        DP_add_0_root_add_0_root_add_223_n60), .A2(
        DP_add_0_root_add_0_root_add_223_n53), .ZN(
        DP_add_0_root_add_0_root_add_223_n51) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U250 ( .B1(
        DP_add_0_root_add_0_root_add_223_n83), .B2(
        DP_add_0_root_add_0_root_add_223_n93), .A(
        DP_add_0_root_add_0_root_add_223_n84), .ZN(
        DP_add_0_root_add_0_root_add_223_n82) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U249 ( .B1(
        DP_add_0_root_add_0_root_add_223_n81), .B2(
        DP_add_0_root_add_0_root_add_223_n102), .A(
        DP_add_0_root_add_0_root_add_223_n82), .ZN(
        DP_add_0_root_add_0_root_add_223_n80) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U248 ( .A(
        DP_add_0_root_add_0_root_add_223_n137), .ZN(
        DP_add_0_root_add_0_root_add_223_n136) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U247 ( .A1(
        DP_add_0_root_add_0_root_add_223_n243), .A2(
        DP_add_0_root_add_0_root_add_223_n27), .ZN(
        DP_add_0_root_add_0_root_add_223_n3) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U246 ( .A1(
        DP_add_0_root_add_0_root_add_223_n110), .A2(
        DP_add_0_root_add_0_root_add_223_n103), .ZN(
        DP_add_0_root_add_0_root_add_223_n101) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U245 ( .A1(
        DP_add_0_root_add_0_root_add_223_n42), .A2(
        DP_add_0_root_add_0_root_add_223_n35), .ZN(
        DP_add_0_root_add_0_root_add_223_n33) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U244 ( .A1(
        DP_add_0_root_add_0_root_add_223_n92), .A2(
        DP_add_0_root_add_0_root_add_223_n83), .ZN(
        DP_add_0_root_add_0_root_add_223_n81) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U243 ( .B1(
        DP_add_0_root_add_0_root_add_223_n35), .B2(
        DP_add_0_root_add_0_root_add_223_n43), .A(
        DP_add_0_root_add_0_root_add_223_n36), .ZN(
        DP_add_0_root_add_0_root_add_223_n34) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U242 ( .B1(
        DP_add_0_root_add_0_root_add_223_n103), .B2(
        DP_add_0_root_add_0_root_add_223_n111), .A(
        DP_add_0_root_add_0_root_add_223_n104), .ZN(
        DP_add_0_root_add_0_root_add_223_n102) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U241 ( .B1(
        DP_add_0_root_add_0_root_add_223_n119), .B2(
        DP_add_0_root_add_0_root_add_223_n131), .A(
        DP_add_0_root_add_0_root_add_223_n120), .ZN(
        DP_add_0_root_add_0_root_add_223_n118) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U240 ( .B1(
        DP_add_0_root_add_0_root_add_223_n118), .B2(
        DP_add_0_root_add_0_root_add_223_n79), .A(
        DP_add_0_root_add_0_root_add_223_n80), .ZN(
        DP_add_0_root_add_0_root_add_223_n78) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U239 ( .A1(
        DP_add_0_root_add_0_root_add_223_n117), .A2(
        DP_add_0_root_add_0_root_add_223_n79), .ZN(
        DP_add_0_root_add_0_root_add_223_n77) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U238 ( .B1(
        DP_add_0_root_add_0_root_add_223_n137), .B2(
        DP_add_0_root_add_0_root_add_223_n77), .A(
        DP_add_0_root_add_0_root_add_223_n78), .ZN(
        DP_add_0_root_add_0_root_add_223_n76) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U237 ( .B1(
        DP_add_0_root_add_0_root_add_223_n71), .B2(
        DP_add_0_root_add_0_root_add_223_n75), .A(
        DP_add_0_root_add_0_root_add_223_n72), .ZN(
        DP_add_0_root_add_0_root_add_223_n70) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U236 ( .A1(
        DP_add_0_root_add_0_root_add_223_n74), .A2(
        DP_add_0_root_add_0_root_add_223_n71), .ZN(
        DP_add_0_root_add_0_root_add_223_n69) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U235 ( .A(
        DP_add_0_root_add_0_root_add_223_n116), .ZN(
        DP_add_0_root_add_0_root_add_223_n114) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U234 ( .A(
        DP_add_0_root_add_0_root_add_223_n115), .ZN(
        DP_add_0_root_add_0_root_add_223_n113) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U233 ( .B1(
        DP_add_0_root_add_0_root_add_223_n136), .B2(
        DP_add_0_root_add_0_root_add_223_n113), .A(
        DP_add_0_root_add_0_root_add_223_n114), .ZN(
        DP_add_0_root_add_0_root_add_223_n112) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U232 ( .A(
        DP_add_0_root_add_0_root_add_223_n33), .ZN(
        DP_add_0_root_add_0_root_add_223_n32) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U231 ( .A(
        DP_add_0_root_add_0_root_add_223_n32), .ZN(
        DP_add_0_root_add_0_root_add_223_n31) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U230 ( .A(
        DP_add_0_root_add_0_root_add_223_n70), .ZN(
        DP_add_0_root_add_0_root_add_223_n68) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U229 ( .A(
        DP_add_0_root_add_0_root_add_223_n68), .ZN(
        DP_add_0_root_add_0_root_add_223_n66) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U228 ( .A1(
        DP_add_0_root_add_0_root_add_223_n33), .A2(
        DP_add_0_root_add_0_root_add_223_n243), .ZN(
        DP_add_0_root_add_0_root_add_223_n22) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U227 ( .A(
        DP_add_0_root_add_0_root_add_223_n101), .ZN(
        DP_add_0_root_add_0_root_add_223_n99) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U226 ( .A(
        DP_add_0_root_add_0_root_add_223_n102), .ZN(
        DP_add_0_root_add_0_root_add_223_n100) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U225 ( .A1(
        DP_add_0_root_add_0_root_add_223_n101), .A2(
        DP_add_0_root_add_0_root_add_223_n81), .ZN(
        DP_add_0_root_add_0_root_add_223_n79) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U224 ( .A1(
        DP_add_0_root_add_0_root_add_223_n69), .A2(
        DP_add_0_root_add_0_root_add_223_n51), .ZN(
        DP_add_0_root_add_0_root_add_223_n49) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U223 ( .A(
        DP_add_0_root_add_0_root_add_223_n99), .ZN(
        DP_add_0_root_add_0_root_add_223_n97) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U222 ( .B1(
        DP_add_0_root_add_0_root_add_223_n116), .B2(
        DP_add_0_root_add_0_root_add_223_n97), .A(
        DP_add_0_root_add_0_root_add_223_n98), .ZN(
        DP_add_0_root_add_0_root_add_223_n96) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U221 ( .A1(
        DP_add_0_root_add_0_root_add_223_n115), .A2(
        DP_add_0_root_add_0_root_add_223_n97), .ZN(
        DP_add_0_root_add_0_root_add_223_n95) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U220 ( .B1(
        DP_add_0_root_add_0_root_add_223_n136), .B2(
        DP_add_0_root_add_0_root_add_223_n95), .A(
        DP_add_0_root_add_0_root_add_223_n96), .ZN(
        DP_add_0_root_add_0_root_add_223_n94) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U219 ( .A1(
        DP_add_0_root_add_0_root_add_223_n99), .A2(
        DP_add_0_root_add_0_root_add_223_n90), .ZN(
        DP_add_0_root_add_0_root_add_223_n88) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U218 ( .B1(
        DP_add_0_root_add_0_root_add_223_n88), .B2(
        DP_add_0_root_add_0_root_add_223_n116), .A(
        DP_add_0_root_add_0_root_add_223_n89), .ZN(
        DP_add_0_root_add_0_root_add_223_n87) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U217 ( .A1(
        DP_add_0_root_add_0_root_add_223_n88), .A2(
        DP_add_0_root_add_0_root_add_223_n115), .ZN(
        DP_add_0_root_add_0_root_add_223_n86) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U216 ( .B1(
        DP_add_0_root_add_0_root_add_223_n136), .B2(
        DP_add_0_root_add_0_root_add_223_n86), .A(
        DP_add_0_root_add_0_root_add_223_n87), .ZN(
        DP_add_0_root_add_0_root_add_223_n85) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U215 ( .A(
        DP_add_0_root_add_0_root_add_223_n66), .ZN(
        DP_add_0_root_add_0_root_add_223_n64) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U214 ( .A(
        DP_add_0_root_add_0_root_add_223_n69), .ZN(
        DP_add_0_root_add_0_root_add_223_n63) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U213 ( .B1(
        DP_add_0_root_add_0_root_add_223_n1), .B2(
        DP_add_0_root_add_0_root_add_223_n63), .A(
        DP_add_0_root_add_0_root_add_223_n64), .ZN(
        DP_add_0_root_add_0_root_add_223_n62) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U212 ( .A(
        DP_add_0_root_add_0_root_add_223_n47), .ZN(
        DP_add_0_root_add_0_root_add_223_n45) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U211 ( .A(
        DP_add_0_root_add_0_root_add_223_n48), .ZN(
        DP_add_0_root_add_0_root_add_223_n46) );
  OAI21_X1 DP_add_0_root_add_0_root_add_223_U210 ( .B1(
        DP_add_0_root_add_0_root_add_223_n1), .B2(
        DP_add_0_root_add_0_root_add_223_n45), .A(
        DP_add_0_root_add_0_root_add_223_n46), .ZN(
        DP_add_0_root_add_0_root_add_223_n44) );
  AOI21_X1 DP_add_0_root_add_0_root_add_223_U209 ( .B1(
        DP_add_0_root_add_0_root_add_223_n48), .B2(
        DP_add_0_root_add_0_root_add_223_n31), .A(
        DP_add_0_root_add_0_root_add_223_n34), .ZN(
        DP_add_0_root_add_0_root_add_223_n30) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U208 ( .A(
        DP_add_0_root_add_0_root_add_223_n117), .ZN(
        DP_add_0_root_add_0_root_add_223_n115) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U207 ( .A(
        DP_add_0_root_add_0_root_add_223_n118), .ZN(
        DP_add_0_root_add_0_root_add_223_n116) );
  NAND2_X1 DP_add_0_root_add_0_root_add_223_U206 ( .A1(
        DP_add_0_root_add_0_root_add_223_n47), .A2(
        DP_add_0_root_add_0_root_add_223_n31), .ZN(
        DP_add_0_root_add_0_root_add_223_n29) );
  OR2_X1 DP_add_0_root_add_0_root_add_223_U205 ( .A1(
        DP_add_0_root_add_0_root_add_223_n49), .A2(
        DP_add_0_root_add_0_root_add_223_n22), .ZN(
        DP_add_0_root_add_0_root_add_223_n244) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U204 ( .A(
        DP_add_0_root_add_0_root_add_223_n100), .ZN(
        DP_add_0_root_add_0_root_add_223_n98) );
  INV_X1 DP_add_0_root_add_0_root_add_223_U203 ( .A(
        DP_add_0_root_add_0_root_add_223_n49), .ZN(
        DP_add_0_root_add_0_root_add_223_n47) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U202 ( .A1(DP_ff_21_), .A2(
        DP_ff_part_21_), .ZN(DP_add_0_root_add_0_root_add_223_n35) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U201 ( .A1(DP_ff_13_), .A2(
        DP_ff_part_13_), .ZN(DP_add_0_root_add_0_root_add_223_n103) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U200 ( .A1(DP_ff_15_), .A2(
        DP_ff_part_15_), .ZN(DP_add_0_root_add_0_root_add_223_n83) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U199 ( .A1(DP_ff_19_), .A2(
        DP_ff_part_19_), .ZN(DP_add_0_root_add_0_root_add_223_n53) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U198 ( .A1(DP_ff_20_), .A2(
        DP_ff_part_20_), .ZN(DP_add_0_root_add_0_root_add_223_n42) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U197 ( .A1(DP_ff_18_), .A2(
        DP_ff_part_18_), .ZN(DP_add_0_root_add_0_root_add_223_n60) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U196 ( .A1(DP_ff_12_), .A2(
        DP_ff_part_12_), .ZN(DP_add_0_root_add_0_root_add_223_n110) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U195 ( .A1(DP_ff_14_), .A2(
        DP_ff_part_14_), .ZN(DP_add_0_root_add_0_root_add_223_n92) );
  NOR2_X1 DP_add_0_root_add_0_root_add_223_U194 ( .A1(DP_ff_16_), .A2(
        DP_ff_part_16_), .ZN(DP_add_0_root_add_0_root_add_223_n74) );
  CLKBUF_X3 DP_add_0_root_add_0_root_add_223_U193 ( .A(
        DP_add_0_root_add_0_root_add_223_n76), .Z(
        DP_add_0_root_add_0_root_add_223_n1) );
  OR2_X1 DP_add_0_root_add_0_root_add_223_U192 ( .A1(DP_ff_22_), .A2(
        DP_ff_part_22_), .ZN(DP_add_0_root_add_0_root_add_223_n243) );
  INV_X1 DP_mult_205_U2828 ( .A(DP_mult_205_n2325), .ZN(DP_mult_205_n2324) );
  INV_X1 DP_mult_205_U2827 ( .A(DP_mult_205_n2317), .ZN(DP_mult_205_n2316) );
  INV_X1 DP_mult_205_U2826 ( .A(DP_mult_205_n2044), .ZN(DP_mult_205_n2300) );
  INV_X1 DP_mult_205_U2825 ( .A(DP_mult_205_n2164), .ZN(DP_mult_205_n2296) );
  INV_X1 DP_mult_205_U2824 ( .A(DP_mult_205_n2286), .ZN(DP_mult_205_n2285) );
  INV_X1 DP_mult_205_U2823 ( .A(DP_mult_205_n2134), .ZN(DP_mult_205_n2279) );
  INV_X1 DP_mult_205_U2822 ( .A(DP_mult_205_n1992), .ZN(DP_mult_205_n2263) );
  INV_X1 DP_mult_205_U2821 ( .A(DP_mult_205_n1986), .ZN(DP_mult_205_n2260) );
  INV_X1 DP_mult_205_U2820 ( .A(DP_mult_205_n2204), .ZN(DP_mult_205_n2257) );
  XNOR2_X1 DP_mult_205_U2819 ( .A(DP_sw1_17_), .B(DP_mult_205_n2292), .ZN(
        DP_mult_205_n1713) );
  XNOR2_X1 DP_mult_205_U2818 ( .A(DP_sw1_19_), .B(DP_mult_205_n2290), .ZN(
        DP_mult_205_n1711) );
  XNOR2_X1 DP_mult_205_U2817 ( .A(DP_sw1_11_), .B(DP_mult_205_n2292), .ZN(
        DP_mult_205_n1719) );
  XNOR2_X1 DP_mult_205_U2816 ( .A(DP_sw1_15_), .B(DP_mult_205_n2291), .ZN(
        DP_mult_205_n1715) );
  XNOR2_X1 DP_mult_205_U2815 ( .A(DP_sw1_21_), .B(DP_mult_205_n2291), .ZN(
        DP_mult_205_n1709) );
  OAI22_X1 DP_mult_205_U2814 ( .A1(DP_mult_205_n2247), .A2(DP_mult_205_n1683), 
        .B1(DP_mult_205_n1682), .B2(DP_mult_205_n1983), .ZN(DP_mult_205_n836)
         );
  XNOR2_X1 DP_mult_205_U2813 ( .A(DP_sw1_13_), .B(DP_mult_205_n2291), .ZN(
        DP_mult_205_n1717) );
  OAI22_X1 DP_mult_205_U2812 ( .A1(DP_mult_205_n1706), .A2(DP_mult_205_n1983), 
        .B1(DP_mult_205_n2171), .B2(DP_mult_205_n2164), .ZN(DP_mult_205_n1190)
         );
  OAI22_X1 DP_mult_205_U2811 ( .A1(DP_mult_205_n2096), .A2(DP_mult_205_n1693), 
        .B1(DP_mult_205_n1692), .B2(DP_mult_205_n1983), .ZN(DP_mult_205_n1396)
         );
  OAI22_X1 DP_mult_205_U2810 ( .A1(DP_mult_205_n2248), .A2(DP_mult_205_n1684), 
        .B1(DP_mult_205_n1982), .B2(DP_mult_205_n1683), .ZN(DP_mult_205_n1387)
         );
  INV_X1 DP_mult_205_U2809 ( .A(DP_mult_205_n836), .ZN(DP_mult_205_n837) );
  OAI22_X1 DP_mult_205_U2808 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1688), 
        .B1(DP_mult_205_n1983), .B2(DP_mult_205_n1687), .ZN(DP_mult_205_n1391)
         );
  OAI22_X1 DP_mult_205_U2807 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1685), 
        .B1(DP_mult_205_n1684), .B2(DP_mult_205_n1982), .ZN(DP_mult_205_n1388)
         );
  OAI22_X1 DP_mult_205_U2806 ( .A1(DP_mult_205_n2095), .A2(DP_mult_205_n1692), 
        .B1(DP_mult_205_n1982), .B2(DP_mult_205_n1691), .ZN(DP_mult_205_n1395)
         );
  OAI22_X1 DP_mult_205_U2805 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1687), 
        .B1(DP_mult_205_n1686), .B2(DP_mult_205_n1982), .ZN(DP_mult_205_n1390)
         );
  OAI22_X1 DP_mult_205_U2804 ( .A1(DP_mult_205_n2096), .A2(DP_mult_205_n1690), 
        .B1(DP_mult_205_n1982), .B2(DP_mult_205_n1689), .ZN(DP_mult_205_n1393)
         );
  OAI22_X1 DP_mult_205_U2803 ( .A1(DP_mult_205_n2095), .A2(DP_mult_205_n1689), 
        .B1(DP_mult_205_n1688), .B2(DP_mult_205_n1983), .ZN(DP_mult_205_n1392)
         );
  OAI22_X1 DP_mult_205_U2802 ( .A1(DP_mult_205_n2248), .A2(DP_mult_205_n1686), 
        .B1(DP_mult_205_n1983), .B2(DP_mult_205_n1685), .ZN(DP_mult_205_n1389)
         );
  OAI22_X1 DP_mult_205_U2801 ( .A1(DP_mult_205_n2096), .A2(DP_mult_205_n1691), 
        .B1(DP_mult_205_n1690), .B2(DP_mult_205_n1982), .ZN(DP_mult_205_n1394)
         );
  NAND2_X1 DP_mult_205_U2800 ( .A1(DP_mult_205_n775), .A2(DP_mult_205_n788), 
        .ZN(DP_mult_205_n474) );
  OAI21_X1 DP_mult_205_U2799 ( .B1(DP_mult_205_n301), .B2(DP_mult_205_n398), 
        .A(DP_mult_205_n399), .ZN(DP_mult_205_n397) );
  OAI21_X1 DP_mult_205_U2798 ( .B1(DP_mult_205_n2230), .B2(DP_mult_205_n389), 
        .A(DP_mult_205_n390), .ZN(DP_mult_205_n388) );
  OAI21_X1 DP_mult_205_U2797 ( .B1(DP_mult_205_n301), .B2(DP_mult_205_n431), 
        .A(DP_mult_205_n432), .ZN(DP_mult_205_n430) );
  OAI21_X1 DP_mult_205_U2796 ( .B1(DP_mult_205_n2230), .B2(DP_mult_205_n411), 
        .A(DP_mult_205_n412), .ZN(DP_mult_205_n410) );
  OAI21_X1 DP_mult_205_U2795 ( .B1(DP_mult_205_n2230), .B2(DP_mult_205_n420), 
        .A(DP_mult_205_n421), .ZN(DP_mult_205_n419) );
  OAI21_X1 DP_mult_205_U2794 ( .B1(DP_mult_205_n301), .B2(DP_mult_205_n343), 
        .A(DP_mult_205_n344), .ZN(DP_mult_205_n342) );
  OAI21_X1 DP_mult_205_U2793 ( .B1(DP_mult_205_n301), .B2(DP_mult_205_n380), 
        .A(DP_mult_205_n381), .ZN(DP_mult_205_n379) );
  OAI21_X1 DP_mult_205_U2792 ( .B1(DP_mult_205_n301), .B2(DP_mult_205_n371), 
        .A(DP_mult_205_n372), .ZN(DP_mult_205_n370) );
  OAI21_X1 DP_mult_205_U2791 ( .B1(DP_mult_205_n301), .B2(DP_mult_205_n354), 
        .A(DP_mult_205_n355), .ZN(DP_mult_205_n353) );
  OAI21_X1 DP_mult_205_U2790 ( .B1(DP_mult_205_n2230), .B2(DP_mult_205_n438), 
        .A(DP_mult_205_n439), .ZN(DP_mult_205_n437) );
  INV_X1 DP_mult_205_U2789 ( .A(DP_mult_205_n2230), .ZN(DP_mult_205_n448) );
  OAI21_X1 DP_mult_205_U2788 ( .B1(DP_mult_205_n2230), .B2(DP_mult_205_n326), 
        .A(DP_mult_205_n327), .ZN(DP_mult_205_n325) );
  XNOR2_X1 DP_mult_205_U2787 ( .A(DP_mult_205_n437), .B(DP_mult_205_n311), 
        .ZN(DP_sw1_coeff_ret1[13]) );
  NAND2_X1 DP_mult_205_U2786 ( .A1(DP_mult_205_n1815), .A2(DP_mult_205_n2156), 
        .ZN(DP_mult_205_n279) );
  XNOR2_X1 DP_mult_205_U2785 ( .A(DP_sw1_13_), .B(DP_mult_205_n2288), .ZN(
        DP_mult_205_n1742) );
  XNOR2_X1 DP_mult_205_U2784 ( .A(DP_sw1_17_), .B(DP_mult_205_n2287), .ZN(
        DP_mult_205_n1738) );
  XNOR2_X1 DP_mult_205_U2783 ( .A(DP_sw1_11_), .B(DP_mult_205_n2288), .ZN(
        DP_mult_205_n1744) );
  XNOR2_X1 DP_mult_205_U2782 ( .A(DP_sw1_19_), .B(DP_mult_205_n2288), .ZN(
        DP_mult_205_n1736) );
  XNOR2_X1 DP_mult_205_U2781 ( .A(DP_sw1_15_), .B(DP_mult_205_n2287), .ZN(
        DP_mult_205_n1740) );
  XNOR2_X1 DP_mult_205_U2780 ( .A(DP_sw1_21_), .B(DP_mult_205_n2287), .ZN(
        DP_mult_205_n1734) );
  OAI22_X1 DP_mult_205_U2779 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1714), 
        .B1(DP_mult_205_n1713), .B2(DP_mult_205_n2043), .ZN(DP_mult_205_n1416)
         );
  OAI22_X1 DP_mult_205_U2778 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1719), 
        .B1(DP_mult_205_n2276), .B2(DP_mult_205_n1718), .ZN(DP_mult_205_n1421)
         );
  OAI22_X1 DP_mult_205_U2777 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1716), 
        .B1(DP_mult_205_n1715), .B2(DP_mult_205_n2042), .ZN(DP_mult_205_n1418)
         );
  OAI22_X1 DP_mult_205_U2776 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1712), 
        .B1(DP_mult_205_n1711), .B2(DP_mult_205_n2276), .ZN(DP_mult_205_n1414)
         );
  OAI22_X1 DP_mult_205_U2775 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1722), 
        .B1(DP_mult_205_n1721), .B2(DP_mult_205_n2042), .ZN(DP_mult_205_n1424)
         );
  OAI22_X1 DP_mult_205_U2774 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1729), 
        .B1(DP_mult_205_n2043), .B2(DP_mult_205_n1728), .ZN(DP_mult_205_n1431)
         );
  OAI22_X1 DP_mult_205_U2773 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1728), 
        .B1(DP_mult_205_n1727), .B2(DP_mult_205_n2043), .ZN(DP_mult_205_n1430)
         );
  OAI22_X1 DP_mult_205_U2772 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1710), 
        .B1(DP_mult_205_n1709), .B2(DP_mult_205_n2276), .ZN(DP_mult_205_n1412)
         );
  OAI22_X1 DP_mult_205_U2771 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1723), 
        .B1(DP_mult_205_n2276), .B2(DP_mult_205_n1722), .ZN(DP_mult_205_n1425)
         );
  OAI22_X1 DP_mult_205_U2770 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1725), 
        .B1(DP_mult_205_n2043), .B2(DP_mult_205_n1724), .ZN(DP_mult_205_n1427)
         );
  OAI22_X1 DP_mult_205_U2769 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1708), 
        .B1(DP_mult_205_n1707), .B2(DP_mult_205_n2276), .ZN(DP_mult_205_n874)
         );
  OAI22_X1 DP_mult_205_U2768 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1730), 
        .B1(DP_mult_205_n1729), .B2(DP_mult_205_n2042), .ZN(DP_mult_205_n1432)
         );
  OAI22_X1 DP_mult_205_U2767 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1726), 
        .B1(DP_mult_205_n1725), .B2(DP_mult_205_n2276), .ZN(DP_mult_205_n1428)
         );
  OAI22_X1 DP_mult_205_U2766 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1718), 
        .B1(DP_mult_205_n1717), .B2(DP_mult_205_n2042), .ZN(DP_mult_205_n1420)
         );
  OAI22_X1 DP_mult_205_U2765 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1721), 
        .B1(DP_mult_205_n2276), .B2(DP_mult_205_n1720), .ZN(DP_mult_205_n1423)
         );
  OAI22_X1 DP_mult_205_U2764 ( .A1(DP_mult_205_n1731), .A2(DP_mult_205_n2042), 
        .B1(DP_mult_205_n2249), .B2(DP_mult_205_n2106), .ZN(DP_mult_205_n1191)
         );
  OAI22_X1 DP_mult_205_U2763 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1720), 
        .B1(DP_mult_205_n1719), .B2(DP_mult_205_n2043), .ZN(DP_mult_205_n1422)
         );
  OAI22_X1 DP_mult_205_U2762 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1727), 
        .B1(DP_mult_205_n2043), .B2(DP_mult_205_n1726), .ZN(DP_mult_205_n1429)
         );
  OAI21_X1 DP_mult_205_U2761 ( .B1(DP_mult_205_n536), .B2(DP_mult_205_n498), 
        .A(DP_mult_205_n499), .ZN(DP_mult_205_n497) );
  OAI21_X1 DP_mult_205_U2760 ( .B1(DP_mult_205_n536), .B2(DP_mult_205_n487), 
        .A(DP_mult_205_n488), .ZN(DP_mult_205_n486) );
  OAI21_X1 DP_mult_205_U2759 ( .B1(DP_mult_205_n536), .B2(DP_mult_205_n476), 
        .A(DP_mult_205_n477), .ZN(DP_mult_205_n475) );
  OAI21_X1 DP_mult_205_U2758 ( .B1(DP_mult_205_n536), .B2(DP_mult_205_n2158), 
        .A(DP_mult_205_n524), .ZN(DP_mult_205_n522) );
  OAI21_X1 DP_mult_205_U2757 ( .B1(DP_mult_205_n536), .B2(DP_mult_205_n463), 
        .A(DP_mult_205_n464), .ZN(DP_mult_205_n462) );
  OAI21_X1 DP_mult_205_U2756 ( .B1(DP_mult_205_n536), .B2(DP_mult_205_n534), 
        .A(DP_mult_205_n2031), .ZN(DP_mult_205_n533) );
  OAI21_X1 DP_mult_205_U2755 ( .B1(DP_mult_205_n536), .B2(DP_mult_205_n516), 
        .A(DP_mult_205_n517), .ZN(DP_mult_205_n515) );
  OAI21_X1 DP_mult_205_U2754 ( .B1(DP_mult_205_n536), .B2(DP_mult_205_n2157), 
        .A(DP_mult_205_n2225), .ZN(DP_mult_205_n504) );
  XNOR2_X1 DP_mult_205_U2753 ( .A(DP_mult_205_n533), .B(DP_mult_205_n320), 
        .ZN(DP_sw1_coeff_ret1[4]) );
  XNOR2_X1 DP_mult_205_U2752 ( .A(DP_sw1_11_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1594) );
  XNOR2_X1 DP_mult_205_U2751 ( .A(DP_sw1_21_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1584) );
  XNOR2_X1 DP_mult_205_U2750 ( .A(DP_sw1_19_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1586) );
  OAI22_X1 DP_mult_205_U2749 ( .A1(DP_mult_205_n2240), .A2(DP_mult_205_n1558), 
        .B1(DP_mult_205_n1557), .B2(DP_mult_205_n2263), .ZN(DP_mult_205_n706)
         );
  XNOR2_X1 DP_mult_205_U2748 ( .A(DP_sw1_15_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1590) );
  XNOR2_X1 DP_mult_205_U2747 ( .A(DP_sw1_13_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1592) );
  XNOR2_X1 DP_mult_205_U2746 ( .A(DP_sw1_17_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1588) );
  OAI22_X1 DP_mult_205_U2745 ( .A1(DP_mult_205_n2179), .A2(DP_mult_205_n1568), 
        .B1(DP_mult_205_n1567), .B2(DP_mult_205_n2262), .ZN(DP_mult_205_n1276)
         );
  OAI22_X1 DP_mult_205_U2744 ( .A1(DP_mult_205_n2240), .A2(DP_mult_205_n1562), 
        .B1(DP_mult_205_n1561), .B2(DP_mult_205_n2263), .ZN(DP_mult_205_n1270)
         );
  OAI22_X1 DP_mult_205_U2743 ( .A1(DP_mult_205_n2239), .A2(DP_mult_205_n1559), 
        .B1(DP_mult_205_n2263), .B2(DP_mult_205_n1558), .ZN(DP_mult_205_n1267)
         );
  OAI22_X1 DP_mult_205_U2742 ( .A1(DP_mult_205_n2180), .A2(DP_mult_205_n1565), 
        .B1(DP_mult_205_n2263), .B2(DP_mult_205_n1564), .ZN(DP_mult_205_n1273)
         );
  OAI22_X1 DP_mult_205_U2741 ( .A1(DP_mult_205_n1581), .A2(DP_mult_205_n2263), 
        .B1(DP_mult_205_n2239), .B2(DP_mult_205_n2317), .ZN(DP_mult_205_n1185)
         );
  OAI22_X1 DP_mult_205_U2740 ( .A1(DP_mult_205_n2240), .A2(DP_mult_205_n1560), 
        .B1(DP_mult_205_n1559), .B2(DP_mult_205_n2262), .ZN(DP_mult_205_n1268)
         );
  OAI22_X1 DP_mult_205_U2739 ( .A1(DP_mult_205_n2180), .A2(DP_mult_205_n1564), 
        .B1(DP_mult_205_n1563), .B2(DP_mult_205_n2263), .ZN(DP_mult_205_n1272)
         );
  OAI22_X1 DP_mult_205_U2738 ( .A1(DP_mult_205_n2239), .A2(DP_mult_205_n1561), 
        .B1(DP_mult_205_n2262), .B2(DP_mult_205_n1560), .ZN(DP_mult_205_n1269)
         );
  OAI22_X1 DP_mult_205_U2737 ( .A1(DP_mult_205_n2239), .A2(DP_mult_205_n1566), 
        .B1(DP_mult_205_n1565), .B2(DP_mult_205_n2262), .ZN(DP_mult_205_n1274)
         );
  OAI22_X1 DP_mult_205_U2736 ( .A1(DP_mult_205_n2240), .A2(DP_mult_205_n1567), 
        .B1(DP_mult_205_n2262), .B2(DP_mult_205_n1566), .ZN(DP_mult_205_n1275)
         );
  OAI22_X1 DP_mult_205_U2735 ( .A1(DP_mult_205_n2180), .A2(DP_mult_205_n1563), 
        .B1(DP_mult_205_n2262), .B2(DP_mult_205_n1562), .ZN(DP_mult_205_n1271)
         );
  NAND2_X1 DP_mult_205_U2734 ( .A1(DP_mult_205_n694), .A2(DP_mult_205_n689), 
        .ZN(DP_mult_205_n378) );
  NAND2_X1 DP_mult_205_U2733 ( .A1(DP_mult_205_n2193), .A2(DP_mult_205_n2195), 
        .ZN(DP_mult_205_n364) );
  NAND2_X1 DP_mult_205_U2732 ( .A1(DP_mult_205_n382), .A2(DP_mult_205_n2193), 
        .ZN(DP_mult_205_n371) );
  AOI21_X1 DP_mult_205_U2731 ( .B1(DP_mult_205_n383), .B2(DP_mult_205_n2193), 
        .A(DP_mult_205_n376), .ZN(DP_mult_205_n372) );
  NAND2_X1 DP_mult_205_U2730 ( .A1(DP_mult_205_n2193), .A2(DP_mult_205_n378), 
        .ZN(DP_mult_205_n305) );
  INV_X1 DP_mult_205_U2729 ( .A(DP_mult_205_n325), .ZN(DP_sw1_coeff_ret1[23])
         );
  OAI21_X1 DP_mult_205_U2728 ( .B1(DP_mult_205_n506), .B2(DP_mult_205_n452), 
        .A(DP_mult_205_n453), .ZN(DP_mult_205_n451) );
  OAI22_X1 DP_mult_205_U2727 ( .A1(DP_mult_205_n2251), .A2(DP_mult_205_n1733), 
        .B1(DP_mult_205_n1732), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n916)
         );
  XNOR2_X1 DP_mult_205_U2726 ( .A(DP_sw1_15_), .B(DP_mult_205_n2302), .ZN(
        DP_mult_205_n1640) );
  XNOR2_X1 DP_mult_205_U2725 ( .A(DP_sw1_13_), .B(DP_mult_205_n2303), .ZN(
        DP_mult_205_n1642) );
  XNOR2_X1 DP_mult_205_U2724 ( .A(DP_sw1_11_), .B(DP_mult_205_n2302), .ZN(
        DP_mult_205_n1644) );
  XNOR2_X1 DP_mult_205_U2723 ( .A(DP_sw1_17_), .B(DP_mult_205_n2303), .ZN(
        DP_mult_205_n1638) );
  OAI22_X1 DP_mult_205_U2722 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1608), 
        .B1(DP_mult_205_n1607), .B2(DP_mult_205_n2267), .ZN(DP_mult_205_n746)
         );
  XNOR2_X1 DP_mult_205_U2721 ( .A(DP_sw1_21_), .B(DP_mult_205_n2303), .ZN(
        DP_mult_205_n1634) );
  XNOR2_X1 DP_mult_205_U2720 ( .A(DP_sw1_19_), .B(DP_mult_205_n2303), .ZN(
        DP_mult_205_n1636) );
  OAI22_X1 DP_mult_205_U2719 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1609), 
        .B1(DP_mult_205_n2267), .B2(DP_mult_205_n1608), .ZN(DP_mult_205_n1315)
         );
  OAI22_X1 DP_mult_205_U2718 ( .A1(DP_mult_205_n1995), .A2(DP_mult_205_n1618), 
        .B1(DP_mult_205_n1617), .B2(DP_mult_205_n2268), .ZN(DP_mult_205_n1324)
         );
  OAI22_X1 DP_mult_205_U2717 ( .A1(DP_mult_205_n1631), .A2(DP_mult_205_n2268), 
        .B1(DP_mult_205_n2130), .B2(DP_mult_205_n1965), .ZN(DP_mult_205_n1187)
         );
  OAI22_X1 DP_mult_205_U2716 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1611), 
        .B1(DP_mult_205_n2268), .B2(DP_mult_205_n1610), .ZN(DP_mult_205_n1317)
         );
  OAI22_X1 DP_mult_205_U2715 ( .A1(DP_mult_205_n2242), .A2(DP_mult_205_n1616), 
        .B1(DP_mult_205_n1615), .B2(DP_mult_205_n2268), .ZN(DP_mult_205_n1322)
         );
  OAI22_X1 DP_mult_205_U2714 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1615), 
        .B1(DP_mult_205_n2267), .B2(DP_mult_205_n1614), .ZN(DP_mult_205_n1321)
         );
  OAI22_X1 DP_mult_205_U2713 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1612), 
        .B1(DP_mult_205_n1611), .B2(DP_mult_205_n2268), .ZN(DP_mult_205_n1318)
         );
  OAI22_X1 DP_mult_205_U2712 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1617), 
        .B1(DP_mult_205_n2268), .B2(DP_mult_205_n1616), .ZN(DP_mult_205_n1323)
         );
  OAI22_X1 DP_mult_205_U2711 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1610), 
        .B1(DP_mult_205_n1609), .B2(DP_mult_205_n2267), .ZN(DP_mult_205_n1316)
         );
  OAI22_X1 DP_mult_205_U2710 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1613), 
        .B1(DP_mult_205_n2267), .B2(DP_mult_205_n1612), .ZN(DP_mult_205_n1319)
         );
  NAND2_X1 DP_mult_205_U2709 ( .A1(DP_mult_205_n717), .A2(DP_mult_205_n726), 
        .ZN(DP_mult_205_n418) );
  AOI21_X1 DP_mult_205_U2708 ( .B1(DP_mult_205_n346), .B2(DP_mult_205_n2197), 
        .A(DP_mult_205_n339), .ZN(DP_mult_205_n337) );
  NAND2_X1 DP_mult_205_U2707 ( .A1(DP_mult_205_n422), .A2(DP_mult_205_n2187), 
        .ZN(DP_mult_205_n411) );
  AOI21_X1 DP_mult_205_U2706 ( .B1(DP_mult_205_n423), .B2(DP_mult_205_n2187), 
        .A(DP_mult_205_n416), .ZN(DP_mult_205_n412) );
  INV_X1 DP_mult_205_U2705 ( .A(DP_mult_205_n346), .ZN(DP_mult_205_n344) );
  NAND2_X1 DP_mult_205_U2704 ( .A1(DP_mult_205_n2187), .A2(DP_mult_205_n418), 
        .ZN(DP_mult_205_n309) );
  OAI22_X1 DP_mult_205_U2703 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1605), 
        .B1(DP_mult_205_n1604), .B2(DP_mult_205_n1933), .ZN(DP_mult_205_n1312)
         );
  NAND2_X1 DP_mult_205_U2702 ( .A1(DP_mult_205_n454), .A2(DP_mult_205_n489), 
        .ZN(DP_mult_205_n452) );
  OAI22_X1 DP_mult_205_U2701 ( .A1(DP_mult_205_n2236), .A2(DP_mult_205_n1528), 
        .B1(DP_mult_205_n1527), .B2(DP_mult_205_n2208), .ZN(DP_mult_205_n1238)
         );
  OAI22_X1 DP_mult_205_U2700 ( .A1(DP_mult_205_n2236), .A2(DP_mult_205_n1527), 
        .B1(DP_mult_205_n2256), .B2(DP_mult_205_n1526), .ZN(DP_mult_205_n1237)
         );
  OAI22_X1 DP_mult_205_U2699 ( .A1(DP_mult_205_n2236), .A2(DP_mult_205_n1530), 
        .B1(DP_mult_205_n1529), .B2(DP_mult_205_n2208), .ZN(DP_mult_205_n1240)
         );
  OAI22_X1 DP_mult_205_U2698 ( .A1(DP_mult_205_n2236), .A2(DP_mult_205_n1526), 
        .B1(DP_mult_205_n1525), .B2(DP_mult_205_n2256), .ZN(DP_mult_205_n1236)
         );
  OAI22_X1 DP_mult_205_U2697 ( .A1(DP_mult_205_n2236), .A2(DP_mult_205_n1529), 
        .B1(DP_mult_205_n2256), .B2(DP_mult_205_n1528), .ZN(DP_mult_205_n1239)
         );
  OAI22_X1 DP_mult_205_U2696 ( .A1(DP_mult_205_n2236), .A2(DP_mult_205_n1524), 
        .B1(DP_mult_205_n1523), .B2(DP_mult_205_n2256), .ZN(DP_mult_205_n1234)
         );
  OAI22_X1 DP_mult_205_U2695 ( .A1(DP_mult_205_n2236), .A2(DP_mult_205_n1523), 
        .B1(DP_mult_205_n2256), .B2(DP_mult_205_n1522), .ZN(DP_mult_205_n1233)
         );
  OAI22_X1 DP_mult_205_U2694 ( .A1(DP_mult_205_n2236), .A2(DP_mult_205_n1525), 
        .B1(DP_mult_205_n2256), .B2(DP_mult_205_n1524), .ZN(DP_mult_205_n1235)
         );
  OAI22_X1 DP_mult_205_U2693 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1519), 
        .B1(DP_mult_205_n2257), .B2(DP_mult_205_n1518), .ZN(DP_mult_205_n1229)
         );
  OAI22_X1 DP_mult_205_U2692 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1520), 
        .B1(DP_mult_205_n1519), .B2(DP_mult_205_n2256), .ZN(DP_mult_205_n1230)
         );
  OAI22_X1 DP_mult_205_U2691 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1521), 
        .B1(DP_mult_205_n2257), .B2(DP_mult_205_n1520), .ZN(DP_mult_205_n1231)
         );
  OAI22_X1 DP_mult_205_U2690 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1522), 
        .B1(DP_mult_205_n1521), .B2(DP_mult_205_n2256), .ZN(DP_mult_205_n1232)
         );
  NOR2_X1 DP_mult_205_U2689 ( .A1(DP_mult_205_n897), .A2(DP_mult_205_n918), 
        .ZN(DP_mult_205_n534) );
  XNOR2_X1 DP_mult_205_U2688 ( .A(DP_mult_205_n430), .B(DP_mult_205_n310), 
        .ZN(DP_sw1_coeff_ret1[14]) );
  XNOR2_X1 DP_mult_205_U2687 ( .A(DP_sw1_13_), .B(DP_mult_205_n2316), .ZN(
        DP_mult_205_n1567) );
  XNOR2_X1 DP_mult_205_U2686 ( .A(DP_sw1_11_), .B(DP_mult_205_n2315), .ZN(
        DP_mult_205_n1569) );
  XNOR2_X1 DP_mult_205_U2685 ( .A(DP_sw1_19_), .B(DP_mult_205_n2314), .ZN(
        DP_mult_205_n1561) );
  XNOR2_X1 DP_mult_205_U2684 ( .A(DP_sw1_15_), .B(DP_mult_205_n2316), .ZN(
        DP_mult_205_n1565) );
  XNOR2_X1 DP_mult_205_U2683 ( .A(DP_sw1_21_), .B(DP_mult_205_n2315), .ZN(
        DP_mult_205_n1559) );
  XNOR2_X1 DP_mult_205_U2682 ( .A(DP_sw1_17_), .B(DP_mult_205_n2313), .ZN(
        DP_mult_205_n1563) );
  OAI22_X1 DP_mult_205_U2681 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1553), 
        .B1(DP_mult_205_n1552), .B2(DP_mult_205_n2259), .ZN(DP_mult_205_n1262)
         );
  OAI22_X1 DP_mult_205_U2680 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1554), 
        .B1(DP_mult_205_n2259), .B2(DP_mult_205_n1553), .ZN(DP_mult_205_n1263)
         );
  OAI22_X1 DP_mult_205_U2679 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1551), 
        .B1(DP_mult_205_n1550), .B2(DP_mult_205_n2260), .ZN(DP_mult_205_n1260)
         );
  OAI22_X1 DP_mult_205_U2678 ( .A1(DP_mult_205_n2172), .A2(DP_mult_205_n1545), 
        .B1(DP_mult_205_n1544), .B2(DP_mult_205_n2259), .ZN(DP_mult_205_n1254)
         );
  OAI22_X1 DP_mult_205_U2677 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1550), 
        .B1(DP_mult_205_n2260), .B2(DP_mult_205_n1549), .ZN(DP_mult_205_n1259)
         );
  OAI22_X1 DP_mult_205_U2676 ( .A1(DP_mult_205_n2237), .A2(DP_mult_205_n1555), 
        .B1(DP_mult_205_n1554), .B2(DP_mult_205_n2260), .ZN(DP_mult_205_n1264)
         );
  OAI22_X1 DP_mult_205_U2675 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1549), 
        .B1(DP_mult_205_n1548), .B2(DP_mult_205_n2259), .ZN(DP_mult_205_n1258)
         );
  OAI22_X1 DP_mult_205_U2674 ( .A1(DP_mult_205_n2172), .A2(DP_mult_205_n1547), 
        .B1(DP_mult_205_n1546), .B2(DP_mult_205_n2259), .ZN(DP_mult_205_n1256)
         );
  OAI22_X1 DP_mult_205_U2673 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1546), 
        .B1(DP_mult_205_n2260), .B2(DP_mult_205_n1545), .ZN(DP_mult_205_n1255)
         );
  OAI22_X1 DP_mult_205_U2672 ( .A1(DP_mult_205_n2172), .A2(DP_mult_205_n1552), 
        .B1(DP_mult_205_n2260), .B2(DP_mult_205_n1551), .ZN(DP_mult_205_n1261)
         );
  OAI22_X1 DP_mult_205_U2671 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1548), 
        .B1(DP_mult_205_n2259), .B2(DP_mult_205_n1547), .ZN(DP_mult_205_n1257)
         );
  OAI22_X1 DP_mult_205_U2670 ( .A1(DP_mult_205_n2237), .A2(DP_mult_205_n1544), 
        .B1(DP_mult_205_n2259), .B2(DP_mult_205_n1543), .ZN(DP_mult_205_n1253)
         );
  OAI22_X1 DP_mult_205_U2669 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1742), 
        .B1(DP_mult_205_n2278), .B2(DP_mult_205_n1741), .ZN(DP_mult_205_n1443)
         );
  OAI22_X1 DP_mult_205_U2668 ( .A1(DP_mult_205_n2251), .A2(DP_mult_205_n1743), 
        .B1(DP_mult_205_n1742), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n1444)
         );
  OAI22_X1 DP_mult_205_U2667 ( .A1(DP_mult_205_n2251), .A2(DP_mult_205_n1737), 
        .B1(DP_mult_205_n1736), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n1438)
         );
  OAI22_X1 DP_mult_205_U2666 ( .A1(DP_mult_205_n1987), .A2(DP_mult_205_n1739), 
        .B1(DP_mult_205_n1738), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n1440)
         );
  OAI22_X1 DP_mult_205_U2665 ( .A1(DP_mult_205_n1987), .A2(DP_mult_205_n1734), 
        .B1(DP_mult_205_n2279), .B2(DP_mult_205_n1733), .ZN(DP_mult_205_n1435)
         );
  OAI22_X1 DP_mult_205_U2664 ( .A1(DP_mult_205_n1987), .A2(DP_mult_205_n1736), 
        .B1(DP_mult_205_n2279), .B2(DP_mult_205_n1735), .ZN(DP_mult_205_n1437)
         );
  INV_X1 DP_mult_205_U2663 ( .A(DP_mult_205_n916), .ZN(DP_mult_205_n917) );
  OAI22_X1 DP_mult_205_U2662 ( .A1(DP_mult_205_n1987), .A2(DP_mult_205_n1735), 
        .B1(DP_mult_205_n1734), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n1436)
         );
  OAI22_X1 DP_mult_205_U2661 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1740), 
        .B1(DP_mult_205_n2278), .B2(DP_mult_205_n1739), .ZN(DP_mult_205_n1441)
         );
  OAI22_X1 DP_mult_205_U2660 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1741), 
        .B1(DP_mult_205_n1740), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n1442)
         );
  OAI22_X1 DP_mult_205_U2659 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1738), 
        .B1(DP_mult_205_n2279), .B2(DP_mult_205_n1737), .ZN(DP_mult_205_n1439)
         );
  OAI22_X1 DP_mult_205_U2658 ( .A1(DP_mult_205_n1756), .A2(DP_mult_205_n1973), 
        .B1(DP_mult_205_n2073), .B2(DP_mult_205_n2289), .ZN(DP_mult_205_n1192)
         );
  OAI22_X1 DP_mult_205_U2657 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1668), 
        .B1(DP_mult_205_n1667), .B2(DP_mult_205_n2274), .ZN(DP_mult_205_n1372)
         );
  OAI22_X1 DP_mult_205_U2656 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1659), 
        .B1(DP_mult_205_n2274), .B2(DP_mult_205_n1658), .ZN(DP_mult_205_n1363)
         );
  OAI22_X1 DP_mult_205_U2655 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1666), 
        .B1(DP_mult_205_n1665), .B2(DP_mult_205_n2274), .ZN(DP_mult_205_n1370)
         );
  OAI22_X1 DP_mult_205_U2654 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1662), 
        .B1(DP_mult_205_n1661), .B2(DP_mult_205_n2273), .ZN(DP_mult_205_n1366)
         );
  OAI22_X1 DP_mult_205_U2653 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1658), 
        .B1(DP_mult_205_n1657), .B2(DP_mult_205_n2273), .ZN(DP_mult_205_n802)
         );
  OAI22_X1 DP_mult_205_U2652 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1665), 
        .B1(DP_mult_205_n2273), .B2(DP_mult_205_n1664), .ZN(DP_mult_205_n1369)
         );
  OAI22_X1 DP_mult_205_U2651 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1667), 
        .B1(DP_mult_205_n2274), .B2(DP_mult_205_n1666), .ZN(DP_mult_205_n1371)
         );
  OAI22_X1 DP_mult_205_U2650 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1664), 
        .B1(DP_mult_205_n1663), .B2(DP_mult_205_n2273), .ZN(DP_mult_205_n1368)
         );
  OAI22_X1 DP_mult_205_U2649 ( .A1(DP_mult_205_n1681), .A2(DP_mult_205_n2274), 
        .B1(DP_mult_205_n2174), .B2(DP_mult_205_n2070), .ZN(DP_mult_205_n1189)
         );
  OAI22_X1 DP_mult_205_U2648 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1663), 
        .B1(DP_mult_205_n2273), .B2(DP_mult_205_n1662), .ZN(DP_mult_205_n1367)
         );
  OAI22_X1 DP_mult_205_U2647 ( .A1(DP_mult_205_n2174), .A2(DP_mult_205_n1660), 
        .B1(DP_mult_205_n1659), .B2(DP_mult_205_n2273), .ZN(DP_mult_205_n1364)
         );
  OAI22_X1 DP_mult_205_U2646 ( .A1(DP_mult_205_n2099), .A2(DP_mult_205_n1661), 
        .B1(DP_mult_205_n2274), .B2(DP_mult_205_n1660), .ZN(DP_mult_205_n1365)
         );
  NAND2_X1 DP_mult_205_U2645 ( .A1(DP_mult_205_n877), .A2(DP_mult_205_n896), 
        .ZN(DP_mult_205_n532) );
  XNOR2_X1 DP_mult_205_U2644 ( .A(DP_mult_205_n419), .B(DP_mult_205_n309), 
        .ZN(DP_sw1_coeff_ret1[15]) );
  XNOR2_X1 DP_mult_205_U2643 ( .A(DP_sw1_15_), .B(DP_mult_205_n2322), .ZN(
        DP_mult_205_n1515) );
  XNOR2_X1 DP_mult_205_U2642 ( .A(DP_sw1_19_), .B(DP_mult_205_n2322), .ZN(
        DP_mult_205_n1511) );
  XNOR2_X1 DP_mult_205_U2641 ( .A(DP_sw1_21_), .B(DP_mult_205_n2323), .ZN(
        DP_mult_205_n1509) );
  XNOR2_X1 DP_mult_205_U2640 ( .A(DP_sw1_13_), .B(DP_mult_205_n2323), .ZN(
        DP_mult_205_n1517) );
  XNOR2_X1 DP_mult_205_U2639 ( .A(DP_sw1_17_), .B(DP_mult_205_n2322), .ZN(
        DP_mult_205_n1513) );
  XNOR2_X1 DP_mult_205_U2638 ( .A(DP_sw1_11_), .B(DP_mult_205_n2322), .ZN(
        DP_mult_205_n1519) );
  OAI22_X1 DP_mult_205_U2637 ( .A1(DP_mult_205_n2177), .A2(DP_mult_205_n1498), 
        .B1(DP_mult_205_n2255), .B2(DP_mult_205_n1497), .ZN(DP_mult_205_n1209)
         );
  OAI22_X1 DP_mult_205_U2636 ( .A1(DP_mult_205_n2233), .A2(DP_mult_205_n1503), 
        .B1(DP_mult_205_n1502), .B2(DP_mult_205_n2254), .ZN(DP_mult_205_n1214)
         );
  OAI22_X1 DP_mult_205_U2635 ( .A1(DP_mult_205_n2177), .A2(DP_mult_205_n1499), 
        .B1(DP_mult_205_n1498), .B2(DP_mult_205_n2255), .ZN(DP_mult_205_n1210)
         );
  OAI22_X1 DP_mult_205_U2634 ( .A1(DP_mult_205_n2234), .A2(DP_mult_205_n1504), 
        .B1(DP_mult_205_n2255), .B2(DP_mult_205_n1503), .ZN(DP_mult_205_n1215)
         );
  OAI22_X1 DP_mult_205_U2633 ( .A1(DP_mult_205_n1506), .A2(DP_mult_205_n2254), 
        .B1(DP_mult_205_n2234), .B2(DP_mult_205_n1939), .ZN(DP_mult_205_n1182)
         );
  OAI22_X1 DP_mult_205_U2632 ( .A1(DP_mult_205_n2178), .A2(DP_mult_205_n1500), 
        .B1(DP_mult_205_n2255), .B2(DP_mult_205_n1499), .ZN(DP_mult_205_n1211)
         );
  OAI22_X1 DP_mult_205_U2631 ( .A1(DP_mult_205_n2234), .A2(DP_mult_205_n1505), 
        .B1(DP_mult_205_n1504), .B2(DP_mult_205_n2254), .ZN(DP_mult_205_n1216)
         );
  OAI22_X1 DP_mult_205_U2630 ( .A1(DP_mult_205_n2233), .A2(DP_mult_205_n1493), 
        .B1(DP_mult_205_n1492), .B2(DP_mult_205_n2254), .ZN(DP_mult_205_n1204)
         );
  OAI22_X1 DP_mult_205_U2629 ( .A1(DP_mult_205_n2234), .A2(DP_mult_205_n1501), 
        .B1(DP_mult_205_n1500), .B2(DP_mult_205_n2254), .ZN(DP_mult_205_n1212)
         );
  OAI22_X1 DP_mult_205_U2628 ( .A1(DP_mult_205_n2177), .A2(DP_mult_205_n1489), 
        .B1(DP_mult_205_n1488), .B2(DP_mult_205_n2255), .ZN(DP_mult_205_n1200)
         );
  OAI22_X1 DP_mult_205_U2627 ( .A1(DP_mult_205_n2177), .A2(DP_mult_205_n1502), 
        .B1(DP_mult_205_n2255), .B2(DP_mult_205_n1501), .ZN(DP_mult_205_n1213)
         );
  OAI22_X1 DP_mult_205_U2626 ( .A1(DP_mult_205_n2178), .A2(DP_mult_205_n1496), 
        .B1(DP_mult_205_n2255), .B2(DP_mult_205_n1495), .ZN(DP_mult_205_n1207)
         );
  OAI22_X1 DP_mult_205_U2625 ( .A1(DP_mult_205_n2178), .A2(DP_mult_205_n1494), 
        .B1(DP_mult_205_n2254), .B2(DP_mult_205_n1493), .ZN(DP_mult_205_n1205)
         );
  OAI22_X1 DP_mult_205_U2624 ( .A1(DP_mult_205_n2233), .A2(DP_mult_205_n1497), 
        .B1(DP_mult_205_n1496), .B2(DP_mult_205_n2255), .ZN(DP_mult_205_n1208)
         );
  OAI22_X1 DP_mult_205_U2623 ( .A1(DP_mult_205_n2177), .A2(DP_mult_205_n1495), 
        .B1(DP_mult_205_n1494), .B2(DP_mult_205_n2254), .ZN(DP_mult_205_n1206)
         );
  OAI22_X1 DP_mult_205_U2622 ( .A1(DP_mult_205_n2178), .A2(DP_mult_205_n1487), 
        .B1(DP_mult_205_n1486), .B2(DP_mult_205_n2255), .ZN(DP_mult_205_n1198)
         );
  OAI22_X1 DP_mult_205_U2621 ( .A1(DP_mult_205_n2233), .A2(DP_mult_205_n1491), 
        .B1(DP_mult_205_n1490), .B2(DP_mult_205_n2254), .ZN(DP_mult_205_n1202)
         );
  OAI22_X1 DP_mult_205_U2620 ( .A1(DP_mult_205_n2233), .A2(DP_mult_205_n1485), 
        .B1(DP_mult_205_n1484), .B2(DP_mult_205_n2254), .ZN(DP_mult_205_n1196)
         );
  NAND2_X1 DP_mult_205_U2619 ( .A1(DP_mult_205_n761), .A2(DP_mult_205_n774), 
        .ZN(DP_mult_205_n461) );
  OAI22_X1 DP_mult_205_U2618 ( .A1(DP_mult_205_n2233), .A2(DP_mult_205_n1483), 
        .B1(DP_mult_205_n1482), .B2(DP_mult_205_n2255), .ZN(DP_mult_205_n676)
         );
  XNOR2_X1 DP_mult_205_U2617 ( .A(DP_mult_205_n410), .B(DP_mult_205_n308), 
        .ZN(DP_sw1_coeff_ret1[16]) );
  XNOR2_X1 DP_mult_205_U2616 ( .A(DP_sw1_17_), .B(DP_mult_205_n2318), .ZN(
        DP_mult_205_n1538) );
  XNOR2_X1 DP_mult_205_U2615 ( .A(DP_sw1_15_), .B(DP_mult_205_n2320), .ZN(
        DP_mult_205_n1540) );
  XNOR2_X1 DP_mult_205_U2614 ( .A(DP_sw1_11_), .B(DP_mult_205_n2319), .ZN(
        DP_mult_205_n1544) );
  XNOR2_X1 DP_mult_205_U2613 ( .A(DP_sw1_13_), .B(DP_mult_205_n2320), .ZN(
        DP_mult_205_n1542) );
  XNOR2_X1 DP_mult_205_U2612 ( .A(DP_sw1_19_), .B(DP_mult_205_n2320), .ZN(
        DP_mult_205_n1536) );
  OR2_X1 DP_mult_205_U2611 ( .A1(DP_mult_205_n1215), .A2(DP_mult_205_n1237), 
        .ZN(DP_mult_205_n938) );
  XNOR2_X1 DP_mult_205_U2610 ( .A(DP_sw1_21_), .B(DP_mult_205_n2318), .ZN(
        DP_mult_205_n1534) );
  XNOR2_X1 DP_mult_205_U2609 ( .A(DP_mult_205_n1215), .B(DP_mult_205_n1237), 
        .ZN(DP_mult_205_n939) );
  INV_X1 DP_mult_205_U2608 ( .A(DP_coeffs_fb_int[46]), .ZN(DP_mult_205_n2286)
         );
  AOI21_X1 DP_mult_205_U2607 ( .B1(DP_mult_205_n2010), .B2(DP_mult_205_n490), 
        .A(DP_mult_205_n455), .ZN(DP_mult_205_n453) );
  OAI22_X1 DP_mult_205_U2606 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1604), 
        .B1(DP_mult_205_n2265), .B2(DP_mult_205_n1603), .ZN(DP_mult_205_n1311)
         );
  OAI22_X1 DP_mult_205_U2605 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1599), 
        .B1(DP_mult_205_n1598), .B2(DP_mult_205_n1933), .ZN(DP_mult_205_n1306)
         );
  OAI22_X1 DP_mult_205_U2604 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1597), 
        .B1(DP_mult_205_n1596), .B2(DP_mult_205_n1933), .ZN(DP_mult_205_n1304)
         );
  OAI22_X1 DP_mult_205_U2603 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1598), 
        .B1(DP_mult_205_n2265), .B2(DP_mult_205_n1597), .ZN(DP_mult_205_n1305)
         );
  OAI22_X1 DP_mult_205_U2602 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1603), 
        .B1(DP_mult_205_n1602), .B2(DP_mult_205_n1933), .ZN(DP_mult_205_n1310)
         );
  OAI22_X1 DP_mult_205_U2601 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1595), 
        .B1(DP_mult_205_n1594), .B2(DP_mult_205_n2265), .ZN(DP_mult_205_n1302)
         );
  OAI22_X1 DP_mult_205_U2600 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1594), 
        .B1(DP_mult_205_n2265), .B2(DP_mult_205_n1593), .ZN(DP_mult_205_n1301)
         );
  OAI22_X1 DP_mult_205_U2599 ( .A1(DP_mult_205_n1601), .A2(DP_mult_205_n289), 
        .B1(DP_mult_205_n1600), .B2(DP_mult_205_n2265), .ZN(DP_mult_205_n1308)
         );
  OAI22_X1 DP_mult_205_U2598 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1596), 
        .B1(DP_mult_205_n1933), .B2(DP_mult_205_n1595), .ZN(DP_mult_205_n1303)
         );
  OAI22_X1 DP_mult_205_U2597 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1600), 
        .B1(DP_mult_205_n1933), .B2(DP_mult_205_n1599), .ZN(DP_mult_205_n1307)
         );
  OAI22_X1 DP_mult_205_U2596 ( .A1(DP_mult_205_n289), .A2(DP_mult_205_n1602), 
        .B1(DP_mult_205_n2265), .B2(DP_mult_205_n1601), .ZN(DP_mult_205_n1309)
         );
  XNOR2_X1 DP_mult_205_U2595 ( .A(DP_sw1_19_), .B(DP_mult_205_n2294), .ZN(
        DP_mult_205_n1686) );
  XNOR2_X1 DP_mult_205_U2594 ( .A(DP_sw1_15_), .B(DP_mult_205_n2294), .ZN(
        DP_mult_205_n1690) );
  XNOR2_X1 DP_mult_205_U2593 ( .A(DP_sw1_11_), .B(DP_mult_205_n2294), .ZN(
        DP_mult_205_n1694) );
  XNOR2_X1 DP_mult_205_U2592 ( .A(DP_sw1_13_), .B(DP_mult_205_n2294), .ZN(
        DP_mult_205_n1692) );
  XNOR2_X1 DP_mult_205_U2591 ( .A(DP_coeffs_fb_int[40]), .B(
        DP_coeffs_fb_int[39]), .ZN(DP_mult_205_n259) );
  OAI22_X1 DP_mult_205_U2590 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1755), 
        .B1(DP_mult_205_n1754), .B2(DP_mult_205_n1973), .ZN(DP_mult_205_n1456)
         );
  OAI22_X1 DP_mult_205_U2589 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1751), 
        .B1(DP_mult_205_n1750), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n1452)
         );
  OAI22_X1 DP_mult_205_U2588 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1752), 
        .B1(DP_mult_205_n2278), .B2(DP_mult_205_n1751), .ZN(DP_mult_205_n1453)
         );
  OAI22_X1 DP_mult_205_U2587 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1754), 
        .B1(DP_mult_205_n1973), .B2(DP_mult_205_n1753), .ZN(DP_mult_205_n1455)
         );
  OAI22_X1 DP_mult_205_U2586 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1746), 
        .B1(DP_mult_205_n2279), .B2(DP_mult_205_n1745), .ZN(DP_mult_205_n1447)
         );
  OAI22_X1 DP_mult_205_U2585 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1744), 
        .B1(DP_mult_205_n2279), .B2(DP_mult_205_n1743), .ZN(DP_mult_205_n1445)
         );
  OAI22_X1 DP_mult_205_U2584 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1748), 
        .B1(DP_mult_205_n1973), .B2(DP_mult_205_n1747), .ZN(DP_mult_205_n1449)
         );
  OAI22_X1 DP_mult_205_U2583 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1749), 
        .B1(DP_mult_205_n1748), .B2(DP_mult_205_n1973), .ZN(DP_mult_205_n1450)
         );
  OAI22_X1 DP_mult_205_U2582 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1745), 
        .B1(DP_mult_205_n1744), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n1446)
         );
  OAI22_X1 DP_mult_205_U2581 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1750), 
        .B1(DP_mult_205_n1973), .B2(DP_mult_205_n1749), .ZN(DP_mult_205_n1451)
         );
  OAI22_X1 DP_mult_205_U2580 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1747), 
        .B1(DP_mult_205_n1746), .B2(DP_mult_205_n1973), .ZN(DP_mult_205_n1448)
         );
  OAI22_X1 DP_mult_205_U2579 ( .A1(DP_mult_205_n2073), .A2(DP_mult_205_n1753), 
        .B1(DP_mult_205_n1752), .B2(DP_mult_205_n1973), .ZN(DP_mult_205_n1454)
         );
  OAI21_X1 DP_mult_205_U2578 ( .B1(DP_mult_205_n594), .B2(DP_mult_205_n582), 
        .A(DP_mult_205_n583), .ZN(DP_mult_205_n581) );
  OAI22_X1 DP_mult_205_U2577 ( .A1(DP_mult_205_n2176), .A2(DP_mult_205_n1646), 
        .B1(DP_mult_205_n2271), .B2(DP_mult_205_n1645), .ZN(DP_mult_205_n1351)
         );
  OAI22_X1 DP_mult_205_U2576 ( .A1(DP_mult_205_n2176), .A2(DP_mult_205_n1651), 
        .B1(DP_mult_205_n1650), .B2(DP_mult_205_n2270), .ZN(DP_mult_205_n1356)
         );
  OAI22_X1 DP_mult_205_U2575 ( .A1(DP_mult_205_n2244), .A2(DP_mult_205_n1644), 
        .B1(DP_mult_205_n2270), .B2(DP_mult_205_n1643), .ZN(DP_mult_205_n1349)
         );
  OAI22_X1 DP_mult_205_U2574 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1645), 
        .B1(DP_mult_205_n1644), .B2(DP_mult_205_n2270), .ZN(DP_mult_205_n1350)
         );
  OAI22_X1 DP_mult_205_U2573 ( .A1(DP_mult_205_n1969), .A2(DP_mult_205_n1650), 
        .B1(DP_mult_205_n2271), .B2(DP_mult_205_n1649), .ZN(DP_mult_205_n1355)
         );
  OAI22_X1 DP_mult_205_U2572 ( .A1(DP_mult_205_n1968), .A2(DP_mult_205_n1647), 
        .B1(DP_mult_205_n1646), .B2(DP_mult_205_n2271), .ZN(DP_mult_205_n1352)
         );
  OAI22_X1 DP_mult_205_U2571 ( .A1(DP_mult_205_n1968), .A2(DP_mult_205_n1655), 
        .B1(DP_mult_205_n1654), .B2(DP_mult_205_n2270), .ZN(DP_mult_205_n1360)
         );
  OAI22_X1 DP_mult_205_U2570 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1648), 
        .B1(DP_mult_205_n2270), .B2(DP_mult_205_n1647), .ZN(DP_mult_205_n1353)
         );
  OAI22_X1 DP_mult_205_U2569 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1654), 
        .B1(DP_mult_205_n2270), .B2(DP_mult_205_n1653), .ZN(DP_mult_205_n1359)
         );
  OAI22_X1 DP_mult_205_U2568 ( .A1(DP_mult_205_n2176), .A2(DP_mult_205_n1649), 
        .B1(DP_mult_205_n1648), .B2(DP_mult_205_n2270), .ZN(DP_mult_205_n1354)
         );
  OAI22_X1 DP_mult_205_U2567 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1652), 
        .B1(DP_mult_205_n2271), .B2(DP_mult_205_n1651), .ZN(DP_mult_205_n1357)
         );
  OAI22_X1 DP_mult_205_U2566 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1653), 
        .B1(DP_mult_205_n1652), .B2(DP_mult_205_n2270), .ZN(DP_mult_205_n1358)
         );
  INV_X1 DP_mult_205_U2565 ( .A(DP_mult_205_n746), .ZN(DP_mult_205_n747) );
  NAND2_X1 DP_mult_205_U2564 ( .A1(DP_mult_205_n709), .A2(DP_mult_205_n716), 
        .ZN(DP_mult_205_n409) );
  NAND2_X1 DP_mult_205_U2563 ( .A1(DP_mult_205_n422), .A2(DP_mult_205_n356), 
        .ZN(DP_mult_205_n354) );
  AOI21_X1 DP_mult_205_U2562 ( .B1(DP_mult_205_n423), .B2(DP_mult_205_n356), 
        .A(DP_mult_205_n359), .ZN(DP_mult_205_n355) );
  NAND2_X1 DP_mult_205_U2561 ( .A1(DP_mult_205_n1816), .A2(DP_mult_205_n2277), 
        .ZN(DP_mult_205_n277) );
  XNOR2_X1 DP_mult_205_U2560 ( .A(DP_sw1_19_), .B(DP_mult_205_n2283), .ZN(
        DP_mult_205_n1761) );
  XNOR2_X1 DP_mult_205_U2559 ( .A(DP_sw1_15_), .B(DP_mult_205_n2283), .ZN(
        DP_mult_205_n1765) );
  XNOR2_X1 DP_mult_205_U2558 ( .A(DP_sw1_21_), .B(DP_mult_205_n2283), .ZN(
        DP_mult_205_n1759) );
  XNOR2_X1 DP_mult_205_U2557 ( .A(DP_sw1_11_), .B(DP_mult_205_n2285), .ZN(
        DP_mult_205_n1769) );
  XNOR2_X1 DP_mult_205_U2556 ( .A(DP_sw1_17_), .B(DP_mult_205_n2283), .ZN(
        DP_mult_205_n1763) );
  XNOR2_X1 DP_mult_205_U2555 ( .A(DP_sw1_13_), .B(DP_mult_205_n2285), .ZN(
        DP_mult_205_n1767) );
  NAND2_X1 DP_mult_205_U2554 ( .A1(DP_mult_205_n805), .A2(DP_mult_205_n1936), 
        .ZN(DP_mult_205_n496) );
  XNOR2_X1 DP_mult_205_U2553 ( .A(DP_mult_205_n397), .B(DP_mult_205_n307), 
        .ZN(DP_sw1_coeff_ret1[17]) );
  OAI22_X1 DP_mult_205_U2552 ( .A1(DP_mult_205_n1968), .A2(DP_mult_205_n1643), 
        .B1(DP_mult_205_n1642), .B2(DP_mult_205_n2270), .ZN(DP_mult_205_n1348)
         );
  OAI22_X1 DP_mult_205_U2551 ( .A1(DP_mult_205_n1969), .A2(DP_mult_205_n1641), 
        .B1(DP_mult_205_n1640), .B2(DP_mult_205_n2271), .ZN(DP_mult_205_n1346)
         );
  OAI22_X1 DP_mult_205_U2550 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1633), 
        .B1(DP_mult_205_n1632), .B2(DP_mult_205_n2271), .ZN(DP_mult_205_n772)
         );
  OAI22_X1 DP_mult_205_U2549 ( .A1(DP_mult_205_n1656), .A2(DP_mult_205_n2270), 
        .B1(DP_mult_205_n2175), .B2(DP_mult_205_n2104), .ZN(DP_mult_205_n1188)
         );
  OAI22_X1 DP_mult_205_U2548 ( .A1(DP_mult_205_n2244), .A2(DP_mult_205_n1642), 
        .B1(DP_mult_205_n2270), .B2(DP_mult_205_n1641), .ZN(DP_mult_205_n1347)
         );
  OAI22_X1 DP_mult_205_U2547 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1640), 
        .B1(DP_mult_205_n2271), .B2(DP_mult_205_n1639), .ZN(DP_mult_205_n1345)
         );
  OAI22_X1 DP_mult_205_U2546 ( .A1(DP_mult_205_n2244), .A2(DP_mult_205_n1639), 
        .B1(DP_mult_205_n1638), .B2(DP_mult_205_n2271), .ZN(DP_mult_205_n1344)
         );
  OAI22_X1 DP_mult_205_U2545 ( .A1(DP_mult_205_n1969), .A2(DP_mult_205_n1638), 
        .B1(DP_mult_205_n2270), .B2(DP_mult_205_n1637), .ZN(DP_mult_205_n1343)
         );
  OAI22_X1 DP_mult_205_U2544 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1635), 
        .B1(DP_mult_205_n1634), .B2(DP_mult_205_n2271), .ZN(DP_mult_205_n1340)
         );
  OAI22_X1 DP_mult_205_U2543 ( .A1(DP_mult_205_n1969), .A2(DP_mult_205_n1634), 
        .B1(DP_mult_205_n2271), .B2(DP_mult_205_n1633), .ZN(DP_mult_205_n1339)
         );
  OAI22_X1 DP_mult_205_U2542 ( .A1(DP_mult_205_n2175), .A2(DP_mult_205_n1636), 
        .B1(DP_mult_205_n2271), .B2(DP_mult_205_n1635), .ZN(DP_mult_205_n1341)
         );
  OAI22_X1 DP_mult_205_U2541 ( .A1(DP_mult_205_n1968), .A2(DP_mult_205_n1637), 
        .B1(DP_mult_205_n1636), .B2(DP_mult_205_n2270), .ZN(DP_mult_205_n1342)
         );
  OAI22_X1 DP_mult_205_U2540 ( .A1(DP_mult_205_n1606), .A2(DP_mult_205_n2265), 
        .B1(DP_mult_205_n2079), .B2(DP_mult_205_n2312), .ZN(DP_mult_205_n1186)
         );
  OAI22_X1 DP_mult_205_U2539 ( .A1(DP_mult_205_n2078), .A2(DP_mult_205_n1586), 
        .B1(DP_mult_205_n2265), .B2(DP_mult_205_n1585), .ZN(DP_mult_205_n1293)
         );
  OAI22_X1 DP_mult_205_U2538 ( .A1(DP_mult_205_n2079), .A2(DP_mult_205_n1591), 
        .B1(DP_mult_205_n1590), .B2(DP_mult_205_n1933), .ZN(DP_mult_205_n1298)
         );
  OAI22_X1 DP_mult_205_U2537 ( .A1(DP_mult_205_n2241), .A2(DP_mult_205_n1587), 
        .B1(DP_mult_205_n1586), .B2(DP_mult_205_n2265), .ZN(DP_mult_205_n1294)
         );
  OAI22_X1 DP_mult_205_U2536 ( .A1(DP_mult_205_n2079), .A2(DP_mult_205_n1592), 
        .B1(DP_mult_205_n1933), .B2(DP_mult_205_n1591), .ZN(DP_mult_205_n1299)
         );
  OAI22_X1 DP_mult_205_U2535 ( .A1(DP_mult_205_n2078), .A2(DP_mult_205_n1583), 
        .B1(DP_mult_205_n1582), .B2(DP_mult_205_n1933), .ZN(DP_mult_205_n724)
         );
  OAI22_X1 DP_mult_205_U2534 ( .A1(DP_mult_205_n2078), .A2(DP_mult_205_n1588), 
        .B1(DP_mult_205_n1933), .B2(DP_mult_205_n1587), .ZN(DP_mult_205_n1295)
         );
  OAI22_X1 DP_mult_205_U2533 ( .A1(DP_mult_205_n2241), .A2(DP_mult_205_n1585), 
        .B1(DP_mult_205_n1584), .B2(DP_mult_205_n2265), .ZN(DP_mult_205_n1292)
         );
  OAI22_X1 DP_mult_205_U2532 ( .A1(DP_mult_205_n2241), .A2(DP_mult_205_n1589), 
        .B1(DP_mult_205_n1588), .B2(DP_mult_205_n2265), .ZN(DP_mult_205_n1296)
         );
  OAI22_X1 DP_mult_205_U2531 ( .A1(DP_mult_205_n2241), .A2(DP_mult_205_n1584), 
        .B1(DP_mult_205_n1933), .B2(DP_mult_205_n1583), .ZN(DP_mult_205_n1291)
         );
  OAI22_X1 DP_mult_205_U2530 ( .A1(DP_mult_205_n2078), .A2(DP_mult_205_n1590), 
        .B1(DP_mult_205_n1933), .B2(DP_mult_205_n1589), .ZN(DP_mult_205_n1297)
         );
  OAI22_X1 DP_mult_205_U2529 ( .A1(DP_mult_205_n2078), .A2(DP_mult_205_n1593), 
        .B1(DP_mult_205_n1592), .B2(DP_mult_205_n1933), .ZN(DP_mult_205_n1300)
         );
  OAI21_X1 DP_mult_205_U2528 ( .B1(DP_mult_205_n2227), .B2(DP_mult_205_n550), 
        .A(DP_mult_205_n543), .ZN(DP_mult_205_n541) );
  OAI21_X1 DP_mult_205_U2527 ( .B1(DP_mult_205_n2072), .B2(DP_mult_205_n538), 
        .A(DP_mult_205_n539), .ZN(DP_mult_205_n537) );
  OAI22_X1 DP_mult_205_U2526 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1628), 
        .B1(DP_mult_205_n1627), .B2(DP_mult_205_n2268), .ZN(DP_mult_205_n1334)
         );
  OAI22_X1 DP_mult_205_U2525 ( .A1(DP_mult_205_n2239), .A2(DP_mult_205_n1574), 
        .B1(DP_mult_205_n1573), .B2(DP_mult_205_n2262), .ZN(DP_mult_205_n1282)
         );
  OAI22_X1 DP_mult_205_U2524 ( .A1(DP_mult_205_n2179), .A2(DP_mult_205_n1576), 
        .B1(DP_mult_205_n1575), .B2(DP_mult_205_n2262), .ZN(DP_mult_205_n1284)
         );
  OAI22_X1 DP_mult_205_U2523 ( .A1(DP_mult_205_n2179), .A2(DP_mult_205_n1572), 
        .B1(DP_mult_205_n1571), .B2(DP_mult_205_n2263), .ZN(DP_mult_205_n1280)
         );
  OAI22_X1 DP_mult_205_U2522 ( .A1(DP_mult_205_n2239), .A2(DP_mult_205_n1578), 
        .B1(DP_mult_205_n1577), .B2(DP_mult_205_n2262), .ZN(DP_mult_205_n1286)
         );
  OAI22_X1 DP_mult_205_U2521 ( .A1(DP_mult_205_n2179), .A2(DP_mult_205_n1577), 
        .B1(DP_mult_205_n2263), .B2(DP_mult_205_n1576), .ZN(DP_mult_205_n1285)
         );
  OAI22_X1 DP_mult_205_U2520 ( .A1(DP_mult_205_n2240), .A2(DP_mult_205_n1579), 
        .B1(DP_mult_205_n2262), .B2(DP_mult_205_n1578), .ZN(DP_mult_205_n1287)
         );
  OAI22_X1 DP_mult_205_U2519 ( .A1(DP_mult_205_n2240), .A2(DP_mult_205_n1569), 
        .B1(DP_mult_205_n2263), .B2(DP_mult_205_n1568), .ZN(DP_mult_205_n1277)
         );
  OAI22_X1 DP_mult_205_U2518 ( .A1(DP_mult_205_n2180), .A2(DP_mult_205_n1573), 
        .B1(DP_mult_205_n2262), .B2(DP_mult_205_n1572), .ZN(DP_mult_205_n1281)
         );
  OAI22_X1 DP_mult_205_U2517 ( .A1(DP_mult_205_n2180), .A2(DP_mult_205_n1580), 
        .B1(DP_mult_205_n1579), .B2(DP_mult_205_n2262), .ZN(DP_mult_205_n1288)
         );
  OAI22_X1 DP_mult_205_U2516 ( .A1(DP_mult_205_n2240), .A2(DP_mult_205_n1571), 
        .B1(DP_mult_205_n2263), .B2(DP_mult_205_n1570), .ZN(DP_mult_205_n1279)
         );
  OAI22_X1 DP_mult_205_U2515 ( .A1(DP_mult_205_n2239), .A2(DP_mult_205_n1570), 
        .B1(DP_mult_205_n1569), .B2(DP_mult_205_n2262), .ZN(DP_mult_205_n1278)
         );
  OAI22_X1 DP_mult_205_U2514 ( .A1(DP_mult_205_n2180), .A2(DP_mult_205_n1575), 
        .B1(DP_mult_205_n2263), .B2(DP_mult_205_n1574), .ZN(DP_mult_205_n1283)
         );
  OAI22_X1 DP_mult_205_U2513 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1516), 
        .B1(DP_mult_205_n1515), .B2(DP_mult_205_n2208), .ZN(DP_mult_205_n1226)
         );
  OAI22_X1 DP_mult_205_U2512 ( .A1(DP_mult_205_n1531), .A2(DP_mult_205_n2208), 
        .B1(DP_mult_205_n2235), .B2(DP_mult_205_n2007), .ZN(DP_mult_205_n1183)
         );
  OAI22_X1 DP_mult_205_U2511 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1517), 
        .B1(DP_mult_205_n2256), .B2(DP_mult_205_n1516), .ZN(DP_mult_205_n1227)
         );
  OAI22_X1 DP_mult_205_U2510 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1512), 
        .B1(DP_mult_205_n1511), .B2(DP_mult_205_n2208), .ZN(DP_mult_205_n1222)
         );
  OAI22_X1 DP_mult_205_U2509 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1509), 
        .B1(DP_mult_205_n2257), .B2(DP_mult_205_n1508), .ZN(DP_mult_205_n1219)
         );
  OAI22_X1 DP_mult_205_U2508 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1510), 
        .B1(DP_mult_205_n1509), .B2(DP_mult_205_n2208), .ZN(DP_mult_205_n1220)
         );
  OAI22_X1 DP_mult_205_U2507 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1515), 
        .B1(DP_mult_205_n2256), .B2(DP_mult_205_n1514), .ZN(DP_mult_205_n1225)
         );
  OAI22_X1 DP_mult_205_U2506 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1514), 
        .B1(DP_mult_205_n1513), .B2(DP_mult_205_n2208), .ZN(DP_mult_205_n1224)
         );
  OAI22_X1 DP_mult_205_U2505 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1511), 
        .B1(DP_mult_205_n2257), .B2(DP_mult_205_n1510), .ZN(DP_mult_205_n1221)
         );
  OAI22_X1 DP_mult_205_U2504 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1518), 
        .B1(DP_mult_205_n1517), .B2(DP_mult_205_n2208), .ZN(DP_mult_205_n1228)
         );
  OAI22_X1 DP_mult_205_U2503 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1513), 
        .B1(DP_mult_205_n2257), .B2(DP_mult_205_n1512), .ZN(DP_mult_205_n1223)
         );
  OAI22_X1 DP_mult_205_U2502 ( .A1(DP_mult_205_n2235), .A2(DP_mult_205_n1508), 
        .B1(DP_mult_205_n1507), .B2(DP_mult_205_n2208), .ZN(DP_mult_205_n682)
         );
  OAI21_X1 DP_mult_205_U2501 ( .B1(DP_mult_205_n421), .B2(DP_mult_205_n402), 
        .A(DP_mult_205_n405), .ZN(DP_mult_205_n401) );
  OAI21_X1 DP_mult_205_U2500 ( .B1(DP_mult_205_n421), .B2(DP_mult_205_n347), 
        .A(DP_mult_205_n348), .ZN(DP_mult_205_n346) );
  INV_X1 DP_mult_205_U2499 ( .A(DP_mult_205_n421), .ZN(DP_mult_205_n423) );
  XNOR2_X1 DP_mult_205_U2498 ( .A(DP_mult_205_n370), .B(DP_mult_205_n304), 
        .ZN(DP_sw1_coeff_ret1[20]) );
  NAND2_X1 DP_mult_205_U2497 ( .A1(DP_mult_205_n540), .A2(DP_mult_205_n552), 
        .ZN(DP_mult_205_n538) );
  NAND2_X1 DP_mult_205_U2496 ( .A1(DP_mult_205_n963), .A2(DP_mult_205_n982), 
        .ZN(DP_mult_205_n559) );
  OAI22_X1 DP_mult_205_U2495 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1697), 
        .B1(DP_mult_205_n1696), .B2(DP_mult_205_n1982), .ZN(DP_mult_205_n1400)
         );
  OAI22_X1 DP_mult_205_U2494 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1703), 
        .B1(DP_mult_205_n1702), .B2(DP_mult_205_n1983), .ZN(DP_mult_205_n1406)
         );
  OAI22_X1 DP_mult_205_U2493 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1694), 
        .B1(DP_mult_205_n1982), .B2(DP_mult_205_n1693), .ZN(DP_mult_205_n1397)
         );
  OAI22_X1 DP_mult_205_U2492 ( .A1(DP_mult_205_n2248), .A2(DP_mult_205_n1696), 
        .B1(DP_mult_205_n1983), .B2(DP_mult_205_n1695), .ZN(DP_mult_205_n1399)
         );
  OAI22_X1 DP_mult_205_U2491 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1699), 
        .B1(DP_mult_205_n1698), .B2(DP_mult_205_n1982), .ZN(DP_mult_205_n1402)
         );
  OAI22_X1 DP_mult_205_U2490 ( .A1(DP_mult_205_n2248), .A2(DP_mult_205_n1705), 
        .B1(DP_mult_205_n1704), .B2(DP_mult_205_n1982), .ZN(DP_mult_205_n1408)
         );
  OAI22_X1 DP_mult_205_U2489 ( .A1(DP_mult_205_n2095), .A2(DP_mult_205_n1700), 
        .B1(DP_mult_205_n1982), .B2(DP_mult_205_n1699), .ZN(DP_mult_205_n1403)
         );
  OAI22_X1 DP_mult_205_U2488 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1698), 
        .B1(DP_mult_205_n1982), .B2(DP_mult_205_n1697), .ZN(DP_mult_205_n1401)
         );
  OAI22_X1 DP_mult_205_U2487 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1702), 
        .B1(DP_mult_205_n1982), .B2(DP_mult_205_n1701), .ZN(DP_mult_205_n1405)
         );
  OAI22_X1 DP_mult_205_U2486 ( .A1(DP_mult_205_n2096), .A2(DP_mult_205_n1701), 
        .B1(DP_mult_205_n1700), .B2(DP_mult_205_n1982), .ZN(DP_mult_205_n1404)
         );
  OAI22_X1 DP_mult_205_U2485 ( .A1(DP_mult_205_n2171), .A2(DP_mult_205_n1704), 
        .B1(DP_mult_205_n1982), .B2(DP_mult_205_n1703), .ZN(DP_mult_205_n1407)
         );
  OAI22_X1 DP_mult_205_U2484 ( .A1(DP_mult_205_n2095), .A2(DP_mult_205_n1695), 
        .B1(DP_mult_205_n1694), .B2(DP_mult_205_n1982), .ZN(DP_mult_205_n1398)
         );
  OAI21_X1 DP_mult_205_U2483 ( .B1(DP_mult_205_n2094), .B2(DP_mult_205_n1990), 
        .A(DP_mult_205_n2333), .ZN(DP_mult_205_n1386) );
  NAND2_X1 DP_mult_205_U2482 ( .A1(DP_mult_205_n1811), .A2(DP_mult_205_n2266), 
        .ZN(DP_mult_205_n287) );
  XNOR2_X1 DP_mult_205_U2481 ( .A(DP_mult_205_n388), .B(DP_mult_205_n306), 
        .ZN(DP_sw1_coeff_ret1[18]) );
  AOI21_X1 DP_mult_205_U2480 ( .B1(DP_mult_205_n2097), .B2(DP_mult_205_n553), 
        .A(DP_mult_205_n541), .ZN(DP_mult_205_n539) );
  XNOR2_X1 DP_mult_205_U2479 ( .A(DP_mult_205_n379), .B(DP_mult_205_n305), 
        .ZN(DP_sw1_coeff_ret1[19]) );
  XNOR2_X1 DP_mult_205_U2478 ( .A(DP_mult_205_n353), .B(DP_mult_205_n303), 
        .ZN(DP_sw1_coeff_ret1[21]) );
  OAI22_X1 DP_mult_205_U2477 ( .A1(DP_mult_205_n2099), .A2(DP_mult_205_n1678), 
        .B1(DP_mult_205_n1677), .B2(DP_mult_205_n2274), .ZN(DP_mult_205_n1382)
         );
  OAI22_X1 DP_mult_205_U2476 ( .A1(DP_mult_205_n2099), .A2(DP_mult_205_n1673), 
        .B1(DP_mult_205_n2273), .B2(DP_mult_205_n1672), .ZN(DP_mult_205_n1377)
         );
  OAI22_X1 DP_mult_205_U2475 ( .A1(DP_mult_205_n2100), .A2(DP_mult_205_n1680), 
        .B1(DP_mult_205_n1679), .B2(DP_mult_205_n2273), .ZN(DP_mult_205_n1384)
         );
  OAI22_X1 DP_mult_205_U2474 ( .A1(DP_mult_205_n2245), .A2(DP_mult_205_n1674), 
        .B1(DP_mult_205_n1673), .B2(DP_mult_205_n2274), .ZN(DP_mult_205_n1378)
         );
  OAI22_X1 DP_mult_205_U2473 ( .A1(DP_mult_205_n2245), .A2(DP_mult_205_n1676), 
        .B1(DP_mult_205_n1675), .B2(DP_mult_205_n2273), .ZN(DP_mult_205_n1380)
         );
  OAI22_X1 DP_mult_205_U2472 ( .A1(DP_mult_205_n2099), .A2(DP_mult_205_n1675), 
        .B1(DP_mult_205_n2274), .B2(DP_mult_205_n1674), .ZN(DP_mult_205_n1379)
         );
  OAI22_X1 DP_mult_205_U2471 ( .A1(DP_mult_205_n2100), .A2(DP_mult_205_n1672), 
        .B1(DP_mult_205_n1671), .B2(DP_mult_205_n2274), .ZN(DP_mult_205_n1376)
         );
  OAI22_X1 DP_mult_205_U2470 ( .A1(DP_mult_205_n2100), .A2(DP_mult_205_n1677), 
        .B1(DP_mult_205_n2273), .B2(DP_mult_205_n1676), .ZN(DP_mult_205_n1381)
         );
  OAI22_X1 DP_mult_205_U2469 ( .A1(DP_mult_205_n2100), .A2(DP_mult_205_n1679), 
        .B1(DP_mult_205_n2274), .B2(DP_mult_205_n1678), .ZN(DP_mult_205_n1383)
         );
  OAI22_X1 DP_mult_205_U2468 ( .A1(DP_mult_205_n2099), .A2(DP_mult_205_n1671), 
        .B1(DP_mult_205_n2274), .B2(DP_mult_205_n1670), .ZN(DP_mult_205_n1375)
         );
  OAI22_X1 DP_mult_205_U2467 ( .A1(DP_mult_205_n2100), .A2(DP_mult_205_n1670), 
        .B1(DP_mult_205_n1669), .B2(DP_mult_205_n2274), .ZN(DP_mult_205_n1374)
         );
  OAI22_X1 DP_mult_205_U2466 ( .A1(DP_mult_205_n2099), .A2(DP_mult_205_n1669), 
        .B1(DP_mult_205_n2273), .B2(DP_mult_205_n1668), .ZN(DP_mult_205_n1373)
         );
  NAND2_X1 DP_mult_205_U2465 ( .A1(DP_mult_205_n1071), .A2(DP_mult_205_n1084), 
        .ZN(DP_mult_205_n591) );
  NOR2_X1 DP_mult_205_U2464 ( .A1(DP_mult_205_n513), .A2(DP_mult_205_n520), 
        .ZN(DP_mult_205_n511) );
  OAI21_X1 DP_mult_205_U2463 ( .B1(DP_mult_205_n2059), .B2(DP_mult_205_n521), 
        .A(DP_mult_205_n514), .ZN(DP_mult_205_n512) );
  OAI22_X1 DP_mult_205_U2462 ( .A1(DP_mult_205_n2237), .A2(DP_mult_205_n1538), 
        .B1(DP_mult_205_n2260), .B2(DP_mult_205_n1537), .ZN(DP_mult_205_n1247)
         );
  OAI22_X1 DP_mult_205_U2461 ( .A1(DP_mult_205_n2173), .A2(DP_mult_205_n1533), 
        .B1(DP_mult_205_n1532), .B2(DP_mult_205_n2260), .ZN(DP_mult_205_n692)
         );
  OAI22_X1 DP_mult_205_U2460 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1540), 
        .B1(DP_mult_205_n2259), .B2(DP_mult_205_n1539), .ZN(DP_mult_205_n1249)
         );
  OAI22_X1 DP_mult_205_U2459 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1541), 
        .B1(DP_mult_205_n1540), .B2(DP_mult_205_n2260), .ZN(DP_mult_205_n1250)
         );
  OAI22_X1 DP_mult_205_U2458 ( .A1(DP_mult_205_n1556), .A2(DP_mult_205_n2259), 
        .B1(DP_mult_205_n2103), .B2(DP_mult_205_n2321), .ZN(DP_mult_205_n1184)
         );
  OAI22_X1 DP_mult_205_U2457 ( .A1(DP_mult_205_n2237), .A2(DP_mult_205_n1543), 
        .B1(DP_mult_205_n1542), .B2(DP_mult_205_n2260), .ZN(DP_mult_205_n1252)
         );
  OAI22_X1 DP_mult_205_U2456 ( .A1(DP_mult_205_n2103), .A2(DP_mult_205_n1542), 
        .B1(DP_mult_205_n2260), .B2(DP_mult_205_n1541), .ZN(DP_mult_205_n1251)
         );
  OAI22_X1 DP_mult_205_U2455 ( .A1(DP_mult_205_n2173), .A2(DP_mult_205_n1539), 
        .B1(DP_mult_205_n1538), .B2(DP_mult_205_n2259), .ZN(DP_mult_205_n1248)
         );
  OAI22_X1 DP_mult_205_U2454 ( .A1(DP_mult_205_n2237), .A2(DP_mult_205_n1537), 
        .B1(DP_mult_205_n1536), .B2(DP_mult_205_n2260), .ZN(DP_mult_205_n1246)
         );
  OAI22_X1 DP_mult_205_U2453 ( .A1(DP_mult_205_n2173), .A2(DP_mult_205_n1534), 
        .B1(DP_mult_205_n2259), .B2(DP_mult_205_n1533), .ZN(DP_mult_205_n1243)
         );
  OAI22_X1 DP_mult_205_U2452 ( .A1(DP_mult_205_n2237), .A2(DP_mult_205_n1535), 
        .B1(DP_mult_205_n1534), .B2(DP_mult_205_n2259), .ZN(DP_mult_205_n1244)
         );
  OAI22_X1 DP_mult_205_U2451 ( .A1(DP_mult_205_n2237), .A2(DP_mult_205_n1536), 
        .B1(DP_mult_205_n2260), .B2(DP_mult_205_n1535), .ZN(DP_mult_205_n1245)
         );
  NAND2_X1 DP_mult_205_U2450 ( .A1(DP_mult_205_n685), .A2(DP_mult_205_n688), 
        .ZN(DP_mult_205_n369) );
  OAI21_X1 DP_mult_205_U2449 ( .B1(DP_mult_205_n364), .B2(DP_mult_205_n387), 
        .A(DP_mult_205_n365), .ZN(DP_mult_205_n363) );
  NAND2_X1 DP_mult_205_U2448 ( .A1(DP_mult_205_n345), .A2(DP_mult_205_n2197), 
        .ZN(DP_mult_205_n336) );
  INV_X1 DP_mult_205_U2447 ( .A(DP_mult_205_n345), .ZN(DP_mult_205_n343) );
  INV_X1 DP_mult_205_U2446 ( .A(DP_coeffs_fb_int[28]), .ZN(DP_mult_205_n2321)
         );
  OAI22_X1 DP_mult_205_U2445 ( .A1(DP_mult_205_n1781), .A2(DP_mult_205_n2280), 
        .B1(DP_mult_205_n1994), .B2(DP_mult_205_n2222), .ZN(DP_mult_205_n1193)
         );
  XNOR2_X1 DP_mult_205_U2444 ( .A(DP_mult_205_n342), .B(DP_mult_205_n302), 
        .ZN(DP_sw1_coeff_ret1[22]) );
  XNOR2_X1 DP_mult_205_U2443 ( .A(DP_sw1_21_), .B(DP_mult_205_n2298), .ZN(
        DP_mult_205_n1659) );
  XNOR2_X1 DP_mult_205_U2442 ( .A(DP_sw1_13_), .B(DP_mult_205_n2298), .ZN(
        DP_mult_205_n1667) );
  XNOR2_X1 DP_mult_205_U2441 ( .A(DP_sw1_15_), .B(DP_mult_205_n2299), .ZN(
        DP_mult_205_n1665) );
  XNOR2_X1 DP_mult_205_U2440 ( .A(DP_sw1_19_), .B(DP_mult_205_n2299), .ZN(
        DP_mult_205_n1661) );
  XNOR2_X1 DP_mult_205_U2439 ( .A(DP_sw1_11_), .B(DP_mult_205_n2298), .ZN(
        DP_mult_205_n1669) );
  XNOR2_X1 DP_mult_205_U2438 ( .A(DP_sw1_17_), .B(DP_mult_205_n2299), .ZN(
        DP_mult_205_n1663) );
  INV_X1 DP_mult_205_U2437 ( .A(DP_mult_205_n772), .ZN(DP_mult_205_n773) );
  OAI21_X1 DP_mult_205_U2436 ( .B1(DP_mult_205_n2021), .B2(DP_mult_205_n2023), 
        .A(DP_mult_205_n2335), .ZN(DP_mult_205_n1338) );
  NAND2_X1 DP_mult_205_U2435 ( .A1(DP_mult_205_n749), .A2(DP_mult_205_n760), 
        .ZN(DP_mult_205_n439) );
  NOR2_X1 DP_mult_205_U2434 ( .A1(DP_mult_205_n749), .A2(DP_mult_205_n760), 
        .ZN(DP_mult_205_n438) );
  XNOR2_X1 DP_mult_205_U2433 ( .A(DP_sw1_21_), .B(DP_mult_205_n2294), .ZN(
        DP_mult_205_n1684) );
  XNOR2_X1 DP_mult_205_U2432 ( .A(DP_sw1_17_), .B(DP_mult_205_n2294), .ZN(
        DP_mult_205_n1688) );
  XNOR2_X1 DP_mult_205_U2431 ( .A(DP_sw1_17_), .B(DP_mult_205_n2308), .ZN(
        DP_mult_205_n1613) );
  XNOR2_X1 DP_mult_205_U2430 ( .A(DP_sw1_13_), .B(DP_mult_205_n2306), .ZN(
        DP_mult_205_n1617) );
  XNOR2_X1 DP_mult_205_U2429 ( .A(DP_sw1_21_), .B(DP_mult_205_n2306), .ZN(
        DP_mult_205_n1609) );
  XNOR2_X1 DP_mult_205_U2428 ( .A(DP_sw1_15_), .B(DP_mult_205_n2308), .ZN(
        DP_mult_205_n1615) );
  XNOR2_X1 DP_mult_205_U2427 ( .A(DP_sw1_11_), .B(DP_mult_205_n2307), .ZN(
        DP_mult_205_n1619) );
  XNOR2_X1 DP_mult_205_U2426 ( .A(DP_sw1_19_), .B(DP_mult_205_n2308), .ZN(
        DP_mult_205_n1611) );
  OAI21_X1 DP_mult_205_U2425 ( .B1(DP_mult_205_n1972), .B2(DP_mult_205_n2205), 
        .A(DP_mult_205_n2337), .ZN(DP_mult_205_n1290) );
  NOR2_X1 DP_mult_205_U2424 ( .A1(DP_mult_205_n420), .A2(DP_mult_205_n347), 
        .ZN(DP_mult_205_n345) );
  NAND2_X1 DP_mult_205_U2423 ( .A1(DP_mult_205_n332), .A2(DP_mult_205_n1959), 
        .ZN(DP_mult_205_n326) );
  INV_X1 DP_mult_205_U2422 ( .A(DP_mult_205_n474), .ZN(DP_mult_205_n472) );
  NAND2_X1 DP_mult_205_U2421 ( .A1(DP_mult_205_n2182), .A2(DP_mult_205_n474), 
        .ZN(DP_mult_205_n314) );
  AOI21_X1 DP_mult_205_U2420 ( .B1(DP_mult_205_n401), .B2(DP_mult_205_n2191), 
        .A(DP_mult_205_n394), .ZN(DP_mult_205_n390) );
  OAI21_X1 DP_mult_205_U2419 ( .B1(DP_mult_205_n390), .B2(DP_mult_205_n384), 
        .A(DP_mult_205_n387), .ZN(DP_mult_205_n383) );
  OAI21_X1 DP_mult_205_U2418 ( .B1(DP_mult_205_n503), .B2(DP_mult_205_n495), 
        .A(DP_mult_205_n496), .ZN(DP_mult_205_n490) );
  XNOR2_X1 DP_mult_205_U2417 ( .A(DP_mult_205_n475), .B(DP_mult_205_n314), 
        .ZN(DP_sw1_coeff_ret1[10]) );
  NAND2_X1 DP_mult_205_U2416 ( .A1(DP_mult_205_n525), .A2(DP_mult_205_n2036), 
        .ZN(DP_mult_205_n505) );
  NAND2_X1 DP_mult_205_U2415 ( .A1(DP_mult_205_n2168), .A2(DP_mult_205_n2169), 
        .ZN(DP_mult_205_n516) );
  OAI22_X1 DP_mult_205_U2414 ( .A1(DP_mult_205_n2242), .A2(DP_mult_205_n1622), 
        .B1(DP_mult_205_n1621), .B2(DP_mult_205_n2268), .ZN(DP_mult_205_n1328)
         );
  OAI22_X1 DP_mult_205_U2413 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1627), 
        .B1(DP_mult_205_n2267), .B2(DP_mult_205_n1626), .ZN(DP_mult_205_n1333)
         );
  AOI21_X1 DP_mult_205_U2412 ( .B1(DP_mult_205_n2229), .B2(DP_mult_205_n2169), 
        .A(DP_mult_205_n2140), .ZN(DP_mult_205_n517) );
  INV_X1 DP_mult_205_U2411 ( .A(DP_mult_205_n2229), .ZN(DP_mult_205_n524) );
  AOI21_X1 DP_mult_205_U2410 ( .B1(DP_mult_205_n2182), .B2(DP_mult_205_n483), 
        .A(DP_mult_205_n472), .ZN(DP_mult_205_n468) );
  NAND2_X1 DP_mult_205_U2409 ( .A1(DP_mult_205_n666), .A2(DP_mult_205_n2182), 
        .ZN(DP_mult_205_n467) );
  OAI22_X1 DP_mult_205_U2408 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1625), 
        .B1(DP_mult_205_n2268), .B2(DP_mult_205_n1624), .ZN(DP_mult_205_n1331)
         );
  OAI22_X1 DP_mult_205_U2407 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1626), 
        .B1(DP_mult_205_n1625), .B2(DP_mult_205_n2267), .ZN(DP_mult_205_n1332)
         );
  OAI22_X1 DP_mult_205_U2406 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1623), 
        .B1(DP_mult_205_n2268), .B2(DP_mult_205_n1622), .ZN(DP_mult_205_n1329)
         );
  OAI22_X1 DP_mult_205_U2405 ( .A1(DP_mult_205_n1995), .A2(DP_mult_205_n1621), 
        .B1(DP_mult_205_n2268), .B2(DP_mult_205_n1620), .ZN(DP_mult_205_n1327)
         );
  OAI22_X1 DP_mult_205_U2404 ( .A1(DP_mult_205_n1995), .A2(DP_mult_205_n1624), 
        .B1(DP_mult_205_n1623), .B2(DP_mult_205_n2267), .ZN(DP_mult_205_n1330)
         );
  OAI22_X1 DP_mult_205_U2403 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1629), 
        .B1(DP_mult_205_n2268), .B2(DP_mult_205_n1628), .ZN(DP_mult_205_n1335)
         );
  OAI22_X1 DP_mult_205_U2402 ( .A1(DP_mult_205_n1995), .A2(DP_mult_205_n1619), 
        .B1(DP_mult_205_n2267), .B2(DP_mult_205_n1618), .ZN(DP_mult_205_n1325)
         );
  OAI22_X1 DP_mult_205_U2401 ( .A1(DP_mult_205_n2130), .A2(DP_mult_205_n1620), 
        .B1(DP_mult_205_n1619), .B2(DP_mult_205_n2267), .ZN(DP_mult_205_n1326)
         );
  OAI22_X1 DP_mult_205_U2400 ( .A1(DP_mult_205_n1995), .A2(DP_mult_205_n1630), 
        .B1(DP_mult_205_n1629), .B2(DP_mult_205_n2268), .ZN(DP_mult_205_n1336)
         );
  NAND2_X1 DP_mult_205_U2399 ( .A1(DP_mult_205_n1813), .A2(DP_mult_205_n2272), 
        .ZN(DP_mult_205_n283) );
  OAI21_X1 DP_mult_205_U2398 ( .B1(DP_mult_205_n492), .B2(DP_mult_205_n467), 
        .A(DP_mult_205_n468), .ZN(DP_mult_205_n466) );
  XNOR2_X1 DP_mult_205_U2397 ( .A(DP_mult_205_n462), .B(DP_mult_205_n313), 
        .ZN(DP_sw1_coeff_ret1[11]) );
  NOR2_X1 DP_mult_205_U2396 ( .A1(DP_mult_205_n737), .A2(DP_mult_205_n748), 
        .ZN(DP_mult_205_n435) );
  AOI21_X1 DP_mult_205_U2395 ( .B1(DP_mult_205_n508), .B2(DP_mult_205_n2167), 
        .A(DP_mult_205_n2223), .ZN(DP_mult_205_n488) );
  AOI21_X1 DP_mult_205_U2394 ( .B1(DP_mult_205_n508), .B2(DP_mult_205_n668), 
        .A(DP_mult_205_n501), .ZN(DP_mult_205_n499) );
  AOI21_X1 DP_mult_205_U2393 ( .B1(DP_mult_205_n508), .B2(DP_mult_205_n465), 
        .A(DP_mult_205_n466), .ZN(DP_mult_205_n464) );
  AOI21_X1 DP_mult_205_U2392 ( .B1(DP_mult_205_n508), .B2(DP_mult_205_n478), 
        .A(DP_mult_205_n479), .ZN(DP_mult_205_n477) );
  XNOR2_X1 DP_mult_205_U2391 ( .A(DP_mult_205_n486), .B(DP_mult_205_n315), 
        .ZN(DP_sw1_coeff_ret1[9]) );
  NOR2_X1 DP_mult_205_U2390 ( .A1(DP_mult_205_n505), .A2(DP_mult_205_n452), 
        .ZN(DP_mult_205_n450) );
  INV_X1 DP_mult_205_U2389 ( .A(DP_mult_205_n451), .ZN(DP_mult_205_n2232) );
  NAND2_X1 DP_mult_205_U2388 ( .A1(DP_mult_205_n537), .A2(DP_mult_205_n450), 
        .ZN(DP_mult_205_n2231) );
  OAI21_X1 DP_mult_205_U2387 ( .B1(DP_mult_205_n428), .B2(DP_mult_205_n436), 
        .A(DP_mult_205_n429), .ZN(DP_mult_205_n427) );
  NOR2_X1 DP_mult_205_U2386 ( .A1(DP_mult_205_n727), .A2(DP_mult_205_n736), 
        .ZN(DP_mult_205_n428) );
  XNOR2_X1 DP_mult_205_U2385 ( .A(DP_mult_205_n522), .B(DP_mult_205_n319), 
        .ZN(DP_sw1_coeff_ret1[5]) );
  OAI21_X1 DP_mult_205_U2384 ( .B1(DP_mult_205_n2252), .B2(DP_mult_205_n2134), 
        .A(DP_mult_205_n2331), .ZN(DP_mult_205_n1434) );
  NAND2_X1 DP_mult_205_U2383 ( .A1(DP_mult_205_n1165), .A2(DP_mult_205_n1170), 
        .ZN(DP_mult_205_n632) );
  XNOR2_X1 DP_mult_205_U2382 ( .A(DP_mult_205_n515), .B(DP_mult_205_n318), 
        .ZN(DP_sw1_coeff_ret1[6]) );
  OAI21_X1 DP_mult_205_U2381 ( .B1(DP_mult_205_n558), .B2(DP_mult_205_n564), 
        .A(DP_mult_205_n559), .ZN(DP_mult_205_n553) );
  INV_X1 DP_mult_205_U2380 ( .A(DP_mult_205_n558), .ZN(DP_mult_205_n675) );
  OAI21_X1 DP_mult_205_U2379 ( .B1(DP_mult_205_n2170), .B2(DP_mult_205_n535), 
        .A(DP_mult_205_n532), .ZN(DP_mult_205_n526) );
  OAI21_X1 DP_mult_205_U2378 ( .B1(DP_mult_205_n535), .B2(DP_mult_205_n2058), 
        .A(DP_mult_205_n2080), .ZN(DP_mult_205_n2229) );
  NAND2_X1 DP_mult_205_U2377 ( .A1(DP_mult_205_n919), .A2(DP_mult_205_n940), 
        .ZN(DP_mult_205_n543) );
  INV_X1 DP_mult_205_U2376 ( .A(DP_mult_205_n706), .ZN(DP_mult_205_n707) );
  NAND2_X1 DP_mult_205_U2375 ( .A1(DP_mult_205_n701), .A2(DP_mult_205_n708), 
        .ZN(DP_mult_205_n396) );
  OAI21_X1 DP_mult_205_U2374 ( .B1(DP_mult_205_n2250), .B2(DP_mult_205_n2202), 
        .A(DP_mult_205_n2332), .ZN(DP_mult_205_n1410) );
  NAND2_X1 DP_mult_205_U2373 ( .A1(DP_mult_205_n1171), .A2(DP_mult_205_n1174), 
        .ZN(DP_mult_205_n634) );
  NOR2_X1 DP_mult_205_U2372 ( .A1(DP_mult_205_n1171), .A2(DP_mult_205_n1174), 
        .ZN(DP_mult_205_n633) );
  INV_X1 DP_mult_205_U2371 ( .A(DP_mult_205_n382), .ZN(DP_mult_205_n380) );
  OR2_X1 DP_mult_205_U2370 ( .A1(DP_mult_205_n727), .A2(DP_mult_205_n736), 
        .ZN(DP_mult_205_n2228) );
  OAI21_X1 DP_mult_205_U2369 ( .B1(DP_mult_205_n572), .B2(DP_mult_205_n569), 
        .A(DP_mult_205_n570), .ZN(DP_mult_205_n568) );
  NOR2_X1 DP_mult_205_U2368 ( .A1(DP_mult_205_n876), .A2(DP_mult_205_n1929), 
        .ZN(DP_mult_205_n520) );
  NAND2_X1 DP_mult_205_U2367 ( .A1(DP_mult_205_n507), .A2(DP_mult_205_n668), 
        .ZN(DP_mult_205_n498) );
  NAND2_X1 DP_mult_205_U2366 ( .A1(DP_mult_205_n465), .A2(DP_mult_205_n507), 
        .ZN(DP_mult_205_n463) );
  NAND2_X1 DP_mult_205_U2365 ( .A1(DP_mult_205_n478), .A2(DP_mult_205_n507), 
        .ZN(DP_mult_205_n476) );
  NAND2_X1 DP_mult_205_U2364 ( .A1(DP_mult_205_n507), .A2(DP_mult_205_n2167), 
        .ZN(DP_mult_205_n487) );
  AOI21_X1 DP_mult_205_U2363 ( .B1(DP_mult_205_n472), .B2(DP_mult_205_n2183), 
        .A(DP_mult_205_n459), .ZN(DP_mult_205_n457) );
  NOR2_X1 DP_mult_205_U2362 ( .A1(DP_mult_205_n456), .A2(DP_mult_205_n480), 
        .ZN(DP_mult_205_n454) );
  NOR2_X1 DP_mult_205_U2361 ( .A1(DP_mult_205_n542), .A2(DP_mult_205_n547), 
        .ZN(DP_mult_205_n540) );
  OAI22_X1 DP_mult_205_U2360 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1770), 
        .B1(DP_mult_205_n1769), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1471)
         );
  INV_X1 DP_mult_205_U2359 ( .A(DP_mult_205_n1941), .ZN(DP_mult_205_n508) );
  NAND2_X1 DP_mult_205_U2358 ( .A1(DP_mult_205_n1003), .A2(DP_mult_205_n1020), 
        .ZN(DP_mult_205_n570) );
  NOR2_X1 DP_mult_205_U2357 ( .A1(DP_mult_205_n1003), .A2(DP_mult_205_n1020), 
        .ZN(DP_mult_205_n569) );
  NOR2_X1 DP_mult_205_U2356 ( .A1(DP_mult_205_n919), .A2(DP_mult_205_n940), 
        .ZN(DP_mult_205_n542) );
  NOR2_X1 DP_mult_205_U2355 ( .A1(DP_mult_205_n919), .A2(DP_mult_205_n940), 
        .ZN(DP_mult_205_n2227) );
  NAND2_X1 DP_mult_205_U2354 ( .A1(DP_mult_205_n426), .A2(DP_mult_205_n663), 
        .ZN(DP_mult_205_n420) );
  NOR2_X1 DP_mult_205_U2353 ( .A1(DP_mult_205_n435), .A2(DP_mult_205_n428), 
        .ZN(DP_mult_205_n426) );
  OAI21_X1 DP_mult_205_U2352 ( .B1(DP_mult_205_n631), .B2(DP_mult_205_n634), 
        .A(DP_mult_205_n632), .ZN(DP_mult_205_n630) );
  NOR2_X1 DP_mult_205_U2351 ( .A1(DP_mult_205_n633), .A2(DP_mult_205_n631), 
        .ZN(DP_mult_205_n629) );
  INV_X1 DP_mult_205_U2350 ( .A(DP_mult_205_n461), .ZN(DP_mult_205_n459) );
  OAI21_X1 DP_mult_205_U2349 ( .B1(DP_mult_205_n456), .B2(DP_mult_205_n481), 
        .A(DP_mult_205_n457), .ZN(DP_mult_205_n455) );
  OR2_X1 DP_mult_205_U2348 ( .A1(DP_mult_205_n940), .A2(DP_mult_205_n1997), 
        .ZN(DP_mult_205_n2226) );
  NAND2_X1 DP_mult_205_U2347 ( .A1(DP_mult_205_n821), .A2(DP_mult_205_n838), 
        .ZN(DP_mult_205_n503) );
  NOR2_X1 DP_mult_205_U2346 ( .A1(DP_mult_205_n821), .A2(DP_mult_205_n838), 
        .ZN(DP_mult_205_n502) );
  INV_X1 DP_mult_205_U2345 ( .A(DP_mult_205_n2167), .ZN(DP_mult_205_n491) );
  INV_X1 DP_mult_205_U2344 ( .A(DP_coeffs_fb_int[26]), .ZN(DP_mult_205_n2325)
         );
  INV_X1 DP_mult_205_U2343 ( .A(DP_mult_205_n2317), .ZN(DP_mult_205_n2315) );
  NOR2_X1 DP_mult_205_U2342 ( .A1(DP_mult_205_n571), .A2(DP_mult_205_n1993), 
        .ZN(DP_mult_205_n567) );
  INV_X1 DP_mult_205_U2341 ( .A(DP_mult_205_n2081), .ZN(DP_mult_205_n492) );
  INV_X1 DP_mult_205_U2340 ( .A(DP_mult_205_n503), .ZN(DP_mult_205_n501) );
  NAND2_X1 DP_mult_205_U2339 ( .A1(DP_mult_205_n668), .A2(DP_mult_205_n503), 
        .ZN(DP_mult_205_n317) );
  NOR2_X1 DP_mult_205_U2338 ( .A1(DP_mult_205_n1181), .A2(DP_mult_205_n1192), 
        .ZN(DP_mult_205_n644) );
  NAND2_X1 DP_mult_205_U2337 ( .A1(DP_mult_205_n1181), .A2(DP_mult_205_n1192), 
        .ZN(DP_mult_205_n645) );
  NAND2_X1 DP_mult_205_U2336 ( .A1(DP_mult_205_n2192), .A2(DP_mult_205_n2189), 
        .ZN(DP_mult_205_n599) );
  OAI21_X1 DP_mult_205_U2335 ( .B1(DP_mult_205_n405), .B2(DP_mult_205_n360), 
        .A(DP_mult_205_n361), .ZN(DP_mult_205_n359) );
  AOI21_X1 DP_mult_205_U2334 ( .B1(DP_mult_205_n359), .B2(DP_mult_205_n2196), 
        .A(DP_mult_205_n350), .ZN(DP_mult_205_n348) );
  NOR2_X1 DP_mult_205_U2333 ( .A1(DP_mult_205_n805), .A2(DP_mult_205_n820), 
        .ZN(DP_mult_205_n495) );
  AOI21_X1 DP_mult_205_U2332 ( .B1(DP_mult_205_n2184), .B2(DP_mult_205_n1946), 
        .A(DP_mult_205_n1956), .ZN(DP_mult_205_n572) );
  NAND2_X1 DP_mult_205_U2331 ( .A1(DP_mult_205_n2184), .A2(DP_mult_205_n2185), 
        .ZN(DP_mult_205_n571) );
  NOR2_X1 DP_mult_205_U2330 ( .A1(DP_mult_205_n1085), .A2(DP_mult_205_n1098), 
        .ZN(DP_mult_205_n592) );
  NAND2_X1 DP_mult_205_U2329 ( .A1(DP_mult_205_n1085), .A2(DP_mult_205_n1098), 
        .ZN(DP_mult_205_n593) );
  OAI21_X1 DP_mult_205_U2328 ( .B1(DP_mult_205_n590), .B2(DP_mult_205_n593), 
        .A(DP_mult_205_n591), .ZN(DP_mult_205_n589) );
  NOR2_X1 DP_mult_205_U2327 ( .A1(DP_mult_205_n590), .A2(DP_mult_205_n592), 
        .ZN(DP_mult_205_n588) );
  NOR2_X1 DP_mult_205_U2326 ( .A1(DP_mult_205_n1071), .A2(DP_mult_205_n1084), 
        .ZN(DP_mult_205_n590) );
  INV_X1 DP_mult_205_U2325 ( .A(DP_mult_205_n502), .ZN(DP_mult_205_n668) );
  NOR2_X1 DP_mult_205_U2324 ( .A1(DP_mult_205_n491), .A2(DP_mult_205_n467), 
        .ZN(DP_mult_205_n465) );
  NOR2_X1 DP_mult_205_U2323 ( .A1(DP_mult_205_n491), .A2(DP_mult_205_n480), 
        .ZN(DP_mult_205_n478) );
  AOI21_X1 DP_mult_205_U2322 ( .B1(DP_mult_205_n526), .B2(DP_mult_205_n511), 
        .A(DP_mult_205_n512), .ZN(DP_mult_205_n506) );
  INV_X1 DP_mult_205_U2321 ( .A(DP_mult_205_n508), .ZN(DP_mult_205_n2225) );
  NAND2_X1 DP_mult_205_U2320 ( .A1(DP_mult_205_n983), .A2(DP_mult_205_n1002), 
        .ZN(DP_mult_205_n564) );
  NOR2_X1 DP_mult_205_U2319 ( .A1(DP_mult_205_n983), .A2(DP_mult_205_n1002), 
        .ZN(DP_mult_205_n563) );
  INV_X1 DP_mult_205_U2318 ( .A(DP_mult_205_n553), .ZN(DP_mult_205_n555) );
  AOI21_X1 DP_mult_205_U2317 ( .B1(DP_mult_205_n565), .B2(DP_mult_205_n2105), 
        .A(DP_mult_205_n1932), .ZN(DP_mult_205_n551) );
  OR2_X1 DP_mult_205_U2316 ( .A1(DP_mult_205_n805), .A2(DP_mult_205_n1936), 
        .ZN(DP_mult_205_n2224) );
  CLKBUF_X1 DP_mult_205_U2315 ( .A(DP_mult_205_n2081), .Z(DP_mult_205_n2223)
         );
  INV_X1 DP_mult_205_U2314 ( .A(DP_mult_205_n2284), .ZN(DP_mult_205_n2222) );
  INV_X1 DP_mult_205_U2313 ( .A(DP_mult_205_n1989), .ZN(DP_mult_205_n565) );
  NAND2_X1 DP_mult_205_U2312 ( .A1(DP_mult_205_n897), .A2(DP_mult_205_n918), 
        .ZN(DP_mult_205_n535) );
  NAND2_X1 DP_mult_205_U2311 ( .A1(DP_mult_205_n2182), .A2(DP_mult_205_n2183), 
        .ZN(DP_mult_205_n456) );
  NOR2_X1 DP_mult_205_U2310 ( .A1(DP_mult_205_n420), .A2(DP_mult_205_n402), 
        .ZN(DP_mult_205_n400) );
  NAND2_X1 DP_mult_205_U2309 ( .A1(DP_mult_205_n1808), .A2(DP_mult_205_n2258), 
        .ZN(DP_mult_205_n293) );
  NAND2_X1 DP_mult_205_U2308 ( .A1(DP_mult_205_n839), .A2(DP_mult_205_n856), 
        .ZN(DP_mult_205_n514) );
  OAI22_X1 DP_mult_205_U2307 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1711), 
        .B1(DP_mult_205_n2276), .B2(DP_mult_205_n1710), .ZN(DP_mult_205_n1413)
         );
  OAI22_X1 DP_mult_205_U2306 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1709), 
        .B1(DP_mult_205_n2276), .B2(DP_mult_205_n1708), .ZN(DP_mult_205_n1411)
         );
  OAI22_X1 DP_mult_205_U2305 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1715), 
        .B1(DP_mult_205_n2276), .B2(DP_mult_205_n1714), .ZN(DP_mult_205_n1417)
         );
  OAI22_X1 DP_mult_205_U2304 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1713), 
        .B1(DP_mult_205_n2276), .B2(DP_mult_205_n1712), .ZN(DP_mult_205_n1415)
         );
  OAI22_X1 DP_mult_205_U2303 ( .A1(DP_mult_205_n1988), .A2(DP_mult_205_n1717), 
        .B1(DP_mult_205_n2042), .B2(DP_mult_205_n1716), .ZN(DP_mult_205_n1419)
         );
  NAND2_X1 DP_mult_205_U2302 ( .A1(DP_mult_205_n1099), .A2(DP_mult_205_n1110), 
        .ZN(DP_mult_205_n598) );
  NAND2_X1 DP_mult_205_U2301 ( .A1(DP_mult_205_n941), .A2(DP_mult_205_n962), 
        .ZN(DP_mult_205_n550) );
  NOR2_X1 DP_mult_205_U2300 ( .A1(DP_mult_205_n554), .A2(DP_mult_205_n2098), 
        .ZN(DP_mult_205_n545) );
  OAI21_X1 DP_mult_205_U2299 ( .B1(DP_mult_205_n555), .B2(DP_mult_205_n2074), 
        .A(DP_mult_205_n2045), .ZN(DP_mult_205_n546) );
  NOR2_X1 DP_mult_205_U2298 ( .A1(DP_mult_205_n495), .A2(DP_mult_205_n502), 
        .ZN(DP_mult_205_n489) );
  NOR2_X1 DP_mult_205_U2297 ( .A1(DP_mult_205_n789), .A2(DP_mult_205_n804), 
        .ZN(DP_mult_205_n480) );
  NAND3_X1 DP_mult_205_U2296 ( .A1(DP_mult_205_n2218), .A2(DP_mult_205_n2219), 
        .A3(DP_mult_205_n2220), .ZN(DP_mult_205_n804) );
  NAND2_X1 DP_mult_205_U2295 ( .A1(DP_mult_205_n807), .A2(DP_mult_205_n809), 
        .ZN(DP_mult_205_n2220) );
  NAND2_X1 DP_mult_205_U2294 ( .A1(DP_mult_205_n822), .A2(DP_mult_205_n809), 
        .ZN(DP_mult_205_n2219) );
  NAND2_X1 DP_mult_205_U2293 ( .A1(DP_mult_205_n822), .A2(DP_mult_205_n807), 
        .ZN(DP_mult_205_n2218) );
  INV_X1 DP_mult_205_U2292 ( .A(DP_mult_205_n505), .ZN(DP_mult_205_n507) );
  NAND2_X1 DP_mult_205_U2291 ( .A1(DP_mult_205_n1159), .A2(DP_mult_205_n1161), 
        .ZN(DP_mult_205_n627) );
  NOR2_X1 DP_mult_205_U2290 ( .A1(DP_mult_205_n1159), .A2(DP_mult_205_n1161), 
        .ZN(DP_mult_205_n626) );
  NAND2_X1 DP_mult_205_U2289 ( .A1(DP_mult_205_n400), .A2(DP_mult_205_n2191), 
        .ZN(DP_mult_205_n389) );
  INV_X1 DP_mult_205_U2288 ( .A(DP_mult_205_n400), .ZN(DP_mult_205_n398) );
  OR2_X1 DP_mult_205_U2287 ( .A1(DP_mult_205_n897), .A2(DP_mult_205_n918), 
        .ZN(DP_mult_205_n2217) );
  NAND3_X1 DP_mult_205_U2286 ( .A1(DP_mult_205_n2214), .A2(DP_mult_205_n2215), 
        .A3(DP_mult_205_n2216), .ZN(DP_mult_205_n898) );
  NAND2_X1 DP_mult_205_U2285 ( .A1(DP_mult_205_n903), .A2(DP_mult_205_n924), 
        .ZN(DP_mult_205_n2216) );
  NAND2_X1 DP_mult_205_U2284 ( .A1(DP_mult_205_n922), .A2(DP_mult_205_n924), 
        .ZN(DP_mult_205_n2215) );
  NAND2_X1 DP_mult_205_U2283 ( .A1(DP_mult_205_n2019), .A2(DP_mult_205_n903), 
        .ZN(DP_mult_205_n2214) );
  XNOR2_X1 DP_mult_205_U2282 ( .A(DP_sw1_7_), .B(DP_mult_205_n2291), .ZN(
        DP_mult_205_n1723) );
  XNOR2_X1 DP_mult_205_U2281 ( .A(DP_mult_205_n2290), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1724) );
  NAND2_X1 DP_mult_205_U2280 ( .A1(DP_mult_205_n2212), .A2(DP_mult_205_n2213), 
        .ZN(DP_mult_205_n1426) );
  OR2_X1 DP_mult_205_U2279 ( .A1(DP_mult_205_n1723), .A2(DP_mult_205_n2043), 
        .ZN(DP_mult_205_n2213) );
  OR2_X1 DP_mult_205_U2278 ( .A1(DP_mult_205_n2249), .A2(DP_mult_205_n1724), 
        .ZN(DP_mult_205_n2212) );
  NAND3_X1 DP_mult_205_U2277 ( .A1(DP_mult_205_n2209), .A2(DP_mult_205_n2210), 
        .A3(DP_mult_205_n2211), .ZN(DP_mult_205_n1110) );
  NAND2_X1 DP_mult_205_U2276 ( .A1(DP_mult_205_n1124), .A2(DP_mult_205_n1115), 
        .ZN(DP_mult_205_n2211) );
  NAND2_X1 DP_mult_205_U2275 ( .A1(DP_mult_205_n1113), .A2(DP_mult_205_n1115), 
        .ZN(DP_mult_205_n2210) );
  NAND2_X1 DP_mult_205_U2274 ( .A1(DP_mult_205_n1113), .A2(DP_mult_205_n1124), 
        .ZN(DP_mult_205_n2209) );
  INV_X1 DP_mult_205_U2273 ( .A(DP_mult_205_n2093), .ZN(DP_mult_205_n2247) );
  OAI22_X1 DP_mult_205_U2272 ( .A1(DP_mult_205_n2177), .A2(DP_mult_205_n1490), 
        .B1(DP_mult_205_n2255), .B2(DP_mult_205_n1489), .ZN(DP_mult_205_n1201)
         );
  OAI22_X1 DP_mult_205_U2271 ( .A1(DP_mult_205_n2233), .A2(DP_mult_205_n1492), 
        .B1(DP_mult_205_n2254), .B2(DP_mult_205_n1491), .ZN(DP_mult_205_n1203)
         );
  OAI22_X1 DP_mult_205_U2270 ( .A1(DP_mult_205_n2177), .A2(DP_mult_205_n1486), 
        .B1(DP_mult_205_n2254), .B2(DP_mult_205_n1485), .ZN(DP_mult_205_n1197)
         );
  OAI22_X1 DP_mult_205_U2269 ( .A1(DP_mult_205_n2178), .A2(DP_mult_205_n1488), 
        .B1(DP_mult_205_n2255), .B2(DP_mult_205_n1487), .ZN(DP_mult_205_n1199)
         );
  OAI22_X1 DP_mult_205_U2268 ( .A1(DP_mult_205_n2178), .A2(DP_mult_205_n1484), 
        .B1(DP_mult_205_n2255), .B2(DP_mult_205_n1483), .ZN(DP_mult_205_n1195)
         );
  NAND2_X1 DP_mult_205_U2267 ( .A1(DP_mult_205_n2169), .A2(DP_mult_205_n521), 
        .ZN(DP_mult_205_n319) );
  AOI21_X1 DP_mult_205_U2266 ( .B1(DP_mult_205_n565), .B2(DP_mult_205_n545), 
        .A(DP_mult_205_n546), .ZN(DP_mult_205_n544) );
  AOI21_X1 DP_mult_205_U2265 ( .B1(DP_mult_205_n565), .B2(DP_mult_205_n561), 
        .A(DP_mult_205_n562), .ZN(DP_mult_205_n560) );
  INV_X1 DP_mult_205_U2264 ( .A(DP_mult_205_n874), .ZN(DP_mult_205_n875) );
  NOR2_X1 DP_mult_205_U2263 ( .A1(DP_mult_205_n384), .A2(DP_mult_205_n364), 
        .ZN(DP_mult_205_n362) );
  AOI21_X1 DP_mult_205_U2262 ( .B1(DP_mult_205_n362), .B2(DP_mult_205_n394), 
        .A(DP_mult_205_n363), .ZN(DP_mult_205_n361) );
  NAND2_X1 DP_mult_205_U2261 ( .A1(DP_mult_205_n362), .A2(DP_mult_205_n2191), 
        .ZN(DP_mult_205_n360) );
  NAND2_X1 DP_mult_205_U2260 ( .A1(DP_mult_205_n356), .A2(DP_mult_205_n2196), 
        .ZN(DP_mult_205_n347) );
  OAI21_X1 DP_mult_205_U2259 ( .B1(DP_mult_205_n2102), .B2(DP_mult_205_n1992), 
        .A(DP_mult_205_n2338), .ZN(DP_mult_205_n1266) );
  OAI21_X1 DP_mult_205_U2258 ( .B1(DP_mult_205_n1940), .B2(DP_mult_205_n2107), 
        .A(DP_mult_205_n2341), .ZN(DP_mult_205_n1194) );
  INV_X1 DP_mult_205_U2257 ( .A(DP_coeffs_fb_int[44]), .ZN(DP_mult_205_n2289)
         );
  XNOR2_X1 DP_mult_205_U2256 ( .A(DP_sw1_23_), .B(DP_mult_205_n2326), .ZN(
        DP_mult_205_n1482) );
  XNOR2_X1 DP_mult_205_U2255 ( .A(DP_mult_205_n448), .B(DP_mult_205_n312), 
        .ZN(DP_sw1_coeff_ret1[12]) );
  NAND2_X1 DP_mult_205_U2254 ( .A1(DP_mult_205_n2183), .A2(DP_mult_205_n461), 
        .ZN(DP_mult_205_n313) );
  NAND2_X1 DP_mult_205_U2253 ( .A1(DP_mult_205_n2069), .A2(DP_mult_205_n2080), 
        .ZN(DP_mult_205_n320) );
  XNOR2_X1 DP_mult_205_U2252 ( .A(DP_mult_205_n504), .B(DP_mult_205_n317), 
        .ZN(DP_sw1_coeff_ret1[7]) );
  INV_X1 DP_mult_205_U2251 ( .A(DP_coeffs_fb_int[47]), .ZN(DP_mult_205_n251)
         );
  XNOR2_X1 DP_mult_205_U2250 ( .A(DP_mult_205_n2311), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1605) );
  XNOR2_X1 DP_mult_205_U2249 ( .A(DP_mult_205_n2288), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1755) );
  OAI22_X1 DP_mult_205_U2248 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1778), 
        .B1(DP_mult_205_n1777), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1479)
         );
  XNOR2_X1 DP_mult_205_U2247 ( .A(DP_mult_205_n2285), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1780) );
  OAI22_X1 DP_mult_205_U2246 ( .A1(DP_mult_205_n1994), .A2(DP_mult_205_n1780), 
        .B1(DP_mult_205_n1779), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1481)
         );
  INV_X1 DP_mult_205_U2245 ( .A(DP_mult_205_n293), .ZN(DP_mult_205_n2238) );
  INV_X1 DP_mult_205_U2244 ( .A(DP_mult_205_n279), .ZN(DP_mult_205_n2250) );
  INV_X1 DP_mult_205_U2243 ( .A(DP_mult_205_n277), .ZN(DP_mult_205_n2252) );
  XNOR2_X1 DP_mult_205_U2242 ( .A(DP_mult_205_n2320), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1555) );
  XNOR2_X1 DP_mult_205_U2241 ( .A(DP_mult_205_n2308), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1630) );
  NAND2_X1 DP_mult_205_U2240 ( .A1(DP_mult_205_n2224), .A2(DP_mult_205_n496), 
        .ZN(DP_mult_205_n316) );
  XNOR2_X1 DP_mult_205_U2239 ( .A(DP_mult_205_n497), .B(DP_mult_205_n316), 
        .ZN(DP_sw1_coeff_ret1[8]) );
  INV_X1 DP_mult_205_U2238 ( .A(DP_mult_205_n283), .ZN(DP_mult_205_n2246) );
  INV_X1 DP_mult_205_U2237 ( .A(DP_mult_205_n287), .ZN(DP_mult_205_n2243) );
  INV_X1 DP_mult_205_U2236 ( .A(DP_mult_205_n1757), .ZN(DP_mult_205_n2330) );
  OAI21_X1 DP_mult_205_U2235 ( .B1(DP_coeffs_fb_int[47]), .B2(
        DP_mult_205_n2082), .A(DP_mult_205_n2330), .ZN(DP_mult_205_n1458) );
  NAND2_X1 DP_mult_205_U2234 ( .A1(DP_mult_205_n666), .A2(DP_mult_205_n481), 
        .ZN(DP_mult_205_n315) );
  NAND2_X1 DP_mult_205_U2233 ( .A1(DP_mult_205_n2166), .A2(DP_mult_205_n1975), 
        .ZN(DP_mult_205_n318) );
  INV_X1 DP_mult_205_U2232 ( .A(DP_mult_205_n259), .ZN(DP_mult_205_n2275) );
  INV_X1 DP_mult_205_U2231 ( .A(DP_coeffs_fb_int[38]), .ZN(DP_mult_205_n2301)
         );
  INV_X1 DP_mult_205_U2230 ( .A(DP_coeffs_fb_int[36]), .ZN(DP_mult_205_n2305)
         );
  INV_X1 DP_mult_205_U2229 ( .A(DP_coeffs_fb_int[40]), .ZN(DP_mult_205_n2297)
         );
  INV_X1 DP_mult_205_U2228 ( .A(DP_coeffs_fb_int[24]), .ZN(DP_mult_205_n2328)
         );
  XNOR2_X1 DP_mult_205_U2227 ( .A(DP_sw1_21_), .B(DP_mult_205_n2326), .ZN(
        DP_mult_205_n1484) );
  XNOR2_X1 DP_mult_205_U2226 ( .A(DP_sw1_19_), .B(DP_mult_205_n2326), .ZN(
        DP_mult_205_n1486) );
  XNOR2_X1 DP_mult_205_U2225 ( .A(DP_sw1_15_), .B(DP_mult_205_n2326), .ZN(
        DP_mult_205_n1490) );
  XNOR2_X1 DP_mult_205_U2224 ( .A(DP_sw1_17_), .B(DP_mult_205_n2326), .ZN(
        DP_mult_205_n1488) );
  XNOR2_X1 DP_mult_205_U2223 ( .A(DP_sw1_11_), .B(DP_mult_205_n2326), .ZN(
        DP_mult_205_n1494) );
  XNOR2_X1 DP_mult_205_U2222 ( .A(DP_sw1_13_), .B(DP_mult_205_n2326), .ZN(
        DP_mult_205_n1492) );
  XNOR2_X1 DP_mult_205_U2221 ( .A(DP_mult_205_n2314), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1580) );
  XOR2_X1 DP_mult_205_U2220 ( .A(DP_coeffs_fb_int[31]), .B(
        DP_coeffs_fb_int[32]), .Z(DP_mult_205_n2199) );
  XNOR2_X1 DP_mult_205_U2219 ( .A(DP_sw1_7_), .B(DP_mult_205_n2304), .ZN(
        DP_mult_205_n1648) );
  XNOR2_X1 DP_mult_205_U2218 ( .A(DP_sw1_7_), .B(DP_mult_205_n2287), .ZN(
        DP_mult_205_n1748) );
  XNOR2_X1 DP_mult_205_U2217 ( .A(DP_sw1_7_), .B(DP_mult_205_n2299), .ZN(
        DP_mult_205_n1673) );
  XNOR2_X1 DP_mult_205_U2216 ( .A(DP_sw1_7_), .B(DP_mult_205_n2327), .ZN(
        DP_mult_205_n1498) );
  XNOR2_X1 DP_mult_205_U2215 ( .A(DP_sw1_7_), .B(DP_mult_205_n2318), .ZN(
        DP_mult_205_n1548) );
  XNOR2_X1 DP_mult_205_U2214 ( .A(DP_sw1_7_), .B(DP_mult_205_n2324), .ZN(
        DP_mult_205_n1523) );
  XNOR2_X1 DP_mult_205_U2213 ( .A(DP_sw1_7_), .B(DP_mult_205_n2307), .ZN(
        DP_mult_205_n1623) );
  XNOR2_X1 DP_mult_205_U2212 ( .A(DP_sw1_7_), .B(DP_mult_205_n2016), .ZN(
        DP_mult_205_n1698) );
  XNOR2_X1 DP_mult_205_U2211 ( .A(DP_sw1_7_), .B(DP_mult_205_n2314), .ZN(
        DP_mult_205_n1573) );
  XNOR2_X1 DP_mult_205_U2210 ( .A(DP_sw1_7_), .B(DP_mult_205_n2310), .ZN(
        DP_mult_205_n1598) );
  XNOR2_X1 DP_mult_205_U2209 ( .A(DP_sw1_9_), .B(DP_mult_205_n2326), .ZN(
        DP_mult_205_n1496) );
  XNOR2_X1 DP_mult_205_U2208 ( .A(DP_sw1_9_), .B(DP_mult_205_n2299), .ZN(
        DP_mult_205_n1671) );
  XNOR2_X1 DP_mult_205_U2207 ( .A(DP_sw1_9_), .B(DP_mult_205_n2323), .ZN(
        DP_mult_205_n1521) );
  XNOR2_X1 DP_mult_205_U2206 ( .A(DP_sw1_5_), .B(DP_mult_205_n2307), .ZN(
        DP_mult_205_n1625) );
  XNOR2_X1 DP_mult_205_U2205 ( .A(DP_sw1_9_), .B(DP_mult_205_n2290), .ZN(
        DP_mult_205_n1721) );
  XNOR2_X1 DP_mult_205_U2204 ( .A(DP_sw1_1_), .B(DP_mult_205_n2313), .ZN(
        DP_mult_205_n1579) );
  XNOR2_X1 DP_mult_205_U2203 ( .A(DP_sw1_5_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1600) );
  XNOR2_X1 DP_mult_205_U2202 ( .A(DP_sw1_5_), .B(DP_mult_205_n2291), .ZN(
        DP_mult_205_n1725) );
  XNOR2_X1 DP_mult_205_U2201 ( .A(DP_sw1_3_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1602) );
  XNOR2_X1 DP_mult_205_U2200 ( .A(DP_sw1_3_), .B(DP_mult_205_n2292), .ZN(
        DP_mult_205_n1727) );
  XNOR2_X1 DP_mult_205_U2199 ( .A(DP_sw1_5_), .B(DP_mult_205_n2327), .ZN(
        DP_mult_205_n1500) );
  XNOR2_X1 DP_mult_205_U2198 ( .A(DP_sw1_1_), .B(DP_mult_205_n2015), .ZN(
        DP_mult_205_n1704) );
  XNOR2_X1 DP_mult_205_U2197 ( .A(DP_sw1_1_), .B(DP_mult_205_n2306), .ZN(
        DP_mult_205_n1629) );
  XNOR2_X1 DP_mult_205_U2196 ( .A(DP_sw1_3_), .B(DP_mult_205_n2313), .ZN(
        DP_mult_205_n1577) );
  XNOR2_X1 DP_mult_205_U2195 ( .A(DP_sw1_3_), .B(DP_mult_205_n2327), .ZN(
        DP_mult_205_n1502) );
  XNOR2_X1 DP_mult_205_U2194 ( .A(DP_sw1_9_), .B(DP_mult_205_n2319), .ZN(
        DP_mult_205_n1546) );
  XNOR2_X1 DP_mult_205_U2193 ( .A(DP_sw1_5_), .B(DP_mult_205_n2324), .ZN(
        DP_mult_205_n1525) );
  XNOR2_X1 DP_mult_205_U2192 ( .A(DP_sw1_1_), .B(DP_mult_205_n2327), .ZN(
        DP_mult_205_n1504) );
  XNOR2_X1 DP_mult_205_U2191 ( .A(DP_sw1_3_), .B(DP_mult_205_n2302), .ZN(
        DP_mult_205_n1652) );
  XNOR2_X1 DP_mult_205_U2190 ( .A(DP_sw1_5_), .B(DP_mult_205_n2303), .ZN(
        DP_mult_205_n1650) );
  XNOR2_X1 DP_mult_205_U2189 ( .A(DP_sw1_5_), .B(DP_mult_205_n2015), .ZN(
        DP_mult_205_n1700) );
  XNOR2_X1 DP_mult_205_U2188 ( .A(DP_sw1_9_), .B(DP_mult_205_n2313), .ZN(
        DP_mult_205_n1571) );
  XNOR2_X1 DP_mult_205_U2187 ( .A(DP_sw1_9_), .B(DP_mult_205_n2288), .ZN(
        DP_mult_205_n1746) );
  XNOR2_X1 DP_mult_205_U2186 ( .A(DP_sw1_9_), .B(DP_mult_205_n2015), .ZN(
        DP_mult_205_n1696) );
  XNOR2_X1 DP_mult_205_U2185 ( .A(DP_sw1_3_), .B(DP_mult_205_n2288), .ZN(
        DP_mult_205_n1752) );
  XNOR2_X1 DP_mult_205_U2184 ( .A(DP_sw1_3_), .B(DP_mult_205_n2298), .ZN(
        DP_mult_205_n1677) );
  XNOR2_X1 DP_mult_205_U2183 ( .A(DP_sw1_9_), .B(DP_mult_205_n2311), .ZN(
        DP_mult_205_n1596) );
  XNOR2_X1 DP_mult_205_U2182 ( .A(DP_sw1_9_), .B(DP_mult_205_n2307), .ZN(
        DP_mult_205_n1621) );
  XNOR2_X1 DP_mult_205_U2181 ( .A(DP_sw1_1_), .B(DP_mult_205_n2290), .ZN(
        DP_mult_205_n1729) );
  XNOR2_X1 DP_mult_205_U2180 ( .A(DP_sw1_5_), .B(DP_mult_205_n2320), .ZN(
        DP_mult_205_n1550) );
  XNOR2_X1 DP_mult_205_U2179 ( .A(DP_sw1_5_), .B(DP_mult_205_n2300), .ZN(
        DP_mult_205_n1675) );
  XNOR2_X1 DP_mult_205_U2178 ( .A(DP_sw1_9_), .B(DP_mult_205_n2303), .ZN(
        DP_mult_205_n1646) );
  XNOR2_X1 DP_mult_205_U2177 ( .A(DP_sw1_1_), .B(DP_mult_205_n2324), .ZN(
        DP_mult_205_n1529) );
  XNOR2_X1 DP_mult_205_U2176 ( .A(DP_sw1_1_), .B(DP_mult_205_n2319), .ZN(
        DP_mult_205_n1554) );
  XNOR2_X1 DP_mult_205_U2175 ( .A(DP_sw1_3_), .B(DP_mult_205_n2319), .ZN(
        DP_mult_205_n1552) );
  XNOR2_X1 DP_mult_205_U2174 ( .A(DP_sw1_1_), .B(DP_mult_205_n2303), .ZN(
        DP_mult_205_n1654) );
  XNOR2_X1 DP_mult_205_U2173 ( .A(DP_sw1_1_), .B(DP_mult_205_n2300), .ZN(
        DP_mult_205_n1679) );
  XNOR2_X1 DP_mult_205_U2172 ( .A(DP_sw1_5_), .B(DP_mult_205_n2313), .ZN(
        DP_mult_205_n1575) );
  XNOR2_X1 DP_mult_205_U2171 ( .A(DP_sw1_3_), .B(DP_mult_205_n2324), .ZN(
        DP_mult_205_n1527) );
  XNOR2_X1 DP_mult_205_U2170 ( .A(DP_sw1_5_), .B(DP_mult_205_n2287), .ZN(
        DP_mult_205_n1750) );
  XNOR2_X1 DP_mult_205_U2169 ( .A(DP_sw1_1_), .B(DP_mult_205_n2310), .ZN(
        DP_mult_205_n1604) );
  XNOR2_X1 DP_mult_205_U2168 ( .A(DP_sw1_3_), .B(DP_mult_205_n2308), .ZN(
        DP_mult_205_n1627) );
  XNOR2_X1 DP_mult_205_U2167 ( .A(DP_sw1_3_), .B(DP_mult_205_n2016), .ZN(
        DP_mult_205_n1702) );
  XNOR2_X1 DP_mult_205_U2166 ( .A(DP_sw1_1_), .B(DP_mult_205_n2287), .ZN(
        DP_mult_205_n1754) );
  XNOR2_X1 DP_mult_205_U2165 ( .A(DP_mult_205_n2296), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1705) );
  XNOR2_X1 DP_mult_205_U2164 ( .A(DP_mult_205_n2291), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1730) );
  OAI22_X1 DP_mult_205_U2163 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1776), 
        .B1(DP_mult_205_n1775), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1477)
         );
  XNOR2_X1 DP_mult_205_U2162 ( .A(DP_sw1_23_), .B(DP_mult_205_n2323), .ZN(
        DP_mult_205_n1507) );
  XNOR2_X1 DP_mult_205_U2161 ( .A(DP_sw1_23_), .B(DP_mult_205_n2320), .ZN(
        DP_mult_205_n1532) );
  XNOR2_X1 DP_mult_205_U2160 ( .A(DP_sw1_23_), .B(DP_mult_205_n2310), .ZN(
        DP_mult_205_n1582) );
  XNOR2_X1 DP_mult_205_U2159 ( .A(DP_sw1_23_), .B(DP_mult_205_n2313), .ZN(
        DP_mult_205_n1557) );
  XNOR2_X1 DP_mult_205_U2158 ( .A(DP_sw1_23_), .B(DP_mult_205_n2299), .ZN(
        DP_mult_205_n1657) );
  XNOR2_X1 DP_mult_205_U2157 ( .A(DP_sw1_23_), .B(DP_mult_205_n2304), .ZN(
        DP_mult_205_n1632) );
  XNOR2_X1 DP_mult_205_U2156 ( .A(DP_sw1_23_), .B(DP_mult_205_n2307), .ZN(
        DP_mult_205_n1607) );
  XNOR2_X1 DP_mult_205_U2155 ( .A(DP_sw1_23_), .B(DP_mult_205_n2292), .ZN(
        DP_mult_205_n1707) );
  XNOR2_X1 DP_mult_205_U2154 ( .A(DP_sw1_23_), .B(DP_mult_205_n2288), .ZN(
        DP_mult_205_n1732) );
  XNOR2_X1 DP_mult_205_U2153 ( .A(DP_sw1_23_), .B(DP_mult_205_n2016), .ZN(
        DP_mult_205_n1682) );
  XNOR2_X1 DP_mult_205_U2152 ( .A(DP_sw1_7_), .B(DP_mult_205_n2284), .ZN(
        DP_mult_205_n1773) );
  XNOR2_X1 DP_mult_205_U2151 ( .A(DP_mult_205_n2299), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1674) );
  XNOR2_X1 DP_mult_205_U2150 ( .A(DP_mult_205_n2288), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1749) );
  XNOR2_X1 DP_mult_205_U2149 ( .A(DP_mult_205_n2323), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1524) );
  XNOR2_X1 DP_mult_205_U2148 ( .A(DP_mult_205_n2302), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1649) );
  XNOR2_X1 DP_mult_205_U2147 ( .A(DP_mult_205_n2326), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1499) );
  XNOR2_X1 DP_mult_205_U2146 ( .A(DP_mult_205_n2319), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1549) );
  XNOR2_X1 DP_mult_205_U2145 ( .A(DP_mult_205_n2308), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1624) );
  XNOR2_X1 DP_mult_205_U2144 ( .A(DP_mult_205_n2295), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1699) );
  XNOR2_X1 DP_mult_205_U2143 ( .A(DP_mult_205_n2315), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1574) );
  XNOR2_X1 DP_mult_205_U2142 ( .A(DP_mult_205_n2311), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1599) );
  XNOR2_X1 DP_mult_205_U2141 ( .A(DP_sw1_23_), .B(DP_mult_205_n2282), .ZN(
        DP_mult_205_n1757) );
  XNOR2_X1 DP_mult_205_U2140 ( .A(DP_mult_205_n2326), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1483) );
  XNOR2_X1 DP_mult_205_U2139 ( .A(DP_mult_205_n2326), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1487) );
  XNOR2_X1 DP_mult_205_U2138 ( .A(DP_mult_205_n2322), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1508) );
  XNOR2_X1 DP_mult_205_U2137 ( .A(DP_mult_205_n2318), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1533) );
  XNOR2_X1 DP_mult_205_U2136 ( .A(DP_mult_205_n2323), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1514) );
  XNOR2_X1 DP_mult_205_U2135 ( .A(DP_mult_205_n2292), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1720) );
  XNOR2_X1 DP_mult_205_U2134 ( .A(DP_mult_205_n2322), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1518) );
  XNOR2_X1 DP_mult_205_U2133 ( .A(DP_mult_205_n2326), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1489) );
  XNOR2_X1 DP_mult_205_U2132 ( .A(DP_mult_205_n2310), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1583) );
  XNOR2_X1 DP_mult_205_U2131 ( .A(DP_mult_205_n2316), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1566) );
  XNOR2_X1 DP_mult_205_U2130 ( .A(DP_mult_205_n2323), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1512) );
  XNOR2_X1 DP_mult_205_U2129 ( .A(DP_mult_205_n2318), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1537) );
  XNOR2_X1 DP_mult_205_U2128 ( .A(DP_mult_205_n2322), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1520) );
  XNOR2_X1 DP_mult_205_U2127 ( .A(DP_mult_205_n2315), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1562) );
  XNOR2_X1 DP_mult_205_U2126 ( .A(DP_mult_205_n2310), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1589) );
  XNOR2_X1 DP_mult_205_U2125 ( .A(DP_mult_205_n2318), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1541) );
  XNOR2_X1 DP_mult_205_U2124 ( .A(DP_mult_205_n2326), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1495) );
  XNOR2_X1 DP_mult_205_U2123 ( .A(DP_mult_205_n2306), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1612) );
  XNOR2_X1 DP_mult_205_U2122 ( .A(DP_mult_205_n2290), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1716) );
  XNOR2_X1 DP_mult_205_U2121 ( .A(DP_mult_205_n2318), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1543) );
  XNOR2_X1 DP_mult_205_U2120 ( .A(DP_mult_205_n2326), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1491) );
  XNOR2_X1 DP_mult_205_U2119 ( .A(DP_mult_205_n2326), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1493) );
  XNOR2_X1 DP_mult_205_U2118 ( .A(DP_mult_205_n2315), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1564) );
  XNOR2_X1 DP_mult_205_U2117 ( .A(DP_mult_205_n2296), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1689) );
  XNOR2_X1 DP_mult_205_U2116 ( .A(DP_mult_205_n2316), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1558) );
  XNOR2_X1 DP_mult_205_U2115 ( .A(DP_mult_205_n2311), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1587) );
  XNOR2_X1 DP_mult_205_U2114 ( .A(DP_mult_205_n2323), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1516) );
  XNOR2_X1 DP_mult_205_U2113 ( .A(DP_mult_205_n2318), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1539) );
  XNOR2_X1 DP_mult_205_U2112 ( .A(DP_mult_205_n2288), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1739) );
  XNOR2_X1 DP_mult_205_U2111 ( .A(DP_mult_205_n2299), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1670) );
  XNOR2_X1 DP_mult_205_U2110 ( .A(DP_mult_205_n2295), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1687) );
  XNOR2_X1 DP_mult_205_U2109 ( .A(DP_mult_205_n2303), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1639) );
  XNOR2_X1 DP_mult_205_U2108 ( .A(DP_mult_205_n2316), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1570) );
  XNOR2_X1 DP_mult_205_U2107 ( .A(DP_mult_205_n2310), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1593) );
  XNOR2_X1 DP_mult_205_U2106 ( .A(DP_mult_205_n2292), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1718) );
  XNOR2_X1 DP_mult_205_U2105 ( .A(DP_mult_205_n2295), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1695) );
  XNOR2_X1 DP_mult_205_U2104 ( .A(DP_mult_205_n2303), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1633) );
  XNOR2_X1 DP_mult_205_U2103 ( .A(DP_mult_205_n2295), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1691) );
  XNOR2_X1 DP_mult_205_U2102 ( .A(DP_mult_205_n2307), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1614) );
  XNOR2_X1 DP_mult_205_U2101 ( .A(DP_mult_205_n2318), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1545) );
  XNOR2_X1 DP_mult_205_U2100 ( .A(DP_mult_205_n2300), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1664) );
  XNOR2_X1 DP_mult_205_U2099 ( .A(DP_mult_205_n2306), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1608) );
  XNOR2_X1 DP_mult_205_U2098 ( .A(DP_mult_205_n2306), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1620) );
  XNOR2_X1 DP_mult_205_U2097 ( .A(DP_mult_205_n2308), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1616) );
  XNOR2_X1 DP_mult_205_U2096 ( .A(DP_mult_205_n2300), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1662) );
  XNOR2_X1 DP_mult_205_U2095 ( .A(DP_mult_205_n2287), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1741) );
  XNOR2_X1 DP_mult_205_U2094 ( .A(DP_mult_205_n2288), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1743) );
  XNOR2_X1 DP_mult_205_U2093 ( .A(DP_mult_205_n2287), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1745) );
  XNOR2_X1 DP_mult_205_U2092 ( .A(DP_mult_205_n2290), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1708) );
  XNOR2_X1 DP_mult_205_U2091 ( .A(DP_mult_205_n2298), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1666) );
  XNOR2_X1 DP_mult_205_U2090 ( .A(DP_mult_205_n2310), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1591) );
  XNOR2_X1 DP_mult_205_U2089 ( .A(DP_mult_205_n2306), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1618) );
  XNOR2_X1 DP_mult_205_U2088 ( .A(DP_mult_205_n2300), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1658) );
  XNOR2_X1 DP_mult_205_U2087 ( .A(DP_mult_205_n2310), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1595) );
  XNOR2_X1 DP_mult_205_U2086 ( .A(DP_mult_205_n2288), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1737) );
  XNOR2_X1 DP_mult_205_U2085 ( .A(DP_mult_205_n2304), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1645) );
  XNOR2_X1 DP_mult_205_U2084 ( .A(DP_mult_205_n2304), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1641) );
  XNOR2_X1 DP_mult_205_U2083 ( .A(DP_mult_205_n2316), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1568) );
  XNOR2_X1 DP_mult_205_U2082 ( .A(DP_mult_205_n2304), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1637) );
  XNOR2_X1 DP_mult_205_U2081 ( .A(DP_mult_205_n2287), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1733) );
  XNOR2_X1 DP_mult_205_U2080 ( .A(DP_mult_205_n2290), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1712) );
  XNOR2_X1 DP_mult_205_U2079 ( .A(DP_mult_205_n2303), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1643) );
  XNOR2_X1 DP_mult_205_U2078 ( .A(DP_mult_205_n2296), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1683) );
  XNOR2_X1 DP_mult_205_U2077 ( .A(DP_mult_205_n2291), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1714) );
  XNOR2_X1 DP_mult_205_U2076 ( .A(DP_mult_205_n2295), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1693) );
  XNOR2_X1 DP_mult_205_U2075 ( .A(DP_mult_205_n2300), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1668) );
  XNOR2_X1 DP_mult_205_U2074 ( .A(DP_sw1_9_), .B(DP_mult_205_n2285), .ZN(
        DP_mult_205_n1771) );
  XNOR2_X1 DP_mult_205_U2073 ( .A(DP_sw1_1_), .B(DP_mult_205_n2282), .ZN(
        DP_mult_205_n1779) );
  XNOR2_X1 DP_mult_205_U2072 ( .A(DP_sw1_5_), .B(DP_mult_205_n2285), .ZN(
        DP_mult_205_n1775) );
  XNOR2_X1 DP_mult_205_U2071 ( .A(DP_sw1_3_), .B(DP_mult_205_n2284), .ZN(
        DP_mult_205_n1777) );
  XNOR2_X1 DP_mult_205_U2070 ( .A(DP_mult_205_n2320), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1535) );
  XNOR2_X1 DP_mult_205_U2069 ( .A(DP_mult_205_n2322), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1510) );
  XNOR2_X1 DP_mult_205_U2068 ( .A(DP_mult_205_n2326), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1485) );
  XNOR2_X1 DP_mult_205_U2067 ( .A(DP_mult_205_n2314), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1560) );
  XNOR2_X1 DP_mult_205_U2066 ( .A(DP_mult_205_n2299), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1660) );
  XNOR2_X1 DP_mult_205_U2065 ( .A(DP_mult_205_n2304), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1635) );
  XNOR2_X1 DP_mult_205_U2064 ( .A(DP_mult_205_n2307), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1610) );
  XNOR2_X1 DP_mult_205_U2063 ( .A(DP_mult_205_n2290), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1726) );
  XNOR2_X1 DP_mult_205_U2062 ( .A(DP_mult_205_n2310), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1585) );
  XNOR2_X1 DP_mult_205_U2061 ( .A(DP_mult_205_n2310), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1601) );
  XNOR2_X1 DP_mult_205_U2060 ( .A(DP_mult_205_n2295), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1701) );
  XNOR2_X1 DP_mult_205_U2059 ( .A(DP_mult_205_n2302), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1647) );
  XNOR2_X1 DP_mult_205_U2058 ( .A(DP_mult_205_n2288), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1747) );
  XNOR2_X1 DP_mult_205_U2057 ( .A(DP_mult_205_n2299), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1672) );
  XNOR2_X1 DP_mult_205_U2056 ( .A(DP_mult_205_n2319), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1547) );
  XNOR2_X1 DP_mult_205_U2055 ( .A(DP_mult_205_n2308), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1626) );
  XNOR2_X1 DP_mult_205_U2054 ( .A(DP_mult_205_n2287), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1753) );
  XNOR2_X1 DP_mult_205_U2053 ( .A(DP_mult_205_n2296), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1685) );
  XNOR2_X1 DP_mult_205_U2052 ( .A(DP_mult_205_n2292), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1722) );
  XNOR2_X1 DP_mult_205_U2051 ( .A(DP_mult_205_n2324), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1522) );
  XNOR2_X1 DP_mult_205_U2050 ( .A(DP_mult_205_n2314), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1578) );
  XNOR2_X1 DP_mult_205_U2049 ( .A(DP_mult_205_n2326), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1501) );
  XNOR2_X1 DP_mult_205_U2048 ( .A(DP_mult_205_n2291), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1728) );
  XNOR2_X1 DP_mult_205_U2047 ( .A(DP_mult_205_n2310), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1603) );
  XNOR2_X1 DP_mult_205_U2046 ( .A(DP_mult_205_n2303), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1651) );
  XNOR2_X1 DP_mult_205_U2045 ( .A(DP_mult_205_n2292), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1710) );
  XNOR2_X1 DP_mult_205_U2044 ( .A(DP_mult_205_n2295), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1697) );
  XNOR2_X1 DP_mult_205_U2043 ( .A(DP_mult_205_n2299), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1678) );
  XNOR2_X1 DP_mult_205_U2042 ( .A(DP_mult_205_n2319), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1551) );
  XNOR2_X1 DP_mult_205_U2041 ( .A(DP_mult_205_n2310), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1597) );
  XNOR2_X1 DP_mult_205_U2040 ( .A(DP_mult_205_n2324), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1526) );
  XNOR2_X1 DP_mult_205_U2039 ( .A(DP_mult_205_n2287), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1735) );
  XNOR2_X1 DP_mult_205_U2038 ( .A(DP_mult_205_n2326), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1497) );
  XNOR2_X1 DP_mult_205_U2037 ( .A(DP_mult_205_n2315), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1572) );
  XNOR2_X1 DP_mult_205_U2036 ( .A(DP_mult_205_n2327), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1503) );
  XNOR2_X1 DP_mult_205_U2035 ( .A(DP_mult_205_n2298), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1676) );
  XNOR2_X1 DP_mult_205_U2034 ( .A(DP_mult_205_n2306), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1622) );
  XNOR2_X1 DP_mult_205_U2033 ( .A(DP_mult_205_n2320), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1553) );
  XNOR2_X1 DP_mult_205_U2032 ( .A(DP_mult_205_n2287), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1751) );
  XNOR2_X1 DP_mult_205_U2031 ( .A(DP_mult_205_n2302), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1653) );
  XNOR2_X1 DP_mult_205_U2030 ( .A(DP_mult_205_n2295), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1703) );
  XNOR2_X1 DP_mult_205_U2029 ( .A(DP_mult_205_n2324), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1528) );
  XNOR2_X1 DP_mult_205_U2028 ( .A(DP_mult_205_n2314), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1576) );
  XNOR2_X1 DP_mult_205_U2027 ( .A(DP_mult_205_n2308), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1628) );
  XNOR2_X1 DP_mult_205_U2026 ( .A(DP_mult_205_n2282), .B(DP_sw1_10_), .ZN(
        DP_mult_205_n1770) );
  XNOR2_X1 DP_mult_205_U2025 ( .A(DP_mult_205_n2326), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1505) );
  XNOR2_X1 DP_mult_205_U2024 ( .A(DP_mult_205_n2323), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1530) );
  XNOR2_X1 DP_mult_205_U2023 ( .A(DP_mult_205_n2299), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1680) );
  XNOR2_X1 DP_mult_205_U2022 ( .A(DP_mult_205_n2282), .B(DP_sw1_6_), .ZN(
        DP_mult_205_n1774) );
  XNOR2_X1 DP_mult_205_U2021 ( .A(DP_mult_205_n2285), .B(DP_sw1_16_), .ZN(
        DP_mult_205_n1764) );
  XNOR2_X1 DP_mult_205_U2020 ( .A(DP_mult_205_n2282), .B(DP_sw1_14_), .ZN(
        DP_mult_205_n1766) );
  XNOR2_X1 DP_mult_205_U2019 ( .A(DP_mult_205_n2284), .B(DP_sw1_22_), .ZN(
        DP_mult_205_n1758) );
  XNOR2_X1 DP_mult_205_U2018 ( .A(DP_mult_205_n2284), .B(DP_sw1_12_), .ZN(
        DP_mult_205_n1768) );
  XNOR2_X1 DP_mult_205_U2017 ( .A(DP_mult_205_n2284), .B(DP_sw1_18_), .ZN(
        DP_mult_205_n1762) );
  XNOR2_X1 DP_mult_205_U2016 ( .A(DP_mult_205_n2285), .B(DP_sw1_20_), .ZN(
        DP_mult_205_n1760) );
  XNOR2_X1 DP_mult_205_U2015 ( .A(DP_mult_205_n2282), .B(DP_sw1_8_), .ZN(
        DP_mult_205_n1772) );
  XNOR2_X1 DP_mult_205_U2014 ( .A(DP_mult_205_n2284), .B(DP_sw1_4_), .ZN(
        DP_mult_205_n1776) );
  XNOR2_X1 DP_mult_205_U2013 ( .A(DP_mult_205_n2285), .B(DP_sw1_2_), .ZN(
        DP_mult_205_n1778) );
  XNOR2_X1 DP_mult_205_U2012 ( .A(DP_mult_205_n2304), .B(DP_sw1_0_), .ZN(
        DP_mult_205_n1655) );
  INV_X1 DP_mult_205_U2011 ( .A(DP_mult_205_n1482), .ZN(DP_mult_205_n2341) );
  INV_X1 DP_mult_205_U2010 ( .A(DP_mult_205_n1582), .ZN(DP_mult_205_n2337) );
  INV_X1 DP_mult_205_U2009 ( .A(DP_mult_205_n1732), .ZN(DP_mult_205_n2331) );
  INV_X1 DP_mult_205_U2008 ( .A(DP_mult_205_n724), .ZN(DP_mult_205_n725) );
  INV_X1 DP_mult_205_U2007 ( .A(DP_mult_205_n1657), .ZN(DP_mult_205_n2334) );
  INV_X1 DP_mult_205_U2006 ( .A(DP_mult_205_n692), .ZN(DP_mult_205_n693) );
  OAI22_X1 DP_mult_205_U2005 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1767), 
        .B1(DP_mult_205_n1766), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1468)
         );
  OAI22_X1 DP_mult_205_U2004 ( .A1(DP_mult_205_n1949), .A2(DP_mult_205_n1762), 
        .B1(DP_mult_205_n1761), .B2(DP_mult_205_n2281), .ZN(DP_mult_205_n1463)
         );
  OAI22_X1 DP_mult_205_U2003 ( .A1(DP_mult_205_n1949), .A2(DP_mult_205_n1759), 
        .B1(DP_mult_205_n1758), .B2(DP_mult_205_n2281), .ZN(DP_mult_205_n1460)
         );
  INV_X1 DP_mult_205_U2002 ( .A(DP_mult_205_n1607), .ZN(DP_mult_205_n2336) );
  OAI21_X1 DP_mult_205_U2001 ( .B1(DP_mult_205_n2243), .B2(DP_mult_205_n1996), 
        .A(DP_mult_205_n2336), .ZN(DP_mult_205_n1314) );
  NOR2_X1 DP_mult_205_U2000 ( .A1(DP_mult_205_n2263), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1289) );
  NOR2_X1 DP_mult_205_U1999 ( .A1(DP_mult_205_n2267), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1337) );
  OAI22_X1 DP_mult_205_U1998 ( .A1(DP_mult_205_n1949), .A2(DP_mult_205_n1765), 
        .B1(DP_mult_205_n1764), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1466)
         );
  OAI22_X1 DP_mult_205_U1997 ( .A1(DP_mult_205_n1949), .A2(DP_mult_205_n1766), 
        .B1(DP_mult_205_n1765), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1467)
         );
  OAI22_X1 DP_mult_205_U1996 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1768), 
        .B1(DP_mult_205_n1767), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1469)
         );
  INV_X1 DP_mult_205_U1995 ( .A(DP_mult_205_n802), .ZN(DP_mult_205_n803) );
  INV_X1 DP_mult_205_U1994 ( .A(DP_mult_205_n1707), .ZN(DP_mult_205_n2332) );
  NOR2_X1 DP_mult_205_U1993 ( .A1(DP_mult_205_n2256), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1241) );
  OAI22_X1 DP_mult_205_U1992 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1771), 
        .B1(DP_mult_205_n1770), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1472)
         );
  NOR2_X1 DP_mult_205_U1991 ( .A1(DP_mult_205_n2259), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1265) );
  OAI22_X1 DP_mult_205_U1990 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1775), 
        .B1(DP_mult_205_n1774), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1476)
         );
  OAI22_X1 DP_mult_205_U1989 ( .A1(DP_mult_205_n1994), .A2(DP_mult_205_n1772), 
        .B1(DP_mult_205_n1771), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1473)
         );
  INV_X1 DP_mult_205_U1988 ( .A(DP_mult_205_n1682), .ZN(DP_mult_205_n2333) );
  INV_X1 DP_mult_205_U1987 ( .A(DP_mult_205_n1557), .ZN(DP_mult_205_n2338) );
  OAI21_X1 DP_mult_205_U1986 ( .B1(DP_mult_205_n1934), .B2(DP_mult_205_n2275), 
        .A(DP_mult_205_n2334), .ZN(DP_mult_205_n1362) );
  OAI22_X1 DP_mult_205_U1985 ( .A1(DP_mult_205_n1949), .A2(DP_mult_205_n1763), 
        .B1(DP_mult_205_n1762), .B2(DP_mult_205_n2281), .ZN(DP_mult_205_n1464)
         );
  OAI22_X1 DP_mult_205_U1984 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1769), 
        .B1(DP_mult_205_n1768), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1470)
         );
  NOR2_X1 DP_mult_205_U1983 ( .A1(DP_mult_205_n2265), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1313) );
  NOR2_X1 DP_mult_205_U1982 ( .A1(DP_mult_205_n2271), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1361) );
  NOR2_X1 DP_mult_205_U1981 ( .A1(DP_mult_205_n2254), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1217) );
  OAI22_X1 DP_mult_205_U1980 ( .A1(DP_mult_205_n1949), .A2(DP_mult_205_n1761), 
        .B1(DP_mult_205_n1760), .B2(DP_mult_205_n2281), .ZN(DP_mult_205_n1462)
         );
  NOR2_X1 DP_mult_205_U1979 ( .A1(DP_mult_205_n1982), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1409) );
  INV_X1 DP_mult_205_U1978 ( .A(DP_mult_205_n1532), .ZN(DP_mult_205_n2339) );
  OAI21_X1 DP_mult_205_U1977 ( .B1(DP_mult_205_n1985), .B2(DP_mult_205_n1986), 
        .A(DP_mult_205_n2339), .ZN(DP_mult_205_n1242) );
  NOR2_X1 DP_mult_205_U1976 ( .A1(DP_mult_205_n2273), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1385) );
  OAI22_X1 DP_mult_205_U1975 ( .A1(DP_mult_205_n1994), .A2(DP_mult_205_n1777), 
        .B1(DP_mult_205_n1776), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1478)
         );
  OAI22_X1 DP_mult_205_U1974 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1764), 
        .B1(DP_mult_205_n1763), .B2(DP_mult_205_n2281), .ZN(DP_mult_205_n1465)
         );
  INV_X1 DP_mult_205_U1973 ( .A(DP_mult_205_n1632), .ZN(DP_mult_205_n2335) );
  NAND2_X1 DP_mult_205_U1972 ( .A1(DP_mult_205_n2299), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1681) );
  NAND2_X1 DP_mult_205_U1971 ( .A1(DP_mult_205_n2323), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1531) );
  NAND2_X1 DP_mult_205_U1970 ( .A1(DP_mult_205_n2310), .A2(DP_mult_205_n2329), 
        .ZN(DP_mult_205_n1606) );
  NAND2_X1 DP_mult_205_U1969 ( .A1(DP_mult_205_n2304), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1656) );
  NAND2_X1 DP_mult_205_U1968 ( .A1(DP_mult_205_n2295), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1706) );
  NAND2_X1 DP_mult_205_U1967 ( .A1(DP_mult_205_n2307), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1631) );
  NAND2_X1 DP_mult_205_U1966 ( .A1(DP_mult_205_n2326), .A2(DP_mult_205_n2329), 
        .ZN(DP_mult_205_n1506) );
  NAND2_X1 DP_mult_205_U1965 ( .A1(DP_mult_205_n2315), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1581) );
  NAND2_X1 DP_mult_205_U1964 ( .A1(DP_mult_205_n2320), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1556) );
  CLKBUF_X1 DP_mult_205_U1963 ( .A(DP_mult_205_n251), .Z(DP_mult_205_n2281) );
  NAND2_X1 DP_mult_205_U1962 ( .A1(DP_mult_205_n2282), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1781) );
  AOI21_X1 DP_mult_205_U1961 ( .B1(DP_mult_205_n1943), .B2(DP_mult_205_n1942), 
        .A(DP_mult_205_n1951), .ZN(DP_mult_205_n646) );
  NOR2_X1 DP_mult_205_U1960 ( .A1(DP_mult_205_n2042), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1433) );
  INV_X1 DP_mult_205_U1959 ( .A(DP_mult_205_n2199), .ZN(DP_mult_205_n2261) );
  INV_X1 DP_mult_205_U1958 ( .A(DP_mult_205_n2205), .ZN(DP_mult_205_n2264) );
  INV_X1 DP_mult_205_U1957 ( .A(DP_mult_205_n2317), .ZN(DP_mult_205_n2313) );
  INV_X1 DP_mult_205_U1956 ( .A(DP_mult_205_n2044), .ZN(DP_mult_205_n2298) );
  INV_X1 DP_mult_205_U1955 ( .A(DP_mult_205_n2305), .ZN(DP_mult_205_n2302) );
  INV_X1 DP_mult_205_U1954 ( .A(DP_mult_205_n2164), .ZN(DP_mult_205_n2294) );
  INV_X1 DP_mult_205_U1953 ( .A(DP_mult_205_n2204), .ZN(DP_mult_205_n2256) );
  INV_X1 DP_mult_205_U1952 ( .A(DP_mult_205_n2275), .ZN(DP_mult_205_n2273) );
  INV_X1 DP_mult_205_U1951 ( .A(DP_mult_205_n1992), .ZN(DP_mult_205_n2262) );
  INV_X1 DP_mult_205_U1950 ( .A(DP_mult_205_n2205), .ZN(DP_mult_205_n2265) );
  INV_X1 DP_mult_205_U1949 ( .A(DP_mult_205_n1940), .ZN(DP_mult_205_n2233) );
  INV_X1 DP_mult_205_U1948 ( .A(DP_mult_205_n2049), .ZN(DP_mult_205_n2234) );
  INV_X1 DP_mult_205_U1947 ( .A(DP_mult_205_n2101), .ZN(DP_mult_205_n2240) );
  NAND2_X1 DP_mult_205_U1946 ( .A1(DP_mult_205_n2292), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1731) );
  INV_X1 DP_mult_205_U1945 ( .A(DP_mult_205_n682), .ZN(DP_mult_205_n683) );
  INV_X1 DP_mult_205_U1944 ( .A(DP_mult_205_n1507), .ZN(DP_mult_205_n2340) );
  OAI21_X1 DP_mult_205_U1943 ( .B1(DP_mult_205_n1971), .B2(DP_mult_205_n2204), 
        .A(DP_mult_205_n2340), .ZN(DP_mult_205_n1218) );
  OAI22_X1 DP_mult_205_U1942 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1774), 
        .B1(DP_mult_205_n1773), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1475)
         );
  OAI22_X1 DP_mult_205_U1941 ( .A1(DP_mult_205_n2253), .A2(DP_mult_205_n1773), 
        .B1(DP_mult_205_n1772), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1474)
         );
  OAI22_X1 DP_mult_205_U1940 ( .A1(DP_mult_205_n1949), .A2(DP_mult_205_n1760), 
        .B1(DP_mult_205_n1759), .B2(DP_mult_205_n2281), .ZN(DP_mult_205_n1461)
         );
  NAND2_X1 DP_mult_205_U1939 ( .A1(DP_mult_205_n2288), .A2(DP_mult_205_n1930), 
        .ZN(DP_mult_205_n1756) );
  NOR2_X1 DP_mult_205_U1938 ( .A1(DP_mult_205_n1973), .A2(DP_mult_205_n1931), 
        .ZN(DP_mult_205_n1457) );
  INV_X1 DP_mult_205_U1937 ( .A(DP_mult_205_n2309), .ZN(DP_mult_205_n2307) );
  INV_X1 DP_mult_205_U1936 ( .A(DP_mult_205_n2164), .ZN(DP_mult_205_n2295) );
  OAI22_X1 DP_mult_205_U1935 ( .A1(DP_mult_205_n1994), .A2(DP_mult_205_n1779), 
        .B1(DP_mult_205_n1778), .B2(DP_mult_205_n2280), .ZN(DP_mult_205_n1480)
         );
  INV_X1 DP_mult_205_U1934 ( .A(DP_mult_205_n2289), .ZN(DP_mult_205_n2287) );
  AND2_X1 DP_mult_205_U1933 ( .A1(DP_mult_205_n1194), .A2(DP_mult_205_n676), 
        .ZN(DP_mult_205_n2198) );
  NAND2_X1 DP_mult_205_U1932 ( .A1(DP_mult_205_n1175), .A2(DP_mult_205_n1178), 
        .ZN(DP_mult_205_n637) );
  NAND2_X1 DP_mult_205_U1931 ( .A1(DP_mult_205_n679), .A2(DP_mult_205_n680), 
        .ZN(DP_mult_205_n341) );
  NAND2_X1 DP_mult_205_U1930 ( .A1(DP_mult_205_n681), .A2(DP_mult_205_n684), 
        .ZN(DP_mult_205_n352) );
  OR2_X1 DP_mult_205_U1929 ( .A1(DP_mult_205_n679), .A2(DP_mult_205_n680), 
        .ZN(DP_mult_205_n2197) );
  OR2_X1 DP_mult_205_U1928 ( .A1(DP_mult_205_n681), .A2(DP_mult_205_n684), 
        .ZN(DP_mult_205_n2196) );
  NOR2_X1 DP_mult_205_U1927 ( .A1(DP_mult_205_n1165), .A2(DP_mult_205_n1170), 
        .ZN(DP_mult_205_n631) );
  NOR2_X1 DP_mult_205_U1926 ( .A1(DP_mult_205_n1175), .A2(DP_mult_205_n1178), 
        .ZN(DP_mult_205_n636) );
  BUF_X1 DP_mult_205_U1925 ( .A(DP_mult_205_n2008), .Z(DP_mult_205_n2208) );
  OR2_X1 DP_mult_205_U1924 ( .A1(DP_mult_205_n685), .A2(DP_mult_205_n688), 
        .ZN(DP_mult_205_n2195) );
  OAI21_X1 DP_mult_205_U1923 ( .B1(DP_mult_205_n646), .B2(DP_mult_205_n644), 
        .A(DP_mult_205_n645), .ZN(DP_mult_205_n643) );
  AOI21_X1 DP_mult_205_U1922 ( .B1(DP_mult_205_n643), .B2(DP_mult_205_n1945), 
        .A(DP_mult_205_n1952), .ZN(DP_mult_205_n638) );
  NOR2_X1 DP_mult_205_U1921 ( .A1(DP_mult_205_n678), .A2(DP_mult_205_n677), 
        .ZN(DP_mult_205_n334) );
  INV_X1 DP_mult_205_U1920 ( .A(DP_mult_205_n341), .ZN(DP_mult_205_n339) );
  NAND2_X1 DP_mult_205_U1919 ( .A1(DP_mult_205_n678), .A2(DP_mult_205_n677), 
        .ZN(DP_mult_205_n335) );
  OAI21_X1 DP_mult_205_U1918 ( .B1(DP_mult_205_n337), .B2(DP_mult_205_n334), 
        .A(DP_mult_205_n335), .ZN(DP_mult_205_n333) );
  INV_X1 DP_mult_205_U1917 ( .A(DP_mult_205_n676), .ZN(DP_mult_205_n677) );
  XNOR2_X1 DP_mult_205_U1916 ( .A(DP_mult_205_n1124), .B(DP_mult_205_n1115), 
        .ZN(DP_mult_205_n2194) );
  XNOR2_X1 DP_mult_205_U1915 ( .A(DP_mult_205_n1113), .B(DP_mult_205_n2194), 
        .ZN(DP_mult_205_n1111) );
  NAND2_X1 DP_mult_205_U1914 ( .A1(DP_mult_205_n2228), .A2(DP_mult_205_n429), 
        .ZN(DP_mult_205_n310) );
  NAND2_X1 DP_mult_205_U1913 ( .A1(DP_mult_205_n2196), .A2(DP_mult_205_n352), 
        .ZN(DP_mult_205_n303) );
  NAND2_X1 DP_mult_205_U1912 ( .A1(DP_mult_205_n2197), .A2(DP_mult_205_n341), 
        .ZN(DP_mult_205_n302) );
  NAND2_X1 DP_mult_205_U1911 ( .A1(DP_mult_205_n2195), .A2(DP_mult_205_n369), 
        .ZN(DP_mult_205_n304) );
  NAND2_X1 DP_mult_205_U1910 ( .A1(DP_mult_205_n1958), .A2(DP_mult_205_n2190), 
        .ZN(DP_mult_205_n610) );
  NAND2_X1 DP_mult_205_U1909 ( .A1(DP_mult_205_n588), .A2(DP_mult_205_n2221), 
        .ZN(DP_mult_205_n582) );
  OR2_X1 DP_mult_205_U1908 ( .A1(DP_mult_205_n694), .A2(DP_mult_205_n689), 
        .ZN(DP_mult_205_n2193) );
  INV_X1 DP_mult_205_U1907 ( .A(DP_mult_205_n369), .ZN(DP_mult_205_n367) );
  NAND2_X1 DP_mult_205_U1906 ( .A1(DP_mult_205_n727), .A2(DP_mult_205_n736), 
        .ZN(DP_mult_205_n429) );
  NAND2_X1 DP_mult_205_U1905 ( .A1(DP_mult_205_n857), .A2(DP_mult_205_n876), 
        .ZN(DP_mult_205_n521) );
  NAND2_X1 DP_mult_205_U1904 ( .A1(DP_mult_205_n695), .A2(DP_mult_205_n700), 
        .ZN(DP_mult_205_n387) );
  OR2_X1 DP_mult_205_U1903 ( .A1(DP_mult_205_n1111), .A2(DP_mult_205_n1122), 
        .ZN(DP_mult_205_n2192) );
  OR2_X1 DP_mult_205_U1902 ( .A1(DP_mult_205_n701), .A2(DP_mult_205_n708), 
        .ZN(DP_mult_205_n2191) );
  OAI21_X1 DP_mult_205_U1901 ( .B1(DP_mult_205_n638), .B2(DP_mult_205_n636), 
        .A(DP_mult_205_n637), .ZN(DP_mult_205_n635) );
  AOI21_X1 DP_mult_205_U1900 ( .B1(DP_mult_205_n629), .B2(DP_mult_205_n635), 
        .A(DP_mult_205_n630), .ZN(DP_mult_205_n628) );
  OR2_X1 DP_mult_205_U1899 ( .A1(DP_mult_205_n1133), .A2(DP_mult_205_n1142), 
        .ZN(DP_mult_205_n2190) );
  AOI21_X1 DP_mult_205_U1898 ( .B1(DP_mult_205_n333), .B2(DP_mult_205_n1959), 
        .A(DP_mult_205_n2198), .ZN(DP_mult_205_n327) );
  AOI21_X1 DP_mult_205_U1897 ( .B1(DP_mult_205_n2190), .B2(DP_mult_205_n1947), 
        .A(DP_mult_205_n1955), .ZN(DP_mult_205_n611) );
  OR2_X1 DP_mult_205_U1896 ( .A1(DP_mult_205_n1123), .A2(DP_mult_205_n1132), 
        .ZN(DP_mult_205_n2189) );
  OAI21_X1 DP_mult_205_U1895 ( .B1(DP_mult_205_n628), .B2(DP_mult_205_n626), 
        .A(DP_mult_205_n627), .ZN(DP_mult_205_n625) );
  AOI21_X1 DP_mult_205_U1894 ( .B1(DP_mult_205_n625), .B2(DP_mult_205_n1957), 
        .A(DP_mult_205_n1948), .ZN(DP_mult_205_n620) );
  NOR2_X1 DP_mult_205_U1893 ( .A1(DP_mult_205_n336), .A2(DP_mult_205_n334), 
        .ZN(DP_mult_205_n332) );
  OR2_X1 DP_mult_205_U1892 ( .A1(DP_mult_205_n709), .A2(DP_mult_205_n716), 
        .ZN(DP_mult_205_n2188) );
  OR2_X1 DP_mult_205_U1891 ( .A1(DP_mult_205_n717), .A2(DP_mult_205_n726), 
        .ZN(DP_mult_205_n2187) );
  NOR2_X1 DP_mult_205_U1890 ( .A1(DP_mult_205_n695), .A2(DP_mult_205_n700), 
        .ZN(DP_mult_205_n384) );
  AOI21_X1 DP_mult_205_U1889 ( .B1(DP_mult_205_n2192), .B2(DP_mult_205_n1953), 
        .A(DP_mult_205_n1944), .ZN(DP_mult_205_n600) );
  AOI21_X1 DP_mult_205_U1888 ( .B1(DP_mult_205_n376), .B2(DP_mult_205_n2195), 
        .A(DP_mult_205_n367), .ZN(DP_mult_205_n365) );
  INV_X1 DP_mult_205_U1887 ( .A(DP_mult_205_n352), .ZN(DP_mult_205_n350) );
  XNOR2_X1 DP_mult_205_U1886 ( .A(DP_mult_205_n807), .B(DP_mult_205_n809), 
        .ZN(DP_mult_205_n2186) );
  XNOR2_X1 DP_mult_205_U1885 ( .A(DP_mult_205_n2186), .B(DP_mult_205_n822), 
        .ZN(DP_mult_205_n805) );
  NOR2_X1 DP_mult_205_U1884 ( .A1(DP_mult_205_n1099), .A2(DP_mult_205_n1110), 
        .ZN(DP_mult_205_n597) );
  NAND2_X1 DP_mult_205_U1883 ( .A1(DP_mult_205_n2191), .A2(DP_mult_205_n396), 
        .ZN(DP_mult_205_n307) );
  NAND2_X1 DP_mult_205_U1882 ( .A1(DP_mult_205_n2188), .A2(DP_mult_205_n409), 
        .ZN(DP_mult_205_n308) );
  OR2_X1 DP_mult_205_U1881 ( .A1(DP_mult_205_n1039), .A2(DP_mult_205_n1054), 
        .ZN(DP_mult_205_n2185) );
  INV_X1 DP_mult_205_U1880 ( .A(DP_mult_205_n396), .ZN(DP_mult_205_n394) );
  INV_X1 DP_mult_205_U1879 ( .A(DP_mult_205_n384), .ZN(DP_mult_205_n657) );
  NAND2_X1 DP_mult_205_U1878 ( .A1(DP_mult_205_n657), .A2(DP_mult_205_n387), 
        .ZN(DP_mult_205_n306) );
  OR2_X1 DP_mult_205_U1877 ( .A1(DP_mult_205_n1021), .A2(DP_mult_205_n1038), 
        .ZN(DP_mult_205_n2184) );
  INV_X1 DP_mult_205_U1876 ( .A(DP_mult_205_n378), .ZN(DP_mult_205_n376) );
  INV_X1 DP_mult_205_U1875 ( .A(DP_mult_205_n418), .ZN(DP_mult_205_n416) );
  NOR2_X1 DP_mult_205_U1874 ( .A1(DP_mult_205_n389), .A2(DP_mult_205_n384), 
        .ZN(DP_mult_205_n382) );
  OR2_X1 DP_mult_205_U1873 ( .A1(DP_mult_205_n761), .A2(DP_mult_205_n774), 
        .ZN(DP_mult_205_n2183) );
  AOI21_X1 DP_mult_205_U1872 ( .B1(DP_mult_205_n589), .B2(DP_mult_205_n2221), 
        .A(DP_mult_205_n1954), .ZN(DP_mult_205_n583) );
  OAI21_X1 DP_mult_205_U1871 ( .B1(DP_mult_205_n600), .B2(DP_mult_205_n597), 
        .A(DP_mult_205_n598), .ZN(DP_mult_205_n596) );
  OAI21_X1 DP_mult_205_U1870 ( .B1(DP_mult_205_n620), .B2(DP_mult_205_n610), 
        .A(DP_mult_205_n611), .ZN(DP_mult_205_n609) );
  NOR2_X1 DP_mult_205_U1869 ( .A1(DP_mult_205_n597), .A2(DP_mult_205_n599), 
        .ZN(DP_mult_205_n595) );
  AOI21_X1 DP_mult_205_U1868 ( .B1(DP_mult_205_n595), .B2(DP_mult_205_n609), 
        .A(DP_mult_205_n596), .ZN(DP_mult_205_n594) );
  NAND2_X1 DP_mult_205_U1867 ( .A1(DP_mult_205_n2187), .A2(DP_mult_205_n2188), 
        .ZN(DP_mult_205_n402) );
  INV_X1 DP_mult_205_U1866 ( .A(DP_mult_205_n409), .ZN(DP_mult_205_n407) );
  AOI21_X1 DP_mult_205_U1865 ( .B1(DP_mult_205_n2188), .B2(DP_mult_205_n416), 
        .A(DP_mult_205_n407), .ZN(DP_mult_205_n405) );
  NAND2_X1 DP_mult_205_U1864 ( .A1(DP_mult_205_n737), .A2(DP_mult_205_n748), 
        .ZN(DP_mult_205_n436) );
  NAND2_X1 DP_mult_205_U1863 ( .A1(DP_mult_205_n789), .A2(DP_mult_205_n804), 
        .ZN(DP_mult_205_n481) );
  INV_X1 DP_mult_205_U1862 ( .A(DP_mult_205_n564), .ZN(DP_mult_205_n562) );
  INV_X1 DP_mult_205_U1861 ( .A(DP_mult_205_n552), .ZN(DP_mult_205_n554) );
  NAND2_X1 DP_mult_205_U1860 ( .A1(DP_mult_205_n662), .A2(DP_mult_205_n436), 
        .ZN(DP_mult_205_n311) );
  INV_X1 DP_mult_205_U1859 ( .A(DP_mult_205_n563), .ZN(DP_mult_205_n561) );
  NAND2_X1 DP_mult_205_U1858 ( .A1(DP_mult_205_n663), .A2(DP_mult_205_n439), 
        .ZN(DP_mult_205_n312) );
  NOR2_X1 DP_mult_205_U1857 ( .A1(DP_mult_205_n402), .A2(DP_mult_205_n360), 
        .ZN(DP_mult_205_n356) );
  INV_X1 DP_mult_205_U1856 ( .A(DP_mult_205_n439), .ZN(DP_mult_205_n445) );
  INV_X1 DP_mult_205_U1855 ( .A(DP_mult_205_n480), .ZN(DP_mult_205_n666) );
  INV_X1 DP_mult_205_U1854 ( .A(DP_mult_205_n438), .ZN(DP_mult_205_n663) );
  INV_X1 DP_mult_205_U1853 ( .A(DP_mult_205_n383), .ZN(DP_mult_205_n381) );
  INV_X1 DP_mult_205_U1852 ( .A(DP_mult_205_n436), .ZN(DP_mult_205_n434) );
  AOI21_X1 DP_mult_205_U1851 ( .B1(DP_mult_205_n662), .B2(DP_mult_205_n445), 
        .A(DP_mult_205_n434), .ZN(DP_mult_205_n432) );
  NAND2_X1 DP_mult_205_U1850 ( .A1(DP_mult_205_n663), .A2(DP_mult_205_n662), 
        .ZN(DP_mult_205_n431) );
  INV_X1 DP_mult_205_U1849 ( .A(DP_mult_205_n481), .ZN(DP_mult_205_n483) );
  OAI21_X1 DP_mult_205_U1848 ( .B1(DP_mult_205_n492), .B2(DP_mult_205_n480), 
        .A(DP_mult_205_n481), .ZN(DP_mult_205_n479) );
  INV_X1 DP_mult_205_U1847 ( .A(DP_mult_205_n435), .ZN(DP_mult_205_n662) );
  NOR2_X1 DP_mult_205_U1846 ( .A1(DP_mult_205_n558), .A2(DP_mult_205_n563), 
        .ZN(DP_mult_205_n552) );
  INV_X1 DP_mult_205_U1845 ( .A(DP_mult_205_n420), .ZN(DP_mult_205_n422) );
  INV_X1 DP_mult_205_U1844 ( .A(DP_mult_205_n401), .ZN(DP_mult_205_n399) );
  INV_X1 DP_mult_205_U1843 ( .A(DP_mult_205_n537), .ZN(DP_mult_205_n536) );
  INV_X1 DP_mult_205_U1842 ( .A(DP_mult_205_n2102), .ZN(DP_mult_205_n2180) );
  INV_X1 DP_mult_205_U1841 ( .A(DP_mult_205_n1940), .ZN(DP_mult_205_n2178) );
  INV_X1 DP_mult_205_U1840 ( .A(DP_mult_205_n2022), .ZN(DP_mult_205_n2176) );
  INV_X1 DP_mult_205_U1839 ( .A(DP_mult_205_n2238), .ZN(DP_mult_205_n2237) );
  INV_X1 DP_mult_205_U1838 ( .A(DP_mult_205_n2238), .ZN(DP_mult_205_n2172) );
  INV_X2 DP_mult_205_U1837 ( .A(DP_mult_205_n2094), .ZN(DP_mult_205_n2171) );
  AND2_X2 DP_mult_205_U1836 ( .A1(DP_mult_205_n2232), .A2(DP_mult_205_n2231), 
        .ZN(DP_mult_205_n2230) );
  AND2_X2 DP_mult_205_U1835 ( .A1(DP_mult_205_n2232), .A2(DP_mult_205_n2231), 
        .ZN(DP_mult_205_n301) );
  XOR2_X1 DP_mult_205_U1834 ( .A(DP_coeffs_fb_int[45]), .B(
        DP_coeffs_fb_int[46]), .Z(DP_mult_205_n2201) );
  NOR2_X1 DP_mult_205_U1833 ( .A1(DP_mult_205_n877), .A2(DP_mult_205_n896), 
        .ZN(DP_mult_205_n531) );
  NOR2_X1 DP_mult_205_U1832 ( .A1(DP_mult_205_n877), .A2(DP_mult_205_n896), 
        .ZN(DP_mult_205_n2170) );
  OR2_X1 DP_mult_205_U1831 ( .A1(DP_mult_205_n876), .A2(DP_mult_205_n857), 
        .ZN(DP_mult_205_n2169) );
  NOR2_X1 DP_mult_205_U1830 ( .A1(DP_mult_205_n531), .A2(DP_mult_205_n534), 
        .ZN(DP_mult_205_n525) );
  INV_X1 DP_mult_205_U1829 ( .A(DP_mult_205_n2158), .ZN(DP_mult_205_n2168) );
  NOR2_X1 DP_mult_205_U1828 ( .A1(DP_mult_205_n502), .A2(DP_mult_205_n2122), 
        .ZN(DP_mult_205_n2167) );
  OR2_X1 DP_mult_205_U1827 ( .A1(DP_mult_205_n2108), .A2(DP_mult_205_n856), 
        .ZN(DP_mult_205_n2166) );
  INV_X2 DP_mult_205_U1826 ( .A(DP_mult_205_n2317), .ZN(DP_mult_205_n2314) );
  INV_X1 DP_mult_205_U1825 ( .A(DP_coeffs_fb_int[40]), .ZN(DP_mult_205_n2164)
         );
  XNOR2_X1 DP_mult_205_U1824 ( .A(DP_mult_205_n903), .B(DP_mult_205_n924), 
        .ZN(DP_mult_205_n2163) );
  XNOR2_X1 DP_mult_205_U1823 ( .A(DP_mult_205_n2020), .B(DP_mult_205_n2163), 
        .ZN(DP_mult_205_n899) );
  NAND3_X1 DP_mult_205_U1822 ( .A1(DP_mult_205_n2160), .A2(DP_mult_205_n2161), 
        .A3(DP_mult_205_n2162), .ZN(DP_mult_205_n974) );
  NAND2_X1 DP_mult_205_U1821 ( .A1(DP_mult_205_n1415), .A2(DP_mult_205_n1393), 
        .ZN(DP_mult_205_n2162) );
  NAND2_X1 DP_mult_205_U1820 ( .A1(DP_mult_205_n1000), .A2(DP_mult_205_n1976), 
        .ZN(DP_mult_205_n2161) );
  NAND2_X1 DP_mult_205_U1819 ( .A1(DP_mult_205_n1000), .A2(DP_mult_205_n1991), 
        .ZN(DP_mult_205_n2160) );
  XNOR2_X1 DP_mult_205_U1818 ( .A(DP_mult_205_n1393), .B(DP_mult_205_n1415), 
        .ZN(DP_mult_205_n2159) );
  XNOR2_X1 DP_mult_205_U1817 ( .A(DP_mult_205_n2159), .B(DP_mult_205_n1000), 
        .ZN(DP_mult_205_n975) );
  NOR2_X1 DP_mult_205_U1816 ( .A1(DP_mult_205_n839), .A2(DP_mult_205_n856), 
        .ZN(DP_mult_205_n513) );
  OR2_X1 DP_mult_205_U1815 ( .A1(DP_mult_205_n531), .A2(DP_mult_205_n534), 
        .ZN(DP_mult_205_n2158) );
  INV_X1 DP_mult_205_U1814 ( .A(DP_mult_205_n507), .ZN(DP_mult_205_n2157) );
  INV_X2 DP_mult_205_U1813 ( .A(DP_mult_205_n2202), .ZN(DP_mult_205_n2276) );
  NAND3_X1 DP_mult_205_U1812 ( .A1(DP_mult_205_n2153), .A2(DP_mult_205_n2154), 
        .A3(DP_mult_205_n2155), .ZN(DP_mult_205_n1022) );
  NAND2_X1 DP_mult_205_U1811 ( .A1(DP_mult_205_n1044), .A2(DP_mult_205_n1966), 
        .ZN(DP_mult_205_n2155) );
  NAND2_X1 DP_mult_205_U1810 ( .A1(DP_mult_205_n1027), .A2(DP_mult_205_n1966), 
        .ZN(DP_mult_205_n2154) );
  NAND2_X1 DP_mult_205_U1809 ( .A1(DP_mult_205_n1027), .A2(DP_mult_205_n1044), 
        .ZN(DP_mult_205_n2153) );
  NAND3_X1 DP_mult_205_U1808 ( .A1(DP_mult_205_n2150), .A2(DP_mult_205_n2151), 
        .A3(DP_mult_205_n2152), .ZN(DP_mult_205_n1042) );
  NAND2_X1 DP_mult_205_U1807 ( .A1(DP_mult_205_n1053), .A2(DP_mult_205_n1060), 
        .ZN(DP_mult_205_n2152) );
  NAND2_X1 DP_mult_205_U1806 ( .A1(DP_mult_205_n1062), .A2(DP_mult_205_n1060), 
        .ZN(DP_mult_205_n2151) );
  NAND2_X1 DP_mult_205_U1805 ( .A1(DP_mult_205_n1062), .A2(DP_mult_205_n1053), 
        .ZN(DP_mult_205_n2150) );
  XOR2_X1 DP_mult_205_U1804 ( .A(DP_mult_205_n2149), .B(DP_mult_205_n1060), 
        .Z(DP_mult_205_n1043) );
  XOR2_X1 DP_mult_205_U1803 ( .A(DP_mult_205_n1062), .B(DP_mult_205_n1053), 
        .Z(DP_mult_205_n2149) );
  OR2_X1 DP_mult_205_U1802 ( .A1(DP_mult_205_n941), .A2(DP_mult_205_n962), 
        .ZN(DP_mult_205_n2148) );
  NAND3_X1 DP_mult_205_U1801 ( .A1(DP_mult_205_n2145), .A2(DP_mult_205_n2146), 
        .A3(DP_mult_205_n2147), .ZN(DP_mult_205_n1012) );
  NAND2_X1 DP_mult_205_U1800 ( .A1(DP_mult_205_n1439), .A2(DP_mult_205_n1032), 
        .ZN(DP_mult_205_n2147) );
  NAND2_X1 DP_mult_205_U1799 ( .A1(DP_mult_205_n1036), .A2(DP_mult_205_n1032), 
        .ZN(DP_mult_205_n2146) );
  NAND2_X1 DP_mult_205_U1798 ( .A1(DP_mult_205_n1036), .A2(DP_mult_205_n1439), 
        .ZN(DP_mult_205_n2145) );
  XOR2_X1 DP_mult_205_U1797 ( .A(DP_mult_205_n2144), .B(DP_mult_205_n1032), 
        .Z(DP_mult_205_n1013) );
  XOR2_X1 DP_mult_205_U1796 ( .A(DP_mult_205_n1036), .B(DP_mult_205_n1439), 
        .Z(DP_mult_205_n2144) );
  NAND3_X1 DP_mult_205_U1795 ( .A1(DP_mult_205_n2141), .A2(DP_mult_205_n2142), 
        .A3(DP_mult_205_n2143), .ZN(DP_mult_205_n1032) );
  NAND2_X1 DP_mult_205_U1794 ( .A1(DP_mult_205_n1396), .A2(DP_mult_205_n1330), 
        .ZN(DP_mult_205_n2143) );
  NAND2_X1 DP_mult_205_U1793 ( .A1(DP_mult_205_n1463), .A2(DP_mult_205_n1330), 
        .ZN(DP_mult_205_n2142) );
  NAND2_X1 DP_mult_205_U1792 ( .A1(DP_mult_205_n1463), .A2(DP_mult_205_n1396), 
        .ZN(DP_mult_205_n2141) );
  AND2_X1 DP_mult_205_U1791 ( .A1(DP_mult_205_n1929), .A2(DP_mult_205_n876), 
        .ZN(DP_mult_205_n2140) );
  NAND3_X1 DP_mult_205_U1790 ( .A1(DP_mult_205_n2137), .A2(DP_mult_205_n2138), 
        .A3(DP_mult_205_n2139), .ZN(DP_mult_205_n954) );
  NAND2_X1 DP_mult_205_U1789 ( .A1(DP_mult_205_n1304), .A2(DP_mult_205_n1282), 
        .ZN(DP_mult_205_n2139) );
  NAND2_X1 DP_mult_205_U1788 ( .A1(DP_mult_205_n1414), .A2(DP_mult_205_n1282), 
        .ZN(DP_mult_205_n2138) );
  NAND2_X1 DP_mult_205_U1787 ( .A1(DP_mult_205_n1414), .A2(DP_mult_205_n1304), 
        .ZN(DP_mult_205_n2137) );
  XOR2_X1 DP_mult_205_U1786 ( .A(DP_mult_205_n2136), .B(DP_mult_205_n1414), 
        .Z(DP_mult_205_n955) );
  XOR2_X1 DP_mult_205_U1785 ( .A(DP_mult_205_n1282), .B(DP_mult_205_n1304), 
        .Z(DP_mult_205_n2136) );
  XNOR2_X1 DP_mult_205_U1784 ( .A(DP_mult_205_n1027), .B(DP_mult_205_n1044), 
        .ZN(DP_mult_205_n2135) );
  XNOR2_X1 DP_mult_205_U1783 ( .A(DP_mult_205_n2135), .B(DP_mult_205_n1042), 
        .ZN(DP_mult_205_n1023) );
  INV_X1 DP_mult_205_U1782 ( .A(DP_mult_205_n2277), .ZN(DP_mult_205_n2134) );
  NAND3_X1 DP_mult_205_U1781 ( .A1(DP_mult_205_n2131), .A2(DP_mult_205_n2132), 
        .A3(DP_mult_205_n2133), .ZN(DP_mult_205_n856) );
  NAND2_X1 DP_mult_205_U1780 ( .A1(DP_mult_205_n878), .A2(DP_mult_205_n861), 
        .ZN(DP_mult_205_n2133) );
  NAND2_X1 DP_mult_205_U1779 ( .A1(DP_mult_205_n859), .A2(DP_mult_205_n861), 
        .ZN(DP_mult_205_n2132) );
  NAND2_X1 DP_mult_205_U1778 ( .A1(DP_mult_205_n859), .A2(DP_mult_205_n878), 
        .ZN(DP_mult_205_n2131) );
  INV_X2 DP_mult_205_U1777 ( .A(DP_mult_205_n2082), .ZN(DP_mult_205_n2253) );
  BUF_X2 DP_mult_205_U1776 ( .A(DP_mult_205_n287), .Z(DP_mult_205_n2130) );
  NAND3_X1 DP_mult_205_U1775 ( .A1(DP_mult_205_n2127), .A2(DP_mult_205_n2128), 
        .A3(DP_mult_205_n2129), .ZN(DP_mult_205_n884) );
  NAND2_X1 DP_mult_205_U1774 ( .A1(DP_mult_205_n891), .A2(DP_mult_205_n895), 
        .ZN(DP_mult_205_n2129) );
  NAND2_X1 DP_mult_205_U1773 ( .A1(DP_mult_205_n908), .A2(DP_mult_205_n895), 
        .ZN(DP_mult_205_n2128) );
  NAND2_X1 DP_mult_205_U1772 ( .A1(DP_mult_205_n908), .A2(DP_mult_205_n891), 
        .ZN(DP_mult_205_n2127) );
  XOR2_X1 DP_mult_205_U1771 ( .A(DP_mult_205_n908), .B(DP_mult_205_n2126), .Z(
        DP_mult_205_n885) );
  XOR2_X1 DP_mult_205_U1770 ( .A(DP_mult_205_n891), .B(DP_mult_205_n895), .Z(
        DP_mult_205_n2126) );
  INV_X1 DP_mult_205_U1769 ( .A(DP_mult_205_n2101), .ZN(DP_mult_205_n2179) );
  NAND3_X1 DP_mult_205_U1768 ( .A1(DP_mult_205_n2123), .A2(DP_mult_205_n2124), 
        .A3(DP_mult_205_n2125), .ZN(DP_mult_205_n820) );
  NAND2_X1 DP_mult_205_U1767 ( .A1(DP_mult_205_n840), .A2(DP_mult_205_n825), 
        .ZN(DP_mult_205_n2125) );
  NAND2_X1 DP_mult_205_U1766 ( .A1(DP_mult_205_n823), .A2(DP_mult_205_n825), 
        .ZN(DP_mult_205_n2124) );
  NAND2_X1 DP_mult_205_U1765 ( .A1(DP_mult_205_n823), .A2(DP_mult_205_n840), 
        .ZN(DP_mult_205_n2123) );
  NOR2_X1 DP_mult_205_U1764 ( .A1(DP_mult_205_n805), .A2(DP_mult_205_n820), 
        .ZN(DP_mult_205_n2122) );
  NAND3_X1 DP_mult_205_U1763 ( .A1(DP_mult_205_n2119), .A2(DP_mult_205_n2120), 
        .A3(DP_mult_205_n2121), .ZN(DP_mult_205_n846) );
  NAND2_X1 DP_mult_205_U1762 ( .A1(DP_mult_205_n868), .A2(DP_mult_205_n870), 
        .ZN(DP_mult_205_n2121) );
  NAND2_X1 DP_mult_205_U1761 ( .A1(DP_mult_205_n851), .A2(DP_mult_205_n870), 
        .ZN(DP_mult_205_n2120) );
  NAND2_X1 DP_mult_205_U1760 ( .A1(DP_mult_205_n851), .A2(DP_mult_205_n868), 
        .ZN(DP_mult_205_n2119) );
  XOR2_X1 DP_mult_205_U1759 ( .A(DP_mult_205_n851), .B(DP_mult_205_n2118), .Z(
        DP_mult_205_n847) );
  XOR2_X1 DP_mult_205_U1758 ( .A(DP_mult_205_n868), .B(DP_mult_205_n870), .Z(
        DP_mult_205_n2118) );
  XNOR2_X1 DP_mult_205_U1757 ( .A(DP_mult_205_n878), .B(DP_mult_205_n861), 
        .ZN(DP_mult_205_n2117) );
  XNOR2_X1 DP_mult_205_U1756 ( .A(DP_mult_205_n859), .B(DP_mult_205_n2117), 
        .ZN(DP_mult_205_n857) );
  NAND3_X1 DP_mult_205_U1755 ( .A1(DP_mult_205_n2114), .A2(DP_mult_205_n2116), 
        .A3(DP_mult_205_n2115), .ZN(DP_mult_205_n834) );
  NAND2_X1 DP_mult_205_U1754 ( .A1(DP_mult_205_n1210), .A2(DP_mult_205_n1276), 
        .ZN(DP_mult_205_n2116) );
  NAND2_X1 DP_mult_205_U1753 ( .A1(DP_mult_205_n837), .A2(DP_mult_205_n1276), 
        .ZN(DP_mult_205_n2115) );
  NAND2_X1 DP_mult_205_U1752 ( .A1(DP_mult_205_n837), .A2(DP_mult_205_n1210), 
        .ZN(DP_mult_205_n2114) );
  XOR2_X1 DP_mult_205_U1751 ( .A(DP_mult_205_n1977), .B(DP_mult_205_n2113), 
        .Z(DP_mult_205_n835) );
  XOR2_X1 DP_mult_205_U1750 ( .A(DP_mult_205_n1210), .B(DP_mult_205_n1276), 
        .Z(DP_mult_205_n2113) );
  NAND3_X1 DP_mult_205_U1749 ( .A1(DP_mult_205_n2110), .A2(DP_mult_205_n2111), 
        .A3(DP_mult_205_n2112), .ZN(DP_mult_205_n922) );
  NAND2_X1 DP_mult_205_U1748 ( .A1(DP_mult_205_n948), .A2(DP_mult_205_n929), 
        .ZN(DP_mult_205_n2112) );
  NAND2_X1 DP_mult_205_U1747 ( .A1(DP_mult_205_n946), .A2(DP_mult_205_n929), 
        .ZN(DP_mult_205_n2111) );
  NAND2_X1 DP_mult_205_U1746 ( .A1(DP_mult_205_n946), .A2(DP_mult_205_n948), 
        .ZN(DP_mult_205_n2110) );
  XOR2_X1 DP_mult_205_U1745 ( .A(DP_mult_205_n2057), .B(DP_mult_205_n2109), 
        .Z(DP_mult_205_n923) );
  XOR2_X1 DP_mult_205_U1744 ( .A(DP_mult_205_n948), .B(DP_mult_205_n929), .Z(
        DP_mult_205_n2109) );
  INV_X1 DP_mult_205_U1743 ( .A(DP_coeffs_fb_int[42]), .ZN(DP_mult_205_n2293)
         );
  CLKBUF_X1 DP_mult_205_U1742 ( .A(DP_mult_205_n839), .Z(DP_mult_205_n2108) );
  INV_X1 DP_mult_205_U1741 ( .A(DP_mult_205_n2254), .ZN(DP_mult_205_n2107) );
  NOR2_X1 DP_mult_205_U1740 ( .A1(DP_mult_205_n941), .A2(DP_mult_205_n962), 
        .ZN(DP_mult_205_n547) );
  INV_X4 DP_mult_205_U1739 ( .A(DP_mult_205_n1939), .ZN(DP_mult_205_n2326) );
  INV_X1 DP_mult_205_U1738 ( .A(DP_mult_205_n2290), .ZN(DP_mult_205_n2106) );
  INV_X1 DP_mult_205_U1737 ( .A(DP_mult_205_n554), .ZN(DP_mult_205_n2105) );
  INV_X2 DP_mult_205_U1736 ( .A(DP_mult_205_n2305), .ZN(DP_mult_205_n2303) );
  INV_X1 DP_mult_205_U1735 ( .A(DP_mult_205_n2302), .ZN(DP_mult_205_n2104) );
  XOR2_X1 DP_mult_205_U1734 ( .A(DP_mult_205_n1238), .B(DP_mult_205_n1216), 
        .Z(DP_mult_205_n961) );
  OR2_X2 DP_mult_205_U1733 ( .A1(DP_mult_205_n775), .A2(DP_mult_205_n788), 
        .ZN(DP_mult_205_n2182) );
  AND2_X1 DP_mult_205_U1732 ( .A1(DP_mult_205_n1809), .A2(DP_mult_205_n2261), 
        .ZN(DP_mult_205_n2101) );
  INV_X2 DP_mult_205_U1731 ( .A(DP_mult_205_n2309), .ZN(DP_mult_205_n2308) );
  INV_X1 DP_mult_205_U1730 ( .A(DP_mult_205_n2246), .ZN(DP_mult_205_n2245) );
  INV_X1 DP_mult_205_U1729 ( .A(DP_mult_205_n2246), .ZN(DP_mult_205_n2099) );
  INV_X1 DP_mult_205_U1728 ( .A(DP_mult_205_n2246), .ZN(DP_mult_205_n2100) );
  NOR2_X1 DP_mult_205_U1727 ( .A1(DP_mult_205_n941), .A2(DP_mult_205_n962), 
        .ZN(DP_mult_205_n2098) );
  NOR2_X1 DP_mult_205_U1726 ( .A1(DP_mult_205_n2098), .A2(DP_mult_205_n542), 
        .ZN(DP_mult_205_n2097) );
  INV_X2 DP_mult_205_U1725 ( .A(DP_mult_205_n2293), .ZN(DP_mult_205_n2292) );
  INV_X1 DP_mult_205_U1724 ( .A(DP_mult_205_n2093), .ZN(DP_mult_205_n2248) );
  INV_X1 DP_mult_205_U1723 ( .A(DP_mult_205_n2093), .ZN(DP_mult_205_n2095) );
  INV_X1 DP_mult_205_U1722 ( .A(DP_mult_205_n2093), .ZN(DP_mult_205_n2096) );
  AND2_X1 DP_mult_205_U1721 ( .A1(DP_mult_205_n1814), .A2(DP_mult_205_n2030), 
        .ZN(DP_mult_205_n2094) );
  AND2_X1 DP_mult_205_U1720 ( .A1(DP_mult_205_n1814), .A2(DP_mult_205_n2030), 
        .ZN(DP_mult_205_n2093) );
  INV_X1 DP_mult_205_U1719 ( .A(DP_mult_205_n2203), .ZN(DP_mult_205_n2258) );
  INV_X2 DP_mult_205_U1718 ( .A(DP_mult_205_n1971), .ZN(DP_mult_205_n2235) );
  NAND3_X1 DP_mult_205_U1717 ( .A1(DP_mult_205_n2090), .A2(DP_mult_205_n2091), 
        .A3(DP_mult_205_n2092), .ZN(DP_mult_205_n796) );
  NAND2_X1 DP_mult_205_U1716 ( .A1(DP_mult_205_n1296), .A2(DP_mult_205_n818), 
        .ZN(DP_mult_205_n2092) );
  NAND2_X1 DP_mult_205_U1715 ( .A1(DP_mult_205_n1274), .A2(DP_mult_205_n818), 
        .ZN(DP_mult_205_n2091) );
  NAND2_X1 DP_mult_205_U1714 ( .A1(DP_mult_205_n1274), .A2(DP_mult_205_n1296), 
        .ZN(DP_mult_205_n2090) );
  XOR2_X1 DP_mult_205_U1713 ( .A(DP_mult_205_n2089), .B(DP_mult_205_n818), .Z(
        DP_mult_205_n797) );
  XOR2_X1 DP_mult_205_U1712 ( .A(DP_mult_205_n1274), .B(DP_mult_205_n1296), 
        .Z(DP_mult_205_n2089) );
  NAND3_X1 DP_mult_205_U1711 ( .A1(DP_mult_205_n2086), .A2(DP_mult_205_n2087), 
        .A3(DP_mult_205_n2088), .ZN(DP_mult_205_n818) );
  NAND2_X1 DP_mult_205_U1710 ( .A1(DP_mult_205_n1209), .A2(DP_mult_205_n2165), 
        .ZN(DP_mult_205_n2088) );
  NAND2_X1 DP_mult_205_U1709 ( .A1(DP_mult_205_n1363), .A2(DP_mult_205_n2165), 
        .ZN(DP_mult_205_n2087) );
  NAND2_X1 DP_mult_205_U1708 ( .A1(DP_mult_205_n1363), .A2(DP_mult_205_n1209), 
        .ZN(DP_mult_205_n2086) );
  XOR2_X1 DP_mult_205_U1707 ( .A(DP_mult_205_n2085), .B(DP_mult_205_n2165), 
        .Z(DP_mult_205_n819) );
  XOR2_X1 DP_mult_205_U1706 ( .A(DP_mult_205_n1209), .B(DP_mult_205_n1363), 
        .Z(DP_mult_205_n2085) );
  INV_X2 DP_mult_205_U1705 ( .A(DP_mult_205_n2102), .ZN(DP_mult_205_n2239) );
  INV_X1 DP_mult_205_U1704 ( .A(DP_mult_205_n2286), .ZN(DP_mult_205_n2283) );
  BUF_X2 DP_mult_205_U1703 ( .A(DP_mult_205_n251), .Z(DP_mult_205_n2280) );
  NAND2_X1 DP_mult_205_U1702 ( .A1(DP_mult_205_n2083), .A2(DP_mult_205_n2084), 
        .ZN(DP_mult_205_n1459) );
  OR2_X1 DP_mult_205_U1701 ( .A1(DP_mult_205_n1757), .A2(DP_mult_205_n2280), 
        .ZN(DP_mult_205_n2084) );
  OR2_X1 DP_mult_205_U1700 ( .A1(DP_mult_205_n1949), .A2(DP_mult_205_n1758), 
        .ZN(DP_mult_205_n2083) );
  AND2_X1 DP_mult_205_U1699 ( .A1(DP_mult_205_n1817), .A2(DP_mult_205_n2280), 
        .ZN(DP_mult_205_n2082) );
  OAI21_X1 DP_mult_205_U1698 ( .B1(DP_mult_205_n503), .B2(DP_mult_205_n2122), 
        .A(DP_mult_205_n496), .ZN(DP_mult_205_n2081) );
  BUF_X1 DP_mult_205_U1697 ( .A(DP_mult_205_n532), .Z(DP_mult_205_n2080) );
  INV_X1 DP_mult_205_U1696 ( .A(DP_mult_205_n1972), .ZN(DP_mult_205_n2241) );
  INV_X1 DP_mult_205_U1695 ( .A(DP_mult_205_n1972), .ZN(DP_mult_205_n2078) );
  INV_X1 DP_mult_205_U1694 ( .A(DP_mult_205_n1972), .ZN(DP_mult_205_n2079) );
  NAND3_X1 DP_mult_205_U1693 ( .A1(DP_mult_205_n2075), .A2(DP_mult_205_n2076), 
        .A3(DP_mult_205_n2077), .ZN(DP_mult_205_n806) );
  NAND2_X1 DP_mult_205_U1692 ( .A1(DP_mult_205_n811), .A2(DP_mult_205_n826), 
        .ZN(DP_mult_205_n2077) );
  NAND2_X1 DP_mult_205_U1691 ( .A1(DP_mult_205_n824), .A2(DP_mult_205_n826), 
        .ZN(DP_mult_205_n2076) );
  NAND2_X1 DP_mult_205_U1690 ( .A1(DP_mult_205_n824), .A2(DP_mult_205_n811), 
        .ZN(DP_mult_205_n2075) );
  INV_X1 DP_mult_205_U1689 ( .A(DP_mult_205_n2200), .ZN(DP_mult_205_n2269) );
  CLKBUF_X1 DP_mult_205_U1688 ( .A(DP_mult_205_n547), .Z(DP_mult_205_n2074) );
  CLKBUF_X3 DP_mult_205_U1687 ( .A(DP_mult_205_n277), .Z(DP_mult_205_n2073) );
  AOI21_X1 DP_mult_205_U1686 ( .B1(DP_mult_205_n581), .B2(DP_mult_205_n567), 
        .A(DP_mult_205_n568), .ZN(DP_mult_205_n2072) );
  XNOR2_X1 DP_mult_205_U1685 ( .A(DP_mult_205_n840), .B(DP_mult_205_n825), 
        .ZN(DP_mult_205_n2071) );
  XNOR2_X1 DP_mult_205_U1684 ( .A(DP_mult_205_n823), .B(DP_mult_205_n2071), 
        .ZN(DP_mult_205_n821) );
  INV_X1 DP_mult_205_U1683 ( .A(DP_mult_205_n2298), .ZN(DP_mult_205_n2070) );
  OR2_X1 DP_mult_205_U1682 ( .A1(DP_mult_205_n877), .A2(DP_mult_205_n896), 
        .ZN(DP_mult_205_n2069) );
  BUF_X1 DP_mult_205_U1681 ( .A(DP_mult_205_n1285), .Z(DP_mult_205_n2068) );
  NAND3_X1 DP_mult_205_U1680 ( .A1(DP_mult_205_n2065), .A2(DP_mult_205_n2066), 
        .A3(DP_mult_205_n2067), .ZN(DP_mult_205_n992) );
  NAND2_X1 DP_mult_205_U1679 ( .A1(DP_mult_205_n1001), .A2(DP_mult_205_n1018), 
        .ZN(DP_mult_205_n2067) );
  NAND2_X1 DP_mult_205_U1678 ( .A1(DP_mult_205_n1394), .A2(DP_mult_205_n1935), 
        .ZN(DP_mult_205_n2066) );
  NAND2_X1 DP_mult_205_U1677 ( .A1(DP_mult_205_n1394), .A2(DP_mult_205_n1001), 
        .ZN(DP_mult_205_n2065) );
  XOR2_X1 DP_mult_205_U1676 ( .A(DP_mult_205_n2064), .B(DP_mult_205_n1018), 
        .Z(DP_mult_205_n993) );
  XOR2_X1 DP_mult_205_U1675 ( .A(DP_mult_205_n1394), .B(DP_mult_205_n1001), 
        .Z(DP_mult_205_n2064) );
  NAND3_X1 DP_mult_205_U1674 ( .A1(DP_mult_205_n2061), .A2(DP_mult_205_n2062), 
        .A3(DP_mult_205_n2063), .ZN(DP_mult_205_n1018) );
  NAND2_X1 DP_mult_205_U1673 ( .A1(DP_mult_205_n1263), .A2(DP_mult_205_n1285), 
        .ZN(DP_mult_205_n2063) );
  NAND2_X1 DP_mult_205_U1672 ( .A1(DP_mult_205_n1351), .A2(DP_mult_205_n1285), 
        .ZN(DP_mult_205_n2062) );
  NAND2_X1 DP_mult_205_U1671 ( .A1(DP_mult_205_n1351), .A2(DP_mult_205_n1263), 
        .ZN(DP_mult_205_n2061) );
  XOR2_X1 DP_mult_205_U1670 ( .A(DP_mult_205_n2060), .B(DP_mult_205_n2068), 
        .Z(DP_mult_205_n1019) );
  XOR2_X1 DP_mult_205_U1669 ( .A(DP_mult_205_n1351), .B(DP_mult_205_n1263), 
        .Z(DP_mult_205_n2060) );
  INV_X1 DP_mult_205_U1668 ( .A(DP_mult_205_n1960), .ZN(DP_mult_205_n2266) );
  NOR2_X1 DP_mult_205_U1667 ( .A1(DP_mult_205_n839), .A2(DP_mult_205_n856), 
        .ZN(DP_mult_205_n2059) );
  INV_X1 DP_mult_205_U1666 ( .A(DP_mult_205_n2156), .ZN(DP_mult_205_n2202) );
  INV_X1 DP_mult_205_U1665 ( .A(DP_mult_205_n2069), .ZN(DP_mult_205_n2058) );
  CLKBUF_X1 DP_mult_205_U1664 ( .A(DP_mult_205_n946), .Z(DP_mult_205_n2057) );
  NAND3_X1 DP_mult_205_U1663 ( .A1(DP_mult_205_n2054), .A2(DP_mult_205_n2055), 
        .A3(DP_mult_205_n2056), .ZN(DP_mult_205_n970) );
  NAND2_X1 DP_mult_205_U1662 ( .A1(DP_mult_205_n979), .A2(DP_mult_205_n977), 
        .ZN(DP_mult_205_n2056) );
  NAND2_X1 DP_mult_205_U1661 ( .A1(DP_mult_205_n998), .A2(DP_mult_205_n977), 
        .ZN(DP_mult_205_n2055) );
  NAND2_X1 DP_mult_205_U1660 ( .A1(DP_mult_205_n998), .A2(DP_mult_205_n979), 
        .ZN(DP_mult_205_n2054) );
  NAND3_X1 DP_mult_205_U1659 ( .A1(DP_mult_205_n2051), .A2(DP_mult_205_n2052), 
        .A3(DP_mult_205_n2053), .ZN(DP_mult_205_n976) );
  NAND2_X1 DP_mult_205_U1658 ( .A1(DP_mult_205_n1437), .A2(DP_mult_205_n1327), 
        .ZN(DP_mult_205_n2053) );
  NAND2_X1 DP_mult_205_U1657 ( .A1(DP_mult_205_n1305), .A2(DP_mult_205_n1327), 
        .ZN(DP_mult_205_n2052) );
  NAND2_X1 DP_mult_205_U1656 ( .A1(DP_mult_205_n1305), .A2(DP_mult_205_n1437), 
        .ZN(DP_mult_205_n2051) );
  XOR2_X1 DP_mult_205_U1655 ( .A(DP_mult_205_n2050), .B(DP_mult_205_n977), .Z(
        DP_mult_205_n971) );
  XOR2_X1 DP_mult_205_U1654 ( .A(DP_mult_205_n998), .B(DP_mult_205_n979), .Z(
        DP_mult_205_n2050) );
  NAND3_X1 DP_mult_205_U1653 ( .A1(DP_mult_205_n2046), .A2(DP_mult_205_n2047), 
        .A3(DP_mult_205_n2048), .ZN(DP_mult_205_n940) );
  NAND2_X1 DP_mult_205_U1652 ( .A1(DP_mult_205_n964), .A2(DP_mult_205_n945), 
        .ZN(DP_mult_205_n2048) );
  NAND2_X1 DP_mult_205_U1651 ( .A1(DP_mult_205_n943), .A2(DP_mult_205_n945), 
        .ZN(DP_mult_205_n2047) );
  NAND2_X1 DP_mult_205_U1650 ( .A1(DP_mult_205_n943), .A2(DP_mult_205_n964), 
        .ZN(DP_mult_205_n2046) );
  BUF_X1 DP_mult_205_U1649 ( .A(DP_mult_205_n550), .Z(DP_mult_205_n2045) );
  XNOR2_X1 DP_mult_205_U1648 ( .A(DP_coeffs_fb_int[31]), .B(DP_mult_205_n2317), 
        .ZN(DP_mult_205_n1809) );
  INV_X1 DP_mult_205_U1647 ( .A(DP_coeffs_fb_int[38]), .ZN(DP_mult_205_n2044)
         );
  INV_X1 DP_mult_205_U1646 ( .A(DP_mult_205_n2201), .ZN(DP_mult_205_n2277) );
  INV_X1 DP_mult_205_U1645 ( .A(DP_mult_205_n2041), .ZN(DP_mult_205_n2042) );
  INV_X1 DP_mult_205_U1644 ( .A(DP_mult_205_n2156), .ZN(DP_mult_205_n2041) );
  INV_X2 DP_mult_205_U1643 ( .A(DP_mult_205_n2312), .ZN(DP_mult_205_n2311) );
  INV_X2 DP_mult_205_U1642 ( .A(DP_mult_205_n2312), .ZN(DP_mult_205_n2310) );
  NAND3_X1 DP_mult_205_U1641 ( .A1(DP_mult_205_n2038), .A2(DP_mult_205_n2039), 
        .A3(DP_mult_205_n2040), .ZN(DP_mult_205_n1058) );
  NAND2_X1 DP_mult_205_U1640 ( .A1(DP_mult_205_n1067), .A2(DP_mult_205_n1065), 
        .ZN(DP_mult_205_n2040) );
  NAND2_X1 DP_mult_205_U1639 ( .A1(DP_mult_205_n1076), .A2(DP_mult_205_n1065), 
        .ZN(DP_mult_205_n2039) );
  NAND2_X1 DP_mult_205_U1638 ( .A1(DP_mult_205_n1076), .A2(DP_mult_205_n1067), 
        .ZN(DP_mult_205_n2038) );
  XOR2_X1 DP_mult_205_U1637 ( .A(DP_mult_205_n1970), .B(DP_mult_205_n2037), 
        .Z(DP_mult_205_n1059) );
  XOR2_X1 DP_mult_205_U1636 ( .A(DP_mult_205_n1067), .B(DP_mult_205_n1065), 
        .Z(DP_mult_205_n2037) );
  XNOR2_X1 DP_mult_205_U1635 ( .A(DP_coeffs_fb_int[43]), .B(
        DP_coeffs_fb_int[44]), .ZN(DP_mult_205_n2156) );
  BUF_X2 DP_mult_205_U1634 ( .A(DP_mult_205_n283), .Z(DP_mult_205_n2174) );
  INV_X2 DP_mult_205_U1633 ( .A(DP_mult_205_n2207), .ZN(DP_mult_205_n2236) );
  NOR2_X1 DP_mult_205_U1632 ( .A1(DP_mult_205_n513), .A2(DP_mult_205_n520), 
        .ZN(DP_mult_205_n2036) );
  NAND3_X1 DP_mult_205_U1631 ( .A1(DP_mult_205_n2033), .A2(DP_mult_205_n2034), 
        .A3(DP_mult_205_n2035), .ZN(DP_mult_205_n956) );
  NAND2_X1 DP_mult_205_U1630 ( .A1(DP_mult_205_n1459), .A2(DP_mult_205_n1436), 
        .ZN(DP_mult_205_n2035) );
  NAND2_X1 DP_mult_205_U1629 ( .A1(DP_mult_205_n1370), .A2(DP_mult_205_n1436), 
        .ZN(DP_mult_205_n2034) );
  NAND2_X1 DP_mult_205_U1628 ( .A1(DP_mult_205_n1370), .A2(DP_mult_205_n1459), 
        .ZN(DP_mult_205_n2033) );
  XOR2_X1 DP_mult_205_U1627 ( .A(DP_mult_205_n2032), .B(DP_mult_205_n1370), 
        .Z(DP_mult_205_n957) );
  XOR2_X1 DP_mult_205_U1626 ( .A(DP_mult_205_n1459), .B(DP_mult_205_n1436), 
        .Z(DP_mult_205_n2032) );
  INV_X1 DP_mult_205_U1625 ( .A(DP_mult_205_n2321), .ZN(DP_mult_205_n2319) );
  INV_X1 DP_mult_205_U1624 ( .A(DP_mult_205_n2293), .ZN(DP_mult_205_n2291) );
  CLKBUF_X1 DP_mult_205_U1623 ( .A(DP_mult_205_n535), .Z(DP_mult_205_n2031) );
  NAND2_X1 DP_mult_205_U1622 ( .A1(DP_mult_205_n2028), .A2(DP_mult_205_n2029), 
        .ZN(DP_mult_205_n1320) );
  OR2_X1 DP_mult_205_U1621 ( .A1(DP_mult_205_n1613), .A2(DP_mult_205_n2267), 
        .ZN(DP_mult_205_n2029) );
  OR2_X1 DP_mult_205_U1620 ( .A1(DP_mult_205_n2242), .A2(DP_mult_205_n1614), 
        .ZN(DP_mult_205_n2028) );
  NAND3_X1 DP_mult_205_U1619 ( .A1(DP_mult_205_n2025), .A2(DP_mult_205_n2026), 
        .A3(DP_mult_205_n2027), .ZN(DP_mult_205_n830) );
  NAND2_X1 DP_mult_205_U1618 ( .A1(DP_mult_205_n1254), .A2(DP_mult_205_n1298), 
        .ZN(DP_mult_205_n2027) );
  NAND2_X1 DP_mult_205_U1617 ( .A1(DP_mult_205_n1298), .A2(DP_mult_205_n1320), 
        .ZN(DP_mult_205_n2026) );
  NAND2_X1 DP_mult_205_U1616 ( .A1(DP_mult_205_n2001), .A2(DP_mult_205_n1254), 
        .ZN(DP_mult_205_n2025) );
  XOR2_X1 DP_mult_205_U1615 ( .A(DP_mult_205_n2001), .B(DP_mult_205_n2024), 
        .Z(DP_mult_205_n831) );
  XOR2_X1 DP_mult_205_U1614 ( .A(DP_mult_205_n1298), .B(DP_mult_205_n1254), 
        .Z(DP_mult_205_n2024) );
  XOR2_X1 DP_mult_205_U1613 ( .A(DP_coeffs_fb_int[37]), .B(
        DP_coeffs_fb_int[38]), .Z(DP_mult_205_n2200) );
  INV_X1 DP_mult_205_U1612 ( .A(DP_mult_205_n2269), .ZN(DP_mult_205_n2023) );
  AND2_X1 DP_mult_205_U1611 ( .A1(DP_mult_205_n1812), .A2(DP_mult_205_n2269), 
        .ZN(DP_mult_205_n2021) );
  NAND3_X1 DP_mult_205_U1610 ( .A1(DP_mult_205_n2110), .A2(DP_mult_205_n2111), 
        .A3(DP_mult_205_n2112), .ZN(DP_mult_205_n2019) );
  NAND3_X1 DP_mult_205_U1609 ( .A1(DP_mult_205_n2110), .A2(DP_mult_205_n2111), 
        .A3(DP_mult_205_n2112), .ZN(DP_mult_205_n2020) );
  XNOR2_X1 DP_mult_205_U1608 ( .A(DP_mult_205_n1463), .B(DP_mult_205_n1396), 
        .ZN(DP_mult_205_n2018) );
  XNOR2_X1 DP_mult_205_U1607 ( .A(DP_mult_205_n2018), .B(DP_mult_205_n1938), 
        .ZN(DP_mult_205_n1033) );
  INV_X2 DP_mult_205_U1606 ( .A(DP_mult_205_n2206), .ZN(DP_mult_205_n2255) );
  INV_X2 DP_mult_205_U1605 ( .A(DP_mult_205_n2206), .ZN(DP_mult_205_n2254) );
  OAI22_X1 DP_mult_205_U1604 ( .A1(DP_mult_205_n1987), .A2(DP_mult_205_n1733), 
        .B1(DP_mult_205_n1732), .B2(DP_mult_205_n2278), .ZN(DP_mult_205_n2017)
         );
  XNOR2_X1 DP_mult_205_U1603 ( .A(DP_coeffs_fb_int[35]), .B(DP_mult_205_n2309), 
        .ZN(DP_mult_205_n1811) );
  INV_X1 DP_mult_205_U1602 ( .A(DP_mult_205_n2297), .ZN(DP_mult_205_n2015) );
  INV_X1 DP_mult_205_U1601 ( .A(DP_mult_205_n2297), .ZN(DP_mult_205_n2016) );
  INV_X1 DP_mult_205_U1600 ( .A(DP_mult_205_n2293), .ZN(DP_mult_205_n2290) );
  INV_X1 DP_mult_205_U1599 ( .A(DP_mult_205_n2328), .ZN(DP_mult_205_n2327) );
  NAND3_X1 DP_mult_205_U1598 ( .A1(DP_mult_205_n2012), .A2(DP_mult_205_n2013), 
        .A3(DP_mult_205_n2014), .ZN(DP_mult_205_n962) );
  NAND2_X1 DP_mult_205_U1597 ( .A1(DP_mult_205_n984), .A2(DP_mult_205_n967), 
        .ZN(DP_mult_205_n2014) );
  NAND2_X1 DP_mult_205_U1596 ( .A1(DP_mult_205_n965), .A2(DP_mult_205_n967), 
        .ZN(DP_mult_205_n2013) );
  NAND2_X1 DP_mult_205_U1595 ( .A1(DP_mult_205_n965), .A2(DP_mult_205_n984), 
        .ZN(DP_mult_205_n2012) );
  XNOR2_X1 DP_mult_205_U1594 ( .A(DP_coeffs_fb_int[45]), .B(DP_mult_205_n2289), 
        .ZN(DP_mult_205_n1816) );
  INV_X1 DP_mult_205_U1593 ( .A(DP_mult_205_n2275), .ZN(DP_mult_205_n2272) );
  XNOR2_X1 DP_mult_205_U1592 ( .A(DP_mult_205_n811), .B(DP_mult_205_n826), 
        .ZN(DP_mult_205_n2011) );
  XNOR2_X1 DP_mult_205_U1591 ( .A(DP_mult_205_n824), .B(DP_mult_205_n2011), 
        .ZN(DP_mult_205_n807) );
  NOR2_X1 DP_mult_205_U1590 ( .A1(DP_mult_205_n456), .A2(DP_mult_205_n480), 
        .ZN(DP_mult_205_n2010) );
  XNOR2_X1 DP_mult_205_U1589 ( .A(DP_mult_205_n984), .B(DP_mult_205_n967), 
        .ZN(DP_mult_205_n2009) );
  XNOR2_X1 DP_mult_205_U1588 ( .A(DP_mult_205_n965), .B(DP_mult_205_n2009), 
        .ZN(DP_mult_205_n963) );
  INV_X1 DP_mult_205_U1587 ( .A(DP_mult_205_n2008), .ZN(DP_mult_205_n2204) );
  XNOR2_X1 DP_mult_205_U1586 ( .A(DP_coeffs_fb_int[27]), .B(
        DP_coeffs_fb_int[28]), .ZN(DP_mult_205_n2008) );
  CLKBUF_X3 DP_mult_205_U1585 ( .A(DP_mult_205_n293), .Z(DP_mult_205_n2103) );
  INV_X1 DP_mult_205_U1584 ( .A(DP_mult_205_n1985), .ZN(DP_mult_205_n2173) );
  XNOR2_X1 DP_mult_205_U1583 ( .A(DP_coeffs_fb_int[43]), .B(DP_mult_205_n2293), 
        .ZN(DP_mult_205_n1815) );
  INV_X1 DP_mult_205_U1582 ( .A(DP_mult_205_n2322), .ZN(DP_mult_205_n2007) );
  INV_X1 DP_mult_205_U1581 ( .A(DP_mult_205_n1961), .ZN(DP_mult_205_n2267) );
  INV_X1 DP_mult_205_U1580 ( .A(DP_mult_205_n2041), .ZN(DP_mult_205_n2043) );
  NAND3_X1 DP_mult_205_U1579 ( .A1(DP_mult_205_n2003), .A2(DP_mult_205_n2004), 
        .A3(DP_mult_205_n2005), .ZN(DP_mult_205_n958) );
  NAND2_X1 DP_mult_205_U1578 ( .A1(DP_mult_205_n1348), .A2(DP_mult_205_n1182), 
        .ZN(DP_mult_205_n2005) );
  NAND2_X1 DP_mult_205_U1577 ( .A1(DP_mult_205_n1260), .A2(DP_mult_205_n1182), 
        .ZN(DP_mult_205_n2004) );
  NAND2_X1 DP_mult_205_U1576 ( .A1(DP_mult_205_n1260), .A2(DP_mult_205_n1348), 
        .ZN(DP_mult_205_n2003) );
  XOR2_X1 DP_mult_205_U1575 ( .A(DP_mult_205_n2002), .B(DP_mult_205_n1260), 
        .Z(DP_mult_205_n959) );
  XOR2_X1 DP_mult_205_U1574 ( .A(DP_mult_205_n1182), .B(DP_mult_205_n1348), 
        .Z(DP_mult_205_n2002) );
  NAND2_X1 DP_mult_205_U1573 ( .A1(DP_mult_205_n2028), .A2(DP_mult_205_n2029), 
        .ZN(DP_mult_205_n2001) );
  XNOR2_X1 DP_mult_205_U1572 ( .A(DP_mult_205_n964), .B(DP_mult_205_n945), 
        .ZN(DP_mult_205_n2000) );
  XNOR2_X1 DP_mult_205_U1571 ( .A(DP_mult_205_n943), .B(DP_mult_205_n2000), 
        .ZN(DP_mult_205_n941) );
  INV_X2 DP_mult_205_U1570 ( .A(DP_mult_205_n2301), .ZN(DP_mult_205_n2299) );
  INV_X1 DP_mult_205_U1569 ( .A(DP_mult_205_n2325), .ZN(DP_mult_205_n2322) );
  XNOR2_X1 DP_mult_205_U1568 ( .A(DP_coeffs_fb_int[29]), .B(DP_mult_205_n2321), 
        .ZN(DP_mult_205_n1808) );
  INV_X2 DP_mult_205_U1567 ( .A(DP_mult_205_n2021), .ZN(DP_mult_205_n2175) );
  XNOR2_X1 DP_mult_205_U1566 ( .A(DP_mult_205_n1305), .B(DP_mult_205_n1437), 
        .ZN(DP_mult_205_n1999) );
  XNOR2_X1 DP_mult_205_U1565 ( .A(DP_mult_205_n1999), .B(DP_mult_205_n1937), 
        .ZN(DP_mult_205_n977) );
  INV_X2 DP_mult_205_U1564 ( .A(DP_mult_205_n2289), .ZN(DP_mult_205_n2288) );
  CLKBUF_X1 DP_mult_205_U1563 ( .A(DP_mult_205_n919), .Z(DP_mult_205_n1997) );
  INV_X1 DP_mult_205_U1562 ( .A(DP_mult_205_n2243), .ZN(DP_mult_205_n2242) );
  INV_X1 DP_mult_205_U1561 ( .A(DP_mult_205_n2268), .ZN(DP_mult_205_n1996) );
  INV_X1 DP_mult_205_U1560 ( .A(DP_mult_205_n2243), .ZN(DP_mult_205_n1995) );
  INV_X1 DP_mult_205_U1559 ( .A(DP_mult_205_n1986), .ZN(DP_mult_205_n2259) );
  XNOR2_X1 DP_mult_205_U1558 ( .A(DP_coeffs_fb_int[33]), .B(DP_mult_205_n2312), 
        .ZN(DP_mult_205_n1810) );
  INV_X1 DP_mult_205_U1557 ( .A(DP_mult_205_n2082), .ZN(DP_mult_205_n1994) );
  NOR2_X1 DP_mult_205_U1556 ( .A1(DP_mult_205_n1003), .A2(DP_mult_205_n1020), 
        .ZN(DP_mult_205_n1993) );
  XNOR2_X1 DP_mult_205_U1555 ( .A(DP_mult_205_n1974), .B(DP_mult_205_n2325), 
        .ZN(DP_mult_205_n2181) );
  XOR2_X1 DP_mult_205_U1554 ( .A(DP_coeffs_fb_int[31]), .B(
        DP_coeffs_fb_int[32]), .Z(DP_mult_205_n1992) );
  XNOR2_X1 DP_mult_205_U1553 ( .A(DP_coeffs_fb_int[37]), .B(DP_mult_205_n2305), 
        .ZN(DP_mult_205_n1812) );
  BUF_X1 DP_mult_205_U1552 ( .A(DP_mult_205_n2201), .Z(DP_mult_205_n1998) );
  INV_X1 DP_mult_205_U1551 ( .A(DP_mult_205_n2286), .ZN(DP_mult_205_n2284) );
  INV_X1 DP_mult_205_U1550 ( .A(DP_mult_205_n2286), .ZN(DP_mult_205_n2282) );
  CLKBUF_X1 DP_mult_205_U1549 ( .A(DP_mult_205_n1415), .Z(DP_mult_205_n1991)
         );
  INV_X2 DP_mult_205_U1548 ( .A(DP_mult_205_n2006), .ZN(DP_mult_205_n2271) );
  INV_X1 DP_mult_205_U1547 ( .A(DP_mult_205_n1982), .ZN(DP_mult_205_n1990) );
  AOI21_X1 DP_mult_205_U1546 ( .B1(DP_mult_205_n581), .B2(DP_mult_205_n567), 
        .A(DP_mult_205_n568), .ZN(DP_mult_205_n1989) );
  BUF_X2 DP_mult_205_U1545 ( .A(DP_mult_205_n279), .Z(DP_mult_205_n1988) );
  INV_X1 DP_mult_205_U1544 ( .A(DP_mult_205_n2021), .ZN(DP_mult_205_n2244) );
  INV_X1 DP_mult_205_U1543 ( .A(DP_mult_205_n2252), .ZN(DP_mult_205_n2251) );
  INV_X1 DP_mult_205_U1542 ( .A(DP_mult_205_n2252), .ZN(DP_mult_205_n1987) );
  INV_X1 DP_mult_205_U1541 ( .A(DP_coeffs_fb_int[34]), .ZN(DP_mult_205_n2309)
         );
  XOR2_X1 DP_mult_205_U1540 ( .A(DP_coeffs_fb_int[29]), .B(
        DP_coeffs_fb_int[30]), .Z(DP_mult_205_n2203) );
  XOR2_X1 DP_mult_205_U1539 ( .A(DP_coeffs_fb_int[29]), .B(
        DP_coeffs_fb_int[30]), .Z(DP_mult_205_n1986) );
  INV_X1 DP_mult_205_U1538 ( .A(DP_mult_205_n2103), .ZN(DP_mult_205_n1985) );
  INV_X2 DP_mult_205_U1537 ( .A(DP_mult_205_n2321), .ZN(DP_mult_205_n2318) );
  INV_X2 DP_mult_205_U1536 ( .A(DP_mult_205_n2321), .ZN(DP_mult_205_n2320) );
  XOR2_X1 DP_mult_205_U1535 ( .A(DP_coeffs_fb_int[25]), .B(DP_mult_205_n2328), 
        .Z(DP_mult_205_n1984) );
  XNOR2_X1 DP_mult_205_U1534 ( .A(DP_coeffs_fb_int[41]), .B(
        DP_coeffs_fb_int[42]), .ZN(DP_mult_205_n2030) );
  BUF_X2 DP_mult_205_U1533 ( .A(DP_mult_205_n2030), .Z(DP_mult_205_n1983) );
  BUF_X4 DP_mult_205_U1532 ( .A(DP_mult_205_n2030), .Z(DP_mult_205_n1982) );
  INV_X1 DP_mult_205_U1531 ( .A(DP_mult_205_n1961), .ZN(DP_mult_205_n2268) );
  INV_X1 DP_mult_205_U1530 ( .A(DP_coeffs_fb_int[34]), .ZN(DP_mult_205_n1979)
         );
  INV_X1 DP_mult_205_U1529 ( .A(DP_coeffs_fb_int[33]), .ZN(DP_mult_205_n1978)
         );
  NAND2_X1 DP_mult_205_U1528 ( .A1(DP_mult_205_n1980), .A2(DP_mult_205_n1981), 
        .ZN(DP_mult_205_n2205) );
  NAND2_X1 DP_mult_205_U1527 ( .A1(DP_mult_205_n1978), .A2(
        DP_coeffs_fb_int[34]), .ZN(DP_mult_205_n1981) );
  NAND2_X1 DP_mult_205_U1526 ( .A1(DP_coeffs_fb_int[33]), .A2(
        DP_mult_205_n1979), .ZN(DP_mult_205_n1980) );
  INV_X2 DP_mult_205_U1525 ( .A(DP_mult_205_n2250), .ZN(DP_mult_205_n2249) );
  BUF_X1 DP_mult_205_U1524 ( .A(DP_mult_205_n836), .Z(DP_mult_205_n2165) );
  INV_X1 DP_mult_205_U1523 ( .A(DP_mult_205_n2165), .ZN(DP_mult_205_n1977) );
  CLKBUF_X1 DP_mult_205_U1522 ( .A(DP_mult_205_n1393), .Z(DP_mult_205_n1976)
         );
  XNOR2_X1 DP_mult_205_U1521 ( .A(DP_coeffs_fb_int[47]), .B(DP_mult_205_n2286), 
        .ZN(DP_mult_205_n1817) );
  BUF_X1 DP_mult_205_U1520 ( .A(DP_mult_205_n514), .Z(DP_mult_205_n1975) );
  CLKBUF_X1 DP_mult_205_U1519 ( .A(DP_coeffs_fb_int[27]), .Z(DP_mult_205_n1974) );
  INV_X1 DP_mult_205_U1518 ( .A(DP_mult_205_n1998), .ZN(DP_mult_205_n2278) );
  INV_X1 DP_mult_205_U1517 ( .A(DP_mult_205_n1998), .ZN(DP_mult_205_n1973) );
  AND2_X1 DP_mult_205_U1516 ( .A1(DP_mult_205_n1812), .A2(DP_mult_205_n2269), 
        .ZN(DP_mult_205_n2022) );
  AND2_X2 DP_mult_205_U1515 ( .A1(DP_mult_205_n1810), .A2(DP_mult_205_n2264), 
        .ZN(DP_mult_205_n1972) );
  AND2_X1 DP_mult_205_U1514 ( .A1(DP_mult_205_n2181), .A2(DP_mult_205_n2008), 
        .ZN(DP_mult_205_n2207) );
  AND2_X1 DP_mult_205_U1513 ( .A1(DP_mult_205_n2181), .A2(DP_mult_205_n2008), 
        .ZN(DP_mult_205_n1971) );
  CLKBUF_X1 DP_mult_205_U1512 ( .A(DP_mult_205_n1076), .Z(DP_mult_205_n1970)
         );
  INV_X1 DP_mult_205_U1511 ( .A(DP_mult_205_n2022), .ZN(DP_mult_205_n1968) );
  INV_X1 DP_mult_205_U1510 ( .A(DP_mult_205_n2022), .ZN(DP_mult_205_n1969) );
  XNOR2_X1 DP_mult_205_U1509 ( .A(DP_coeffs_fb_int[41]), .B(DP_mult_205_n2297), 
        .ZN(DP_mult_205_n1814) );
  AND2_X1 DP_mult_205_U1508 ( .A1(DP_mult_205_n2217), .A2(DP_mult_205_n535), 
        .ZN(DP_mult_205_n1967) );
  XNOR2_X1 DP_mult_205_U1507 ( .A(DP_mult_205_n536), .B(DP_mult_205_n1967), 
        .ZN(DP_sw1_coeff_ret1[3]) );
  NOR2_X1 DP_mult_205_U1506 ( .A1(DP_mult_205_n963), .A2(DP_mult_205_n982), 
        .ZN(DP_mult_205_n558) );
  INV_X2 DP_mult_205_U1505 ( .A(DP_mult_205_n2309), .ZN(DP_mult_205_n2306) );
  NAND3_X1 DP_mult_205_U1504 ( .A1(DP_mult_205_n2150), .A2(DP_mult_205_n2151), 
        .A3(DP_mult_205_n2152), .ZN(DP_mult_205_n1966) );
  INV_X1 DP_mult_205_U1503 ( .A(DP_mult_205_n2306), .ZN(DP_mult_205_n1965) );
  AND2_X1 DP_mult_205_U1502 ( .A1(DP_mult_205_n2148), .A2(DP_mult_205_n2045), 
        .ZN(DP_mult_205_n1964) );
  XNOR2_X1 DP_mult_205_U1501 ( .A(DP_mult_205_n551), .B(DP_mult_205_n1964), 
        .ZN(DP_sw1_coeff_ret1[1]) );
  AND2_X1 DP_mult_205_U1500 ( .A1(DP_mult_205_n2226), .A2(DP_mult_205_n543), 
        .ZN(DP_mult_205_n1963) );
  XNOR2_X1 DP_mult_205_U1499 ( .A(DP_mult_205_n544), .B(DP_mult_205_n1963), 
        .ZN(DP_sw1_coeff_ret1[2]) );
  AND2_X1 DP_mult_205_U1498 ( .A1(DP_mult_205_n675), .A2(DP_mult_205_n559), 
        .ZN(DP_mult_205_n1962) );
  XNOR2_X1 DP_mult_205_U1497 ( .A(DP_mult_205_n560), .B(DP_mult_205_n1962), 
        .ZN(DP_sw1_coeff_ret1[0]) );
  XOR2_X1 DP_mult_205_U1496 ( .A(DP_coeffs_fb_int[35]), .B(
        DP_coeffs_fb_int[36]), .Z(DP_mult_205_n1961) );
  XOR2_X1 DP_mult_205_U1495 ( .A(DP_coeffs_fb_int[35]), .B(
        DP_coeffs_fb_int[36]), .Z(DP_mult_205_n1960) );
  OR2_X1 DP_mult_205_U1494 ( .A1(DP_mult_205_n1194), .A2(DP_mult_205_n676), 
        .ZN(DP_mult_205_n1959) );
  OR2_X1 DP_mult_205_U1493 ( .A1(DP_mult_205_n1143), .A2(DP_mult_205_n1150), 
        .ZN(DP_mult_205_n1958) );
  OR2_X1 DP_mult_205_U1492 ( .A1(DP_mult_205_n1151), .A2(DP_mult_205_n1158), 
        .ZN(DP_mult_205_n1957) );
  AND2_X1 DP_mult_205_U1491 ( .A1(DP_mult_205_n1021), .A2(DP_mult_205_n1038), 
        .ZN(DP_mult_205_n1956) );
  AND2_X1 DP_mult_205_U1490 ( .A1(DP_mult_205_n1133), .A2(DP_mult_205_n1142), 
        .ZN(DP_mult_205_n1955) );
  AND2_X1 DP_mult_205_U1489 ( .A1(DP_mult_205_n1055), .A2(DP_mult_205_n1070), 
        .ZN(DP_mult_205_n1954) );
  AND2_X1 DP_mult_205_U1488 ( .A1(DP_mult_205_n1123), .A2(DP_mult_205_n1132), 
        .ZN(DP_mult_205_n1953) );
  AND2_X1 DP_mult_205_U1487 ( .A1(DP_mult_205_n1179), .A2(DP_mult_205_n1433), 
        .ZN(DP_mult_205_n1952) );
  AND2_X1 DP_mult_205_U1486 ( .A1(DP_mult_205_n1457), .A2(DP_mult_205_n1480), 
        .ZN(DP_mult_205_n1951) );
  AND2_X1 DP_mult_205_U1485 ( .A1(DP_mult_205_n1238), .A2(DP_mult_205_n1216), 
        .ZN(DP_mult_205_n1950) );
  NAND2_X1 DP_mult_205_U1484 ( .A1(DP_mult_205_n1817), .A2(DP_mult_205_n2280), 
        .ZN(DP_mult_205_n1949) );
  INV_X1 DP_mult_205_U1483 ( .A(DP_coeffs_fb_int[32]), .ZN(DP_mult_205_n2312)
         );
  AND2_X1 DP_mult_205_U1482 ( .A1(DP_mult_205_n1151), .A2(DP_mult_205_n1158), 
        .ZN(DP_mult_205_n1948) );
  AND2_X1 DP_mult_205_U1481 ( .A1(DP_mult_205_n1143), .A2(DP_mult_205_n1150), 
        .ZN(DP_mult_205_n1947) );
  AND2_X1 DP_mult_205_U1480 ( .A1(DP_mult_205_n1039), .A2(DP_mult_205_n1054), 
        .ZN(DP_mult_205_n1946) );
  OR2_X1 DP_mult_205_U1479 ( .A1(DP_mult_205_n1179), .A2(DP_mult_205_n1433), 
        .ZN(DP_mult_205_n1945) );
  AND2_X1 DP_mult_205_U1478 ( .A1(DP_mult_205_n1111), .A2(DP_mult_205_n1122), 
        .ZN(DP_mult_205_n1944) );
  OR2_X1 DP_mult_205_U1477 ( .A1(DP_mult_205_n1457), .A2(DP_mult_205_n1480), 
        .ZN(DP_mult_205_n1943) );
  AND2_X1 DP_mult_205_U1476 ( .A1(DP_mult_205_n1193), .A2(DP_mult_205_n1481), 
        .ZN(DP_mult_205_n1942) );
  OR2_X1 DP_mult_205_U1475 ( .A1(DP_mult_205_n1055), .A2(DP_mult_205_n1070), 
        .ZN(DP_mult_205_n2221) );
  INV_X1 DP_mult_205_U1474 ( .A(DP_mult_205_n2049), .ZN(DP_mult_205_n2177) );
  AND2_X1 DP_mult_205_U1473 ( .A1(DP_mult_205_n1809), .A2(DP_mult_205_n2261), 
        .ZN(DP_mult_205_n2102) );
  INV_X1 DP_mult_205_U1472 ( .A(DP_coeffs_fb_int[30]), .ZN(DP_mult_205_n2317)
         );
  AOI21_X1 DP_mult_205_U1471 ( .B1(DP_mult_205_n526), .B2(DP_mult_205_n511), 
        .A(DP_mult_205_n512), .ZN(DP_mult_205_n1941) );
  AOI21_X2 DP_mult_205_U1470 ( .B1(DP_mult_205_n426), .B2(DP_mult_205_n445), 
        .A(DP_mult_205_n427), .ZN(DP_mult_205_n421) );
  NOR2_X1 DP_mult_205_U1469 ( .A1(DP_mult_205_n1984), .A2(DP_mult_205_n2206), 
        .ZN(DP_mult_205_n2049) );
  NOR2_X1 DP_mult_205_U1468 ( .A1(DP_mult_205_n1984), .A2(DP_mult_205_n2206), 
        .ZN(DP_mult_205_n1940) );
  INV_X1 DP_mult_205_U1467 ( .A(DP_coeffs_fb_int[24]), .ZN(DP_mult_205_n1939)
         );
  BUF_X1 DP_mult_205_U1466 ( .A(DP_mult_205_n1330), .Z(DP_mult_205_n1938) );
  BUF_X1 DP_mult_205_U1465 ( .A(DP_mult_205_n1327), .Z(DP_mult_205_n1937) );
  NAND3_X1 DP_mult_205_U1464 ( .A1(DP_mult_205_n2123), .A2(DP_mult_205_n2124), 
        .A3(DP_mult_205_n2125), .ZN(DP_mult_205_n1936) );
  INV_X1 DP_mult_205_U1463 ( .A(DP_mult_205_n2325), .ZN(DP_mult_205_n2323) );
  NAND3_X1 DP_mult_205_U1462 ( .A1(DP_mult_205_n2061), .A2(DP_mult_205_n2062), 
        .A3(DP_mult_205_n2063), .ZN(DP_mult_205_n1935) );
  XOR2_X1 DP_mult_205_U1461 ( .A(DP_coeffs_fb_int[25]), .B(
        DP_coeffs_fb_int[26]), .Z(DP_mult_205_n2206) );
  BUF_X1 DP_mult_205_U1460 ( .A(DP_mult_205_n2200), .Z(DP_mult_205_n2006) );
  INV_X2 DP_mult_205_U1459 ( .A(DP_mult_205_n2305), .ZN(DP_mult_205_n2304) );
  INV_X1 DP_mult_205_U1458 ( .A(DP_mult_205_n2275), .ZN(DP_mult_205_n2274) );
  INV_X1 DP_mult_205_U1457 ( .A(DP_mult_205_n2100), .ZN(DP_mult_205_n1934) );
  XNOR2_X1 DP_mult_205_U1456 ( .A(DP_coeffs_fb_int[39]), .B(DP_mult_205_n2301), 
        .ZN(DP_mult_205_n1813) );
  AND2_X2 DP_mult_205_U1455 ( .A1(DP_mult_205_n1980), .A2(DP_mult_205_n1981), 
        .ZN(DP_mult_205_n1933) );
  INV_X1 DP_mult_205_U1454 ( .A(DP_mult_205_n555), .ZN(DP_mult_205_n1932) );
  NAND2_X2 DP_mult_205_U1453 ( .A1(DP_mult_205_n1810), .A2(DP_mult_205_n2264), 
        .ZN(DP_mult_205_n289) );
  INV_X2 DP_mult_205_U1452 ( .A(DP_mult_205_n2006), .ZN(DP_mult_205_n2270) );
  INV_X1 DP_mult_205_U1451 ( .A(DP_sw1_0_), .ZN(DP_mult_205_n2329) );
  INV_X1 DP_mult_205_U1450 ( .A(DP_sw1_0_), .ZN(DP_mult_205_n1930) );
  INV_X1 DP_mult_205_U1449 ( .A(DP_sw1_0_), .ZN(DP_mult_205_n1931) );
  XNOR2_X1 DP_mult_205_U1448 ( .A(DP_mult_205_n859), .B(DP_mult_205_n2117), 
        .ZN(DP_mult_205_n1929) );
  HA_X1 DP_mult_205_U798 ( .A(DP_mult_205_n1456), .B(DP_mult_205_n1479), .CO(
        DP_mult_205_n1180), .S(DP_mult_205_n1181) );
  FA_X1 DP_mult_205_U797 ( .A(DP_mult_205_n1455), .B(DP_mult_205_n1478), .CI(
        DP_mult_205_n1180), .CO(DP_mult_205_n1178), .S(DP_mult_205_n1179) );
  HA_X1 DP_mult_205_U796 ( .A(DP_mult_205_n1432), .B(DP_mult_205_n1477), .CO(
        DP_mult_205_n1176), .S(DP_mult_205_n1177) );
  FA_X1 DP_mult_205_U795 ( .A(DP_mult_205_n1191), .B(DP_mult_205_n1454), .CI(
        DP_mult_205_n1177), .CO(DP_mult_205_n1174), .S(DP_mult_205_n1175) );
  FA_X1 DP_mult_205_U794 ( .A(DP_mult_205_n1476), .B(DP_mult_205_n1453), .CI(
        DP_mult_205_n1431), .CO(DP_mult_205_n1172), .S(DP_mult_205_n1173) );
  FA_X1 DP_mult_205_U793 ( .A(DP_mult_205_n1409), .B(DP_mult_205_n1176), .CI(
        DP_mult_205_n1173), .CO(DP_mult_205_n1170), .S(DP_mult_205_n1171) );
  HA_X1 DP_mult_205_U792 ( .A(DP_mult_205_n1408), .B(DP_mult_205_n1430), .CO(
        DP_mult_205_n1168), .S(DP_mult_205_n1169) );
  FA_X1 DP_mult_205_U791 ( .A(DP_mult_205_n1452), .B(DP_mult_205_n1475), .CI(
        DP_mult_205_n1190), .CO(DP_mult_205_n1166), .S(DP_mult_205_n1167) );
  FA_X1 DP_mult_205_U790 ( .A(DP_mult_205_n1172), .B(DP_mult_205_n1169), .CI(
        DP_mult_205_n1167), .CO(DP_mult_205_n1164), .S(DP_mult_205_n1165) );
  FA_X1 DP_mult_205_U789 ( .A(DP_mult_205_n1451), .B(DP_mult_205_n1474), .CI(
        DP_mult_205_n1407), .CO(DP_mult_205_n1162), .S(DP_mult_205_n1163) );
  FA_X1 DP_mult_205_U788 ( .A(DP_mult_205_n1168), .B(DP_mult_205_n1429), .CI(
        DP_mult_205_n1166), .CO(DP_mult_205_n1160), .S(DP_mult_205_n1161) );
  FA_X1 DP_mult_205_U787 ( .A(DP_mult_205_n1163), .B(DP_mult_205_n1385), .CI(
        DP_mult_205_n1164), .CO(DP_mult_205_n1158), .S(DP_mult_205_n1159) );
  HA_X1 DP_mult_205_U786 ( .A(DP_mult_205_n1384), .B(DP_mult_205_n1406), .CO(
        DP_mult_205_n1156), .S(DP_mult_205_n1157) );
  FA_X1 DP_mult_205_U785 ( .A(DP_mult_205_n1450), .B(DP_mult_205_n1428), .CI(
        DP_mult_205_n1189), .CO(DP_mult_205_n1154), .S(DP_mult_205_n1155) );
  FA_X1 DP_mult_205_U784 ( .A(DP_mult_205_n1157), .B(DP_mult_205_n1473), .CI(
        DP_mult_205_n1162), .CO(DP_mult_205_n1152), .S(DP_mult_205_n1153) );
  FA_X1 DP_mult_205_U783 ( .A(DP_mult_205_n1160), .B(DP_mult_205_n1155), .CI(
        DP_mult_205_n1153), .CO(DP_mult_205_n1150), .S(DP_mult_205_n1151) );
  FA_X1 DP_mult_205_U782 ( .A(DP_mult_205_n1383), .B(DP_mult_205_n1472), .CI(
        DP_mult_205_n1405), .CO(DP_mult_205_n1148), .S(DP_mult_205_n1149) );
  FA_X1 DP_mult_205_U781 ( .A(DP_mult_205_n1427), .B(DP_mult_205_n1449), .CI(
        DP_mult_205_n1156), .CO(DP_mult_205_n1146), .S(DP_mult_205_n1147) );
  FA_X1 DP_mult_205_U780 ( .A(DP_mult_205_n1361), .B(DP_mult_205_n1154), .CI(
        DP_mult_205_n1149), .CO(DP_mult_205_n1144), .S(DP_mult_205_n1145) );
  FA_X1 DP_mult_205_U779 ( .A(DP_mult_205_n1152), .B(DP_mult_205_n1147), .CI(
        DP_mult_205_n1145), .CO(DP_mult_205_n1142), .S(DP_mult_205_n1143) );
  HA_X1 DP_mult_205_U778 ( .A(DP_mult_205_n1382), .B(DP_mult_205_n1360), .CO(
        DP_mult_205_n1140), .S(DP_mult_205_n1141) );
  FA_X1 DP_mult_205_U777 ( .A(DP_mult_205_n1471), .B(DP_mult_205_n1426), .CI(
        DP_mult_205_n1188), .CO(DP_mult_205_n1138), .S(DP_mult_205_n1139) );
  FA_X1 DP_mult_205_U776 ( .A(DP_mult_205_n1404), .B(DP_mult_205_n1448), .CI(
        DP_mult_205_n1141), .CO(DP_mult_205_n1136), .S(DP_mult_205_n1137) );
  FA_X1 DP_mult_205_U775 ( .A(DP_mult_205_n1146), .B(DP_mult_205_n1148), .CI(
        DP_mult_205_n1139), .CO(DP_mult_205_n1134), .S(DP_mult_205_n1135) );
  FA_X1 DP_mult_205_U774 ( .A(DP_mult_205_n1144), .B(DP_mult_205_n1137), .CI(
        DP_mult_205_n1135), .CO(DP_mult_205_n1132), .S(DP_mult_205_n1133) );
  FA_X1 DP_mult_205_U773 ( .A(DP_mult_205_n1359), .B(DP_mult_205_n1470), .CI(
        DP_mult_205_n1381), .CO(DP_mult_205_n1130), .S(DP_mult_205_n1131) );
  FA_X1 DP_mult_205_U772 ( .A(DP_mult_205_n1403), .B(DP_mult_205_n1447), .CI(
        DP_mult_205_n1425), .CO(DP_mult_205_n1128), .S(DP_mult_205_n1129) );
  FA_X1 DP_mult_205_U771 ( .A(DP_mult_205_n1138), .B(DP_mult_205_n1140), .CI(
        DP_mult_205_n1337), .CO(DP_mult_205_n1126), .S(DP_mult_205_n1127) );
  FA_X1 DP_mult_205_U770 ( .A(DP_mult_205_n1131), .B(DP_mult_205_n1129), .CI(
        DP_mult_205_n1136), .CO(DP_mult_205_n1124), .S(DP_mult_205_n1125) );
  FA_X1 DP_mult_205_U769 ( .A(DP_mult_205_n1127), .B(DP_mult_205_n1134), .CI(
        DP_mult_205_n1125), .CO(DP_mult_205_n1122), .S(DP_mult_205_n1123) );
  HA_X1 DP_mult_205_U768 ( .A(DP_mult_205_n1336), .B(DP_mult_205_n1358), .CO(
        DP_mult_205_n1120), .S(DP_mult_205_n1121) );
  FA_X1 DP_mult_205_U767 ( .A(DP_mult_205_n1380), .B(DP_mult_205_n1402), .CI(
        DP_mult_205_n1187), .CO(DP_mult_205_n1118), .S(DP_mult_205_n1119) );
  FA_X1 DP_mult_205_U766 ( .A(DP_mult_205_n1424), .B(DP_mult_205_n1469), .CI(
        DP_mult_205_n1446), .CO(DP_mult_205_n1116), .S(DP_mult_205_n1117) );
  FA_X1 DP_mult_205_U765 ( .A(DP_mult_205_n1130), .B(DP_mult_205_n1121), .CI(
        DP_mult_205_n1128), .CO(DP_mult_205_n1114), .S(DP_mult_205_n1115) );
  FA_X1 DP_mult_205_U764 ( .A(DP_mult_205_n1119), .B(DP_mult_205_n1117), .CI(
        DP_mult_205_n1126), .CO(DP_mult_205_n1112), .S(DP_mult_205_n1113) );
  FA_X1 DP_mult_205_U762 ( .A(DP_mult_205_n1335), .B(DP_mult_205_n1468), .CI(
        DP_mult_205_n1357), .CO(DP_mult_205_n1108), .S(DP_mult_205_n1109) );
  FA_X1 DP_mult_205_U761 ( .A(DP_mult_205_n1401), .B(DP_mult_205_n1445), .CI(
        DP_mult_205_n1379), .CO(DP_mult_205_n1106), .S(DP_mult_205_n1107) );
  FA_X1 DP_mult_205_U760 ( .A(DP_mult_205_n1120), .B(DP_mult_205_n1423), .CI(
        DP_mult_205_n1118), .CO(DP_mult_205_n1104), .S(DP_mult_205_n1105) );
  FA_X1 DP_mult_205_U759 ( .A(DP_mult_205_n1313), .B(DP_mult_205_n1116), .CI(
        DP_mult_205_n1107), .CO(DP_mult_205_n1102), .S(DP_mult_205_n1103) );
  FA_X1 DP_mult_205_U758 ( .A(DP_mult_205_n1114), .B(DP_mult_205_n1109), .CI(
        DP_mult_205_n1105), .CO(DP_mult_205_n1100), .S(DP_mult_205_n1101) );
  FA_X1 DP_mult_205_U757 ( .A(DP_mult_205_n1103), .B(DP_mult_205_n1112), .CI(
        DP_mult_205_n1101), .CO(DP_mult_205_n1098), .S(DP_mult_205_n1099) );
  HA_X1 DP_mult_205_U756 ( .A(DP_mult_205_n1334), .B(DP_mult_205_n1312), .CO(
        DP_mult_205_n1096), .S(DP_mult_205_n1097) );
  FA_X1 DP_mult_205_U755 ( .A(DP_mult_205_n1467), .B(DP_mult_205_n1186), .CI(
        DP_mult_205_n1400), .CO(DP_mult_205_n1094), .S(DP_mult_205_n1095) );
  FA_X1 DP_mult_205_U754 ( .A(DP_mult_205_n1444), .B(DP_mult_205_n1356), .CI(
        DP_mult_205_n1378), .CO(DP_mult_205_n1092), .S(DP_mult_205_n1093) );
  FA_X1 DP_mult_205_U753 ( .A(DP_mult_205_n1097), .B(DP_mult_205_n1422), .CI(
        DP_mult_205_n1108), .CO(DP_mult_205_n1090), .S(DP_mult_205_n1091) );
  FA_X1 DP_mult_205_U752 ( .A(DP_mult_205_n1093), .B(DP_mult_205_n1106), .CI(
        DP_mult_205_n1095), .CO(DP_mult_205_n1088), .S(DP_mult_205_n1089) );
  FA_X1 DP_mult_205_U751 ( .A(DP_mult_205_n1102), .B(DP_mult_205_n1104), .CI(
        DP_mult_205_n1091), .CO(DP_mult_205_n1086), .S(DP_mult_205_n1087) );
  FA_X1 DP_mult_205_U750 ( .A(DP_mult_205_n1100), .B(DP_mult_205_n1089), .CI(
        DP_mult_205_n1087), .CO(DP_mult_205_n1084), .S(DP_mult_205_n1085) );
  FA_X1 DP_mult_205_U749 ( .A(DP_mult_205_n1311), .B(DP_mult_205_n1466), .CI(
        DP_mult_205_n1333), .CO(DP_mult_205_n1082), .S(DP_mult_205_n1083) );
  FA_X1 DP_mult_205_U748 ( .A(DP_mult_205_n1355), .B(DP_mult_205_n1443), .CI(
        DP_mult_205_n1377), .CO(DP_mult_205_n1080), .S(DP_mult_205_n1081) );
  FA_X1 DP_mult_205_U747 ( .A(DP_mult_205_n1399), .B(DP_mult_205_n1421), .CI(
        DP_mult_205_n1096), .CO(DP_mult_205_n1078), .S(DP_mult_205_n1079) );
  FA_X1 DP_mult_205_U746 ( .A(DP_mult_205_n1092), .B(DP_mult_205_n1289), .CI(
        DP_mult_205_n1094), .CO(DP_mult_205_n1076), .S(DP_mult_205_n1077) );
  FA_X1 DP_mult_205_U745 ( .A(DP_mult_205_n1083), .B(DP_mult_205_n1081), .CI(
        DP_mult_205_n1079), .CO(DP_mult_205_n1074), .S(DP_mult_205_n1075) );
  FA_X1 DP_mult_205_U744 ( .A(DP_mult_205_n1088), .B(DP_mult_205_n1090), .CI(
        DP_mult_205_n1077), .CO(DP_mult_205_n1072), .S(DP_mult_205_n1073) );
  FA_X1 DP_mult_205_U743 ( .A(DP_mult_205_n1086), .B(DP_mult_205_n1075), .CI(
        DP_mult_205_n1073), .CO(DP_mult_205_n1070), .S(DP_mult_205_n1071) );
  HA_X1 DP_mult_205_U742 ( .A(DP_mult_205_n1288), .B(DP_mult_205_n1310), .CO(
        DP_mult_205_n1068), .S(DP_mult_205_n1069) );
  FA_X1 DP_mult_205_U741 ( .A(DP_mult_205_n1185), .B(DP_mult_205_n1376), .CI(
        DP_mult_205_n1465), .CO(DP_mult_205_n1066), .S(DP_mult_205_n1067) );
  FA_X1 DP_mult_205_U740 ( .A(DP_mult_205_n1332), .B(DP_mult_205_n1354), .CI(
        DP_mult_205_n1442), .CO(DP_mult_205_n1064), .S(DP_mult_205_n1065) );
  FA_X1 DP_mult_205_U739 ( .A(DP_mult_205_n1398), .B(DP_mult_205_n1420), .CI(
        DP_mult_205_n1069), .CO(DP_mult_205_n1062), .S(DP_mult_205_n1063) );
  FA_X1 DP_mult_205_U738 ( .A(DP_mult_205_n1080), .B(DP_mult_205_n1082), .CI(
        DP_mult_205_n1078), .CO(DP_mult_205_n1060), .S(DP_mult_205_n1061) );
  FA_X1 DP_mult_205_U736 ( .A(DP_mult_205_n1061), .B(DP_mult_205_n1063), .CI(
        DP_mult_205_n1074), .CO(DP_mult_205_n1056), .S(DP_mult_205_n1057) );
  FA_X1 DP_mult_205_U735 ( .A(DP_mult_205_n1072), .B(DP_mult_205_n1059), .CI(
        DP_mult_205_n1057), .CO(DP_mult_205_n1054), .S(DP_mult_205_n1055) );
  FA_X1 DP_mult_205_U734 ( .A(DP_mult_205_n1287), .B(DP_mult_205_n1464), .CI(
        DP_mult_205_n1309), .CO(DP_mult_205_n1052), .S(DP_mult_205_n1053) );
  FA_X1 DP_mult_205_U733 ( .A(DP_mult_205_n1331), .B(DP_mult_205_n1353), .CI(
        DP_mult_205_n1375), .CO(DP_mult_205_n1050), .S(DP_mult_205_n1051) );
  FA_X1 DP_mult_205_U732 ( .A(DP_mult_205_n1397), .B(DP_mult_205_n1441), .CI(
        DP_mult_205_n1419), .CO(DP_mult_205_n1048), .S(DP_mult_205_n1049) );
  FA_X1 DP_mult_205_U731 ( .A(DP_mult_205_n1064), .B(DP_mult_205_n1068), .CI(
        DP_mult_205_n1066), .CO(DP_mult_205_n1046), .S(DP_mult_205_n1047) );
  FA_X1 DP_mult_205_U730 ( .A(DP_mult_205_n1049), .B(DP_mult_205_n1265), .CI(
        DP_mult_205_n1051), .CO(DP_mult_205_n1044), .S(DP_mult_205_n1045) );
  FA_X1 DP_mult_205_U728 ( .A(DP_mult_205_n1058), .B(DP_mult_205_n1047), .CI(
        DP_mult_205_n1045), .CO(DP_mult_205_n1040), .S(DP_mult_205_n1041) );
  FA_X1 DP_mult_205_U727 ( .A(DP_mult_205_n1056), .B(DP_mult_205_n1043), .CI(
        DP_mult_205_n1041), .CO(DP_mult_205_n1038), .S(DP_mult_205_n1039) );
  HA_X1 DP_mult_205_U726 ( .A(DP_mult_205_n1286), .B(DP_mult_205_n1264), .CO(
        DP_mult_205_n1036), .S(DP_mult_205_n1037) );
  FA_X1 DP_mult_205_U725 ( .A(DP_mult_205_n1308), .B(DP_mult_205_n1184), .CI(
        DP_mult_205_n1374), .CO(DP_mult_205_n1034), .S(DP_mult_205_n1035) );
  FA_X1 DP_mult_205_U723 ( .A(DP_mult_205_n1418), .B(DP_mult_205_n1440), .CI(
        DP_mult_205_n1352), .CO(DP_mult_205_n1030), .S(DP_mult_205_n1031) );
  FA_X1 DP_mult_205_U722 ( .A(DP_mult_205_n1052), .B(DP_mult_205_n1037), .CI(
        DP_mult_205_n1050), .CO(DP_mult_205_n1028), .S(DP_mult_205_n1029) );
  FA_X1 DP_mult_205_U721 ( .A(DP_mult_205_n1031), .B(DP_mult_205_n1048), .CI(
        DP_mult_205_n1033), .CO(DP_mult_205_n1026), .S(DP_mult_205_n1027) );
  FA_X1 DP_mult_205_U720 ( .A(DP_mult_205_n1046), .B(DP_mult_205_n1035), .CI(
        DP_mult_205_n1029), .CO(DP_mult_205_n1024), .S(DP_mult_205_n1025) );
  FA_X1 DP_mult_205_U718 ( .A(DP_mult_205_n1040), .B(DP_mult_205_n1025), .CI(
        DP_mult_205_n1023), .CO(DP_mult_205_n1020), .S(DP_mult_205_n1021) );
  FA_X1 DP_mult_205_U716 ( .A(DP_mult_205_n1307), .B(DP_mult_205_n1329), .CI(
        DP_mult_205_n1373), .CO(DP_mult_205_n1016), .S(DP_mult_205_n1017) );
  FA_X1 DP_mult_205_U715 ( .A(DP_mult_205_n1417), .B(DP_mult_205_n1462), .CI(
        DP_mult_205_n1395), .CO(DP_mult_205_n1014), .S(DP_mult_205_n1015) );
  FA_X1 DP_mult_205_U713 ( .A(DP_mult_205_n1030), .B(DP_mult_205_n1034), .CI(
        DP_mult_205_n1241), .CO(DP_mult_205_n1010), .S(DP_mult_205_n1011) );
  FA_X1 DP_mult_205_U712 ( .A(DP_mult_205_n1019), .B(DP_mult_205_n1015), .CI(
        DP_mult_205_n1017), .CO(DP_mult_205_n1008), .S(DP_mult_205_n1009) );
  FA_X1 DP_mult_205_U711 ( .A(DP_mult_205_n1013), .B(DP_mult_205_n1028), .CI(
        DP_mult_205_n1026), .CO(DP_mult_205_n1006), .S(DP_mult_205_n1007) );
  FA_X1 DP_mult_205_U710 ( .A(DP_mult_205_n1009), .B(DP_mult_205_n1011), .CI(
        DP_mult_205_n1024), .CO(DP_mult_205_n1004), .S(DP_mult_205_n1005) );
  FA_X1 DP_mult_205_U709 ( .A(DP_mult_205_n1022), .B(DP_mult_205_n1007), .CI(
        DP_mult_205_n1005), .CO(DP_mult_205_n1002), .S(DP_mult_205_n1003) );
  HA_X1 DP_mult_205_U708 ( .A(DP_mult_205_n1240), .B(DP_mult_205_n1262), .CO(
        DP_mult_205_n1000), .S(DP_mult_205_n1001) );
  FA_X1 DP_mult_205_U707 ( .A(DP_mult_205_n1461), .B(DP_mult_205_n1350), .CI(
        DP_mult_205_n1183), .CO(DP_mult_205_n998), .S(DP_mult_205_n999) );
  FA_X1 DP_mult_205_U706 ( .A(DP_mult_205_n1438), .B(DP_mult_205_n1284), .CI(
        DP_mult_205_n1372), .CO(DP_mult_205_n996), .S(DP_mult_205_n997) );
  FA_X1 DP_mult_205_U705 ( .A(DP_mult_205_n1328), .B(DP_mult_205_n1416), .CI(
        DP_mult_205_n1306), .CO(DP_mult_205_n994), .S(DP_mult_205_n995) );
  FA_X1 DP_mult_205_U703 ( .A(DP_mult_205_n1014), .B(DP_mult_205_n1016), .CI(
        DP_mult_205_n995), .CO(DP_mult_205_n990), .S(DP_mult_205_n991) );
  FA_X1 DP_mult_205_U702 ( .A(DP_mult_205_n999), .B(DP_mult_205_n997), .CI(
        DP_mult_205_n1012), .CO(DP_mult_205_n988), .S(DP_mult_205_n989) );
  FA_X1 DP_mult_205_U701 ( .A(DP_mult_205_n993), .B(DP_mult_205_n1010), .CI(
        DP_mult_205_n1008), .CO(DP_mult_205_n986), .S(DP_mult_205_n987) );
  FA_X1 DP_mult_205_U700 ( .A(DP_mult_205_n989), .B(DP_mult_205_n991), .CI(
        DP_mult_205_n1006), .CO(DP_mult_205_n984), .S(DP_mult_205_n985) );
  FA_X1 DP_mult_205_U699 ( .A(DP_mult_205_n1004), .B(DP_mult_205_n987), .CI(
        DP_mult_205_n985), .CO(DP_mult_205_n982), .S(DP_mult_205_n983) );
  FA_X1 DP_mult_205_U698 ( .A(DP_mult_205_n1239), .B(DP_mult_205_n1261), .CI(
        DP_mult_205_n1349), .CO(DP_mult_205_n980), .S(DP_mult_205_n981) );
  FA_X1 DP_mult_205_U697 ( .A(DP_mult_205_n1460), .B(DP_mult_205_n1283), .CI(
        DP_mult_205_n1371), .CO(DP_mult_205_n978), .S(DP_mult_205_n979) );
  FA_X1 DP_mult_205_U694 ( .A(DP_mult_205_n994), .B(DP_mult_205_n996), .CI(
        DP_mult_205_n1217), .CO(DP_mult_205_n972), .S(DP_mult_205_n973) );
  FA_X1 DP_mult_205_U692 ( .A(DP_mult_205_n975), .B(DP_mult_205_n981), .CI(
        DP_mult_205_n992), .CO(DP_mult_205_n968), .S(DP_mult_205_n969) );
  FA_X1 DP_mult_205_U691 ( .A(DP_mult_205_n973), .B(DP_mult_205_n990), .CI(
        DP_mult_205_n988), .CO(DP_mult_205_n966), .S(DP_mult_205_n967) );
  FA_X1 DP_mult_205_U690 ( .A(DP_mult_205_n969), .B(DP_mult_205_n971), .CI(
        DP_mult_205_n986), .CO(DP_mult_205_n964), .S(DP_mult_205_n965) );
  FA_X1 DP_mult_205_U684 ( .A(DP_mult_205_n1326), .B(DP_mult_205_n1392), .CI(
        DP_mult_205_n961), .CO(DP_mult_205_n952), .S(DP_mult_205_n953) );
  FA_X1 DP_mult_205_U683 ( .A(DP_mult_205_n980), .B(DP_mult_205_n976), .CI(
        DP_mult_205_n978), .CO(DP_mult_205_n950), .S(DP_mult_205_n951) );
  FA_X1 DP_mult_205_U682 ( .A(DP_mult_205_n955), .B(DP_mult_205_n974), .CI(
        DP_mult_205_n957), .CO(DP_mult_205_n948), .S(DP_mult_205_n949) );
  FA_X1 DP_mult_205_U681 ( .A(DP_mult_205_n972), .B(DP_mult_205_n959), .CI(
        DP_mult_205_n953), .CO(DP_mult_205_n946), .S(DP_mult_205_n947) );
  FA_X1 DP_mult_205_U680 ( .A(DP_mult_205_n951), .B(DP_mult_205_n970), .CI(
        DP_mult_205_n968), .CO(DP_mult_205_n944), .S(DP_mult_205_n945) );
  FA_X1 DP_mult_205_U679 ( .A(DP_mult_205_n947), .B(DP_mult_205_n949), .CI(
        DP_mult_205_n966), .CO(DP_mult_205_n942), .S(DP_mult_205_n943) );
  FA_X1 DP_mult_205_U675 ( .A(DP_mult_205_n1259), .B(DP_mult_205_n1347), .CI(
        DP_mult_205_n1303), .CO(DP_mult_205_n936), .S(DP_mult_205_n937) );
  FA_X1 DP_mult_205_U674 ( .A(DP_mult_205_n1281), .B(DP_mult_205_n1369), .CI(
        DP_mult_205_n1391), .CO(DP_mult_205_n934), .S(DP_mult_205_n935) );
  FA_X1 DP_mult_205_U673 ( .A(DP_mult_205_n1435), .B(DP_mult_205_n1413), .CI(
        DP_mult_205_n1325), .CO(DP_mult_205_n932), .S(DP_mult_205_n933) );
  FA_X1 DP_mult_205_U672 ( .A(DP_mult_205_n939), .B(DP_mult_205_n1950), .CI(
        DP_mult_205_n1458), .CO(DP_mult_205_n930), .S(DP_mult_205_n931) );
  FA_X1 DP_mult_205_U671 ( .A(DP_mult_205_n958), .B(DP_mult_205_n954), .CI(
        DP_mult_205_n956), .CO(DP_mult_205_n928), .S(DP_mult_205_n929) );
  FA_X1 DP_mult_205_U670 ( .A(DP_mult_205_n937), .B(DP_mult_205_n933), .CI(
        DP_mult_205_n952), .CO(DP_mult_205_n926), .S(DP_mult_205_n927) );
  FA_X1 DP_mult_205_U669 ( .A(DP_mult_205_n950), .B(DP_mult_205_n935), .CI(
        DP_mult_205_n931), .CO(DP_mult_205_n924), .S(DP_mult_205_n925) );
  FA_X1 DP_mult_205_U667 ( .A(DP_mult_205_n925), .B(DP_mult_205_n927), .CI(
        DP_mult_205_n944), .CO(DP_mult_205_n920), .S(DP_mult_205_n921) );
  FA_X1 DP_mult_205_U666 ( .A(DP_mult_205_n942), .B(DP_mult_205_n923), .CI(
        DP_mult_205_n921), .CO(DP_mult_205_n918), .S(DP_mult_205_n919) );
  FA_X1 DP_mult_205_U664 ( .A(DP_mult_205_n917), .B(DP_mult_205_n1302), .CI(
        DP_mult_205_n1214), .CO(DP_mult_205_n914), .S(DP_mult_205_n915) );
  FA_X1 DP_mult_205_U663 ( .A(DP_mult_205_n1412), .B(DP_mult_205_n1236), .CI(
        DP_mult_205_n1258), .CO(DP_mult_205_n912), .S(DP_mult_205_n913) );
  FA_X1 DP_mult_205_U662 ( .A(DP_mult_205_n1346), .B(DP_mult_205_n1280), .CI(
        DP_mult_205_n1324), .CO(DP_mult_205_n910), .S(DP_mult_205_n911) );
  FA_X1 DP_mult_205_U661 ( .A(DP_mult_205_n1368), .B(DP_mult_205_n1390), .CI(
        DP_mult_205_n938), .CO(DP_mult_205_n908), .S(DP_mult_205_n909) );
  FA_X1 DP_mult_205_U660 ( .A(DP_mult_205_n932), .B(DP_mult_205_n936), .CI(
        DP_mult_205_n934), .CO(DP_mult_205_n906), .S(DP_mult_205_n907) );
  FA_X1 DP_mult_205_U659 ( .A(DP_mult_205_n911), .B(DP_mult_205_n913), .CI(
        DP_mult_205_n915), .CO(DP_mult_205_n904), .S(DP_mult_205_n905) );
  FA_X1 DP_mult_205_U658 ( .A(DP_mult_205_n909), .B(DP_mult_205_n930), .CI(
        DP_mult_205_n928), .CO(DP_mult_205_n902), .S(DP_mult_205_n903) );
  FA_X1 DP_mult_205_U657 ( .A(DP_mult_205_n926), .B(DP_mult_205_n907), .CI(
        DP_mult_205_n905), .CO(DP_mult_205_n900), .S(DP_mult_205_n901) );
  FA_X1 DP_mult_205_U655 ( .A(DP_mult_205_n920), .B(DP_mult_205_n901), .CI(
        DP_mult_205_n899), .CO(DP_mult_205_n896), .S(DP_mult_205_n897) );
  FA_X1 DP_mult_205_U654 ( .A(DP_mult_205_n1411), .B(DP_mult_205_n1235), .CI(
        DP_mult_205_n1213), .CO(DP_mult_205_n894), .S(DP_mult_205_n895) );
  FA_X1 DP_mult_205_U653 ( .A(DP_mult_205_n1279), .B(DP_mult_205_n1323), .CI(
        DP_mult_205_n2017), .CO(DP_mult_205_n892), .S(DP_mult_205_n893) );
  FA_X1 DP_mult_205_U652 ( .A(DP_mult_205_n1257), .B(DP_mult_205_n1301), .CI(
        DP_mult_205_n1345), .CO(DP_mult_205_n890), .S(DP_mult_205_n891) );
  FA_X1 DP_mult_205_U651 ( .A(DP_mult_205_n1367), .B(DP_mult_205_n1389), .CI(
        DP_mult_205_n1434), .CO(DP_mult_205_n888), .S(DP_mult_205_n889) );
  FA_X1 DP_mult_205_U650 ( .A(DP_mult_205_n910), .B(DP_mult_205_n912), .CI(
        DP_mult_205_n914), .CO(DP_mult_205_n886), .S(DP_mult_205_n887) );
  FA_X1 DP_mult_205_U648 ( .A(DP_mult_205_n889), .B(DP_mult_205_n893), .CI(
        DP_mult_205_n906), .CO(DP_mult_205_n882), .S(DP_mult_205_n883) );
  FA_X1 DP_mult_205_U647 ( .A(DP_mult_205_n887), .B(DP_mult_205_n904), .CI(
        DP_mult_205_n902), .CO(DP_mult_205_n880), .S(DP_mult_205_n881) );
  FA_X1 DP_mult_205_U646 ( .A(DP_mult_205_n883), .B(DP_mult_205_n885), .CI(
        DP_mult_205_n900), .CO(DP_mult_205_n878), .S(DP_mult_205_n879) );
  FA_X1 DP_mult_205_U645 ( .A(DP_mult_205_n898), .B(DP_mult_205_n881), .CI(
        DP_mult_205_n879), .CO(DP_mult_205_n876), .S(DP_mult_205_n877) );
  FA_X1 DP_mult_205_U643 ( .A(DP_mult_205_n1388), .B(DP_mult_205_n1278), .CI(
        DP_mult_205_n875), .CO(DP_mult_205_n872), .S(DP_mult_205_n873) );
  FA_X1 DP_mult_205_U642 ( .A(DP_mult_205_n1212), .B(DP_mult_205_n1344), .CI(
        DP_mult_205_n1366), .CO(DP_mult_205_n870), .S(DP_mult_205_n871) );
  FA_X1 DP_mult_205_U641 ( .A(DP_mult_205_n1256), .B(DP_mult_205_n1322), .CI(
        DP_mult_205_n1234), .CO(DP_mult_205_n868), .S(DP_mult_205_n869) );
  FA_X1 DP_mult_205_U640 ( .A(DP_mult_205_n894), .B(DP_mult_205_n1300), .CI(
        DP_mult_205_n892), .CO(DP_mult_205_n866), .S(DP_mult_205_n867) );
  FA_X1 DP_mult_205_U639 ( .A(DP_mult_205_n890), .B(DP_mult_205_n869), .CI(
        DP_mult_205_n871), .CO(DP_mult_205_n864), .S(DP_mult_205_n865) );
  FA_X1 DP_mult_205_U638 ( .A(DP_mult_205_n888), .B(DP_mult_205_n873), .CI(
        DP_mult_205_n886), .CO(DP_mult_205_n862), .S(DP_mult_205_n863) );
  FA_X1 DP_mult_205_U637 ( .A(DP_mult_205_n884), .B(DP_mult_205_n867), .CI(
        DP_mult_205_n865), .CO(DP_mult_205_n860), .S(DP_mult_205_n861) );
  FA_X1 DP_mult_205_U636 ( .A(DP_mult_205_n863), .B(DP_mult_205_n882), .CI(
        DP_mult_205_n880), .CO(DP_mult_205_n858), .S(DP_mult_205_n859) );
  FA_X1 DP_mult_205_U634 ( .A(DP_mult_205_n1387), .B(DP_mult_205_n1233), .CI(
        DP_mult_205_n1211), .CO(DP_mult_205_n854), .S(DP_mult_205_n855) );
  FA_X1 DP_mult_205_U633 ( .A(DP_mult_205_n874), .B(DP_mult_205_n1321), .CI(
        DP_mult_205_n1255), .CO(DP_mult_205_n852), .S(DP_mult_205_n853) );
  FA_X1 DP_mult_205_U632 ( .A(DP_mult_205_n1343), .B(DP_mult_205_n1299), .CI(
        DP_mult_205_n1277), .CO(DP_mult_205_n850), .S(DP_mult_205_n851) );
  FA_X1 DP_mult_205_U631 ( .A(DP_mult_205_n1410), .B(DP_mult_205_n1365), .CI(
        DP_mult_205_n872), .CO(DP_mult_205_n848), .S(DP_mult_205_n849) );
  FA_X1 DP_mult_205_U629 ( .A(DP_mult_205_n855), .B(DP_mult_205_n853), .CI(
        DP_mult_205_n866), .CO(DP_mult_205_n844), .S(DP_mult_205_n845) );
  FA_X1 DP_mult_205_U628 ( .A(DP_mult_205_n864), .B(DP_mult_205_n849), .CI(
        DP_mult_205_n862), .CO(DP_mult_205_n842), .S(DP_mult_205_n843) );
  FA_X1 DP_mult_205_U627 ( .A(DP_mult_205_n845), .B(DP_mult_205_n847), .CI(
        DP_mult_205_n860), .CO(DP_mult_205_n840), .S(DP_mult_205_n841) );
  FA_X1 DP_mult_205_U626 ( .A(DP_mult_205_n858), .B(DP_mult_205_n843), .CI(
        DP_mult_205_n841), .CO(DP_mult_205_n838), .S(DP_mult_205_n839) );
  FA_X1 DP_mult_205_U623 ( .A(DP_mult_205_n1232), .B(DP_mult_205_n1364), .CI(
        DP_mult_205_n1342), .CO(DP_mult_205_n832), .S(DP_mult_205_n833) );
  FA_X1 DP_mult_205_U621 ( .A(DP_mult_205_n854), .B(DP_mult_205_n850), .CI(
        DP_mult_205_n852), .CO(DP_mult_205_n828), .S(DP_mult_205_n829) );
  FA_X1 DP_mult_205_U620 ( .A(DP_mult_205_n835), .B(DP_mult_205_n831), .CI(
        DP_mult_205_n833), .CO(DP_mult_205_n826), .S(DP_mult_205_n827) );
  FA_X1 DP_mult_205_U619 ( .A(DP_mult_205_n846), .B(DP_mult_205_n848), .CI(
        DP_mult_205_n829), .CO(DP_mult_205_n824), .S(DP_mult_205_n825) );
  FA_X1 DP_mult_205_U618 ( .A(DP_mult_205_n827), .B(DP_mult_205_n844), .CI(
        DP_mult_205_n842), .CO(DP_mult_205_n822), .S(DP_mult_205_n823) );
  FA_X1 DP_mult_205_U615 ( .A(DP_mult_205_n1231), .B(DP_mult_205_n1297), .CI(
        DP_mult_205_n1275), .CO(DP_mult_205_n816), .S(DP_mult_205_n817) );
  FA_X1 DP_mult_205_U614 ( .A(DP_mult_205_n1319), .B(DP_mult_205_n1253), .CI(
        DP_mult_205_n1341), .CO(DP_mult_205_n814), .S(DP_mult_205_n815) );
  FA_X1 DP_mult_205_U613 ( .A(DP_mult_205_n834), .B(DP_mult_205_n1386), .CI(
        DP_mult_205_n830), .CO(DP_mult_205_n812), .S(DP_mult_205_n813) );
  FA_X1 DP_mult_205_U612 ( .A(DP_mult_205_n815), .B(DP_mult_205_n832), .CI(
        DP_mult_205_n817), .CO(DP_mult_205_n810), .S(DP_mult_205_n811) );
  FA_X1 DP_mult_205_U611 ( .A(DP_mult_205_n828), .B(DP_mult_205_n819), .CI(
        DP_mult_205_n813), .CO(DP_mult_205_n808), .S(DP_mult_205_n809) );
  FA_X1 DP_mult_205_U607 ( .A(DP_mult_205_n1340), .B(DP_mult_205_n1252), .CI(
        DP_mult_205_n803), .CO(DP_mult_205_n800), .S(DP_mult_205_n801) );
  FA_X1 DP_mult_205_U606 ( .A(DP_mult_205_n1208), .B(DP_mult_205_n1318), .CI(
        DP_mult_205_n1230), .CO(DP_mult_205_n798), .S(DP_mult_205_n799) );
  FA_X1 DP_mult_205_U604 ( .A(DP_mult_205_n814), .B(DP_mult_205_n816), .CI(
        DP_mult_205_n799), .CO(DP_mult_205_n794), .S(DP_mult_205_n795) );
  FA_X1 DP_mult_205_U603 ( .A(DP_mult_205_n797), .B(DP_mult_205_n801), .CI(
        DP_mult_205_n812), .CO(DP_mult_205_n792), .S(DP_mult_205_n793) );
  FA_X1 DP_mult_205_U602 ( .A(DP_mult_205_n795), .B(DP_mult_205_n810), .CI(
        DP_mult_205_n808), .CO(DP_mult_205_n790), .S(DP_mult_205_n791) );
  FA_X1 DP_mult_205_U601 ( .A(DP_mult_205_n806), .B(DP_mult_205_n793), .CI(
        DP_mult_205_n791), .CO(DP_mult_205_n788), .S(DP_mult_205_n789) );
  FA_X1 DP_mult_205_U600 ( .A(DP_mult_205_n1251), .B(DP_mult_205_n1207), .CI(
        DP_mult_205_n802), .CO(DP_mult_205_n786), .S(DP_mult_205_n787) );
  FA_X1 DP_mult_205_U599 ( .A(DP_mult_205_n1273), .B(DP_mult_205_n1317), .CI(
        DP_mult_205_n1295), .CO(DP_mult_205_n784), .S(DP_mult_205_n785) );
  FA_X1 DP_mult_205_U598 ( .A(DP_mult_205_n1339), .B(DP_mult_205_n1229), .CI(
        DP_mult_205_n1362), .CO(DP_mult_205_n782), .S(DP_mult_205_n783) );
  FA_X1 DP_mult_205_U597 ( .A(DP_mult_205_n798), .B(DP_mult_205_n800), .CI(
        DP_mult_205_n785), .CO(DP_mult_205_n780), .S(DP_mult_205_n781) );
  FA_X1 DP_mult_205_U596 ( .A(DP_mult_205_n796), .B(DP_mult_205_n787), .CI(
        DP_mult_205_n783), .CO(DP_mult_205_n778), .S(DP_mult_205_n779) );
  FA_X1 DP_mult_205_U595 ( .A(DP_mult_205_n781), .B(DP_mult_205_n794), .CI(
        DP_mult_205_n792), .CO(DP_mult_205_n776), .S(DP_mult_205_n777) );
  FA_X1 DP_mult_205_U594 ( .A(DP_mult_205_n790), .B(DP_mult_205_n779), .CI(
        DP_mult_205_n777), .CO(DP_mult_205_n774), .S(DP_mult_205_n775) );
  FA_X1 DP_mult_205_U592 ( .A(DP_mult_205_n1316), .B(DP_mult_205_n1250), .CI(
        DP_mult_205_n773), .CO(DP_mult_205_n770), .S(DP_mult_205_n771) );
  FA_X1 DP_mult_205_U591 ( .A(DP_mult_205_n1294), .B(DP_mult_205_n1206), .CI(
        DP_mult_205_n1272), .CO(DP_mult_205_n768), .S(DP_mult_205_n769) );
  FA_X1 DP_mult_205_U590 ( .A(DP_mult_205_n786), .B(DP_mult_205_n1228), .CI(
        DP_mult_205_n784), .CO(DP_mult_205_n766), .S(DP_mult_205_n767) );
  FA_X1 DP_mult_205_U589 ( .A(DP_mult_205_n771), .B(DP_mult_205_n769), .CI(
        DP_mult_205_n782), .CO(DP_mult_205_n764), .S(DP_mult_205_n765) );
  FA_X1 DP_mult_205_U588 ( .A(DP_mult_205_n767), .B(DP_mult_205_n780), .CI(
        DP_mult_205_n778), .CO(DP_mult_205_n762), .S(DP_mult_205_n763) );
  FA_X1 DP_mult_205_U587 ( .A(DP_mult_205_n776), .B(DP_mult_205_n765), .CI(
        DP_mult_205_n763), .CO(DP_mult_205_n760), .S(DP_mult_205_n761) );
  FA_X1 DP_mult_205_U586 ( .A(DP_mult_205_n772), .B(DP_mult_205_n1205), .CI(
        DP_mult_205_n1227), .CO(DP_mult_205_n758), .S(DP_mult_205_n759) );
  FA_X1 DP_mult_205_U585 ( .A(DP_mult_205_n1315), .B(DP_mult_205_n1293), .CI(
        DP_mult_205_n1249), .CO(DP_mult_205_n756), .S(DP_mult_205_n757) );
  FA_X1 DP_mult_205_U584 ( .A(DP_mult_205_n1338), .B(DP_mult_205_n1271), .CI(
        DP_mult_205_n770), .CO(DP_mult_205_n754), .S(DP_mult_205_n755) );
  FA_X1 DP_mult_205_U583 ( .A(DP_mult_205_n757), .B(DP_mult_205_n768), .CI(
        DP_mult_205_n759), .CO(DP_mult_205_n752), .S(DP_mult_205_n753) );
  FA_X1 DP_mult_205_U582 ( .A(DP_mult_205_n755), .B(DP_mult_205_n766), .CI(
        DP_mult_205_n764), .CO(DP_mult_205_n750), .S(DP_mult_205_n751) );
  FA_X1 DP_mult_205_U581 ( .A(DP_mult_205_n762), .B(DP_mult_205_n753), .CI(
        DP_mult_205_n751), .CO(DP_mult_205_n748), .S(DP_mult_205_n749) );
  FA_X1 DP_mult_205_U579 ( .A(DP_mult_205_n1292), .B(DP_mult_205_n1248), .CI(
        DP_mult_205_n747), .CO(DP_mult_205_n744), .S(DP_mult_205_n745) );
  FA_X1 DP_mult_205_U578 ( .A(DP_mult_205_n1226), .B(DP_mult_205_n1204), .CI(
        DP_mult_205_n1270), .CO(DP_mult_205_n742), .S(DP_mult_205_n743) );
  FA_X1 DP_mult_205_U577 ( .A(DP_mult_205_n756), .B(DP_mult_205_n758), .CI(
        DP_mult_205_n743), .CO(DP_mult_205_n740), .S(DP_mult_205_n741) );
  FA_X1 DP_mult_205_U576 ( .A(DP_mult_205_n754), .B(DP_mult_205_n745), .CI(
        DP_mult_205_n752), .CO(DP_mult_205_n738), .S(DP_mult_205_n739) );
  FA_X1 DP_mult_205_U575 ( .A(DP_mult_205_n750), .B(DP_mult_205_n741), .CI(
        DP_mult_205_n739), .CO(DP_mult_205_n736), .S(DP_mult_205_n737) );
  FA_X1 DP_mult_205_U574 ( .A(DP_mult_205_n746), .B(DP_mult_205_n1203), .CI(
        DP_mult_205_n1247), .CO(DP_mult_205_n734), .S(DP_mult_205_n735) );
  FA_X1 DP_mult_205_U573 ( .A(DP_mult_205_n1225), .B(DP_mult_205_n1291), .CI(
        DP_mult_205_n1269), .CO(DP_mult_205_n732), .S(DP_mult_205_n733) );
  FA_X1 DP_mult_205_U572 ( .A(DP_mult_205_n744), .B(DP_mult_205_n1314), .CI(
        DP_mult_205_n742), .CO(DP_mult_205_n730), .S(DP_mult_205_n731) );
  FA_X1 DP_mult_205_U571 ( .A(DP_mult_205_n735), .B(DP_mult_205_n733), .CI(
        DP_mult_205_n740), .CO(DP_mult_205_n728), .S(DP_mult_205_n729) );
  FA_X1 DP_mult_205_U570 ( .A(DP_mult_205_n738), .B(DP_mult_205_n731), .CI(
        DP_mult_205_n729), .CO(DP_mult_205_n726), .S(DP_mult_205_n727) );
  FA_X1 DP_mult_205_U568 ( .A(DP_mult_205_n1268), .B(DP_mult_205_n1224), .CI(
        DP_mult_205_n725), .CO(DP_mult_205_n722), .S(DP_mult_205_n723) );
  FA_X1 DP_mult_205_U567 ( .A(DP_mult_205_n1202), .B(DP_mult_205_n1246), .CI(
        DP_mult_205_n734), .CO(DP_mult_205_n720), .S(DP_mult_205_n721) );
  FA_X1 DP_mult_205_U566 ( .A(DP_mult_205_n723), .B(DP_mult_205_n732), .CI(
        DP_mult_205_n730), .CO(DP_mult_205_n718), .S(DP_mult_205_n719) );
  FA_X1 DP_mult_205_U565 ( .A(DP_mult_205_n728), .B(DP_mult_205_n721), .CI(
        DP_mult_205_n719), .CO(DP_mult_205_n716), .S(DP_mult_205_n717) );
  FA_X1 DP_mult_205_U564 ( .A(DP_mult_205_n1267), .B(DP_mult_205_n1201), .CI(
        DP_mult_205_n724), .CO(DP_mult_205_n714), .S(DP_mult_205_n715) );
  FA_X1 DP_mult_205_U563 ( .A(DP_mult_205_n1245), .B(DP_mult_205_n1223), .CI(
        DP_mult_205_n1290), .CO(DP_mult_205_n712), .S(DP_mult_205_n713) );
  FA_X1 DP_mult_205_U562 ( .A(DP_mult_205_n715), .B(DP_mult_205_n722), .CI(
        DP_mult_205_n720), .CO(DP_mult_205_n710), .S(DP_mult_205_n711) );
  FA_X1 DP_mult_205_U561 ( .A(DP_mult_205_n718), .B(DP_mult_205_n713), .CI(
        DP_mult_205_n711), .CO(DP_mult_205_n708), .S(DP_mult_205_n709) );
  FA_X1 DP_mult_205_U559 ( .A(DP_mult_205_n1222), .B(DP_mult_205_n1200), .CI(
        DP_mult_205_n707), .CO(DP_mult_205_n704), .S(DP_mult_205_n705) );
  FA_X1 DP_mult_205_U558 ( .A(DP_mult_205_n714), .B(DP_mult_205_n1244), .CI(
        DP_mult_205_n705), .CO(DP_mult_205_n702), .S(DP_mult_205_n703) );
  FA_X1 DP_mult_205_U557 ( .A(DP_mult_205_n710), .B(DP_mult_205_n712), .CI(
        DP_mult_205_n703), .CO(DP_mult_205_n700), .S(DP_mult_205_n701) );
  FA_X1 DP_mult_205_U556 ( .A(DP_mult_205_n1221), .B(DP_mult_205_n1199), .CI(
        DP_mult_205_n706), .CO(DP_mult_205_n698), .S(DP_mult_205_n699) );
  FA_X1 DP_mult_205_U555 ( .A(DP_mult_205_n1266), .B(DP_mult_205_n1243), .CI(
        DP_mult_205_n704), .CO(DP_mult_205_n696), .S(DP_mult_205_n697) );
  FA_X1 DP_mult_205_U554 ( .A(DP_mult_205_n702), .B(DP_mult_205_n699), .CI(
        DP_mult_205_n697), .CO(DP_mult_205_n694), .S(DP_mult_205_n695) );
  FA_X1 DP_mult_205_U552 ( .A(DP_mult_205_n1198), .B(DP_mult_205_n1220), .CI(
        DP_mult_205_n693), .CO(DP_mult_205_n690), .S(DP_mult_205_n691) );
  FA_X1 DP_mult_205_U551 ( .A(DP_mult_205_n691), .B(DP_mult_205_n698), .CI(
        DP_mult_205_n696), .CO(DP_mult_205_n688), .S(DP_mult_205_n689) );
  FA_X1 DP_mult_205_U550 ( .A(DP_mult_205_n1219), .B(DP_mult_205_n692), .CI(
        DP_mult_205_n1197), .CO(DP_mult_205_n686), .S(DP_mult_205_n687) );
  FA_X1 DP_mult_205_U549 ( .A(DP_mult_205_n690), .B(DP_mult_205_n1242), .CI(
        DP_mult_205_n687), .CO(DP_mult_205_n684), .S(DP_mult_205_n685) );
  FA_X1 DP_mult_205_U547 ( .A(DP_mult_205_n683), .B(DP_mult_205_n1196), .CI(
        DP_mult_205_n686), .CO(DP_mult_205_n680), .S(DP_mult_205_n681) );
  FA_X1 DP_mult_205_U546 ( .A(DP_mult_205_n1195), .B(DP_mult_205_n682), .CI(
        DP_mult_205_n1218), .CO(DP_mult_205_n678), .S(DP_mult_205_n679) );
  INV_X1 DP_mult_204_U2901 ( .A(DP_mult_204_n2210), .ZN(DP_mult_204_n2360) );
  INV_X1 DP_mult_204_U2900 ( .A(DP_mult_204_n2207), .ZN(DP_mult_204_n2357) );
  INV_X1 DP_mult_204_U2899 ( .A(DP_mult_204_n2203), .ZN(DP_mult_204_n2354) );
  INV_X1 DP_mult_204_U2898 ( .A(DP_mult_204_n2243), .ZN(DP_mult_204_n2338) );
  INV_X2 DP_mult_204_U2897 ( .A(DP_mult_204_n1987), .ZN(DP_mult_204_n2311) );
  XNOR2_X1 DP_mult_204_U2896 ( .A(DP_sw0_17_), .B(DP_mult_204_n2351), .ZN(
        DP_mult_204_n1713) );
  XNOR2_X1 DP_mult_204_U2895 ( .A(DP_sw0_19_), .B(DP_mult_204_n2350), .ZN(
        DP_mult_204_n1711) );
  XNOR2_X1 DP_mult_204_U2894 ( .A(DP_sw0_11_), .B(DP_mult_204_n2351), .ZN(
        DP_mult_204_n1719) );
  XNOR2_X1 DP_mult_204_U2893 ( .A(DP_sw0_15_), .B(DP_mult_204_n2350), .ZN(
        DP_mult_204_n1715) );
  XNOR2_X1 DP_mult_204_U2892 ( .A(DP_sw0_21_), .B(DP_mult_204_n2351), .ZN(
        DP_mult_204_n1709) );
  OAI22_X1 DP_mult_204_U2891 ( .A1(DP_mult_204_n2313), .A2(DP_mult_204_n1683), 
        .B1(DP_mult_204_n1682), .B2(DP_mult_204_n2338), .ZN(DP_mult_204_n836)
         );
  XNOR2_X1 DP_mult_204_U2890 ( .A(DP_sw0_13_), .B(DP_mult_204_n2350), .ZN(
        DP_mult_204_n1717) );
  OAI22_X1 DP_mult_204_U2889 ( .A1(DP_mult_204_n1706), .A2(DP_mult_204_n2338), 
        .B1(DP_mult_204_n2185), .B2(DP_mult_204_n2203), .ZN(DP_mult_204_n1190)
         );
  OAI22_X1 DP_mult_204_U2888 ( .A1(DP_mult_204_n2313), .A2(DP_mult_204_n1693), 
        .B1(DP_mult_204_n1692), .B2(DP_mult_204_n2337), .ZN(DP_mult_204_n1396)
         );
  OAI22_X1 DP_mult_204_U2887 ( .A1(DP_mult_204_n2314), .A2(DP_mult_204_n1684), 
        .B1(DP_mult_204_n2338), .B2(DP_mult_204_n1683), .ZN(DP_mult_204_n1387)
         );
  INV_X1 DP_mult_204_U2886 ( .A(DP_mult_204_n836), .ZN(DP_mult_204_n837) );
  OAI22_X1 DP_mult_204_U2885 ( .A1(DP_mult_204_n2314), .A2(DP_mult_204_n1688), 
        .B1(DP_mult_204_n2338), .B2(DP_mult_204_n1687), .ZN(DP_mult_204_n1391)
         );
  OAI22_X1 DP_mult_204_U2884 ( .A1(DP_mult_204_n2186), .A2(DP_mult_204_n1685), 
        .B1(DP_mult_204_n1684), .B2(DP_mult_204_n2337), .ZN(DP_mult_204_n1388)
         );
  OAI22_X1 DP_mult_204_U2883 ( .A1(DP_mult_204_n2186), .A2(DP_mult_204_n1692), 
        .B1(DP_mult_204_n2337), .B2(DP_mult_204_n1691), .ZN(DP_mult_204_n1395)
         );
  OAI22_X1 DP_mult_204_U2882 ( .A1(DP_mult_204_n2186), .A2(DP_mult_204_n1687), 
        .B1(DP_mult_204_n1686), .B2(DP_mult_204_n2338), .ZN(DP_mult_204_n1390)
         );
  OAI22_X1 DP_mult_204_U2881 ( .A1(DP_mult_204_n2185), .A2(DP_mult_204_n1690), 
        .B1(DP_mult_204_n2338), .B2(DP_mult_204_n1689), .ZN(DP_mult_204_n1393)
         );
  OAI22_X1 DP_mult_204_U2880 ( .A1(DP_mult_204_n2314), .A2(DP_mult_204_n1689), 
        .B1(DP_mult_204_n1688), .B2(DP_mult_204_n2338), .ZN(DP_mult_204_n1392)
         );
  OAI22_X1 DP_mult_204_U2879 ( .A1(DP_mult_204_n2186), .A2(DP_mult_204_n1686), 
        .B1(DP_mult_204_n2338), .B2(DP_mult_204_n1685), .ZN(DP_mult_204_n1389)
         );
  OAI22_X1 DP_mult_204_U2878 ( .A1(DP_mult_204_n2314), .A2(DP_mult_204_n1691), 
        .B1(DP_mult_204_n1690), .B2(DP_mult_204_n2337), .ZN(DP_mult_204_n1394)
         );
  NAND2_X1 DP_mult_204_U2877 ( .A1(DP_mult_204_n775), .A2(DP_mult_204_n788), 
        .ZN(DP_mult_204_n474) );
  OAI21_X1 DP_mult_204_U2876 ( .B1(DP_mult_204_n2148), .B2(DP_mult_204_n398), 
        .A(DP_mult_204_n399), .ZN(DP_mult_204_n397) );
  OAI21_X1 DP_mult_204_U2875 ( .B1(DP_mult_204_n2218), .B2(DP_mult_204_n389), 
        .A(DP_mult_204_n390), .ZN(DP_mult_204_n388) );
  OAI21_X1 DP_mult_204_U2874 ( .B1(DP_mult_204_n2219), .B2(DP_mult_204_n431), 
        .A(DP_mult_204_n432), .ZN(DP_mult_204_n430) );
  OAI21_X1 DP_mult_204_U2873 ( .B1(DP_mult_204_n2218), .B2(DP_mult_204_n411), 
        .A(DP_mult_204_n412), .ZN(DP_mult_204_n410) );
  OAI21_X1 DP_mult_204_U2872 ( .B1(DP_mult_204_n2003), .B2(DP_mult_204_n420), 
        .A(DP_mult_204_n421), .ZN(DP_mult_204_n419) );
  OAI21_X1 DP_mult_204_U2871 ( .B1(DP_mult_204_n2148), .B2(DP_mult_204_n343), 
        .A(DP_mult_204_n344), .ZN(DP_mult_204_n342) );
  OAI21_X1 DP_mult_204_U2870 ( .B1(DP_mult_204_n2218), .B2(DP_mult_204_n380), 
        .A(DP_mult_204_n381), .ZN(DP_mult_204_n379) );
  OAI21_X1 DP_mult_204_U2869 ( .B1(DP_mult_204_n2219), .B2(DP_mult_204_n371), 
        .A(DP_mult_204_n372), .ZN(DP_mult_204_n370) );
  OAI21_X1 DP_mult_204_U2868 ( .B1(DP_mult_204_n2148), .B2(DP_mult_204_n354), 
        .A(DP_mult_204_n355), .ZN(DP_mult_204_n353) );
  OAI21_X1 DP_mult_204_U2867 ( .B1(DP_mult_204_n2003), .B2(DP_mult_204_n438), 
        .A(DP_mult_204_n439), .ZN(DP_mult_204_n437) );
  OAI21_X1 DP_mult_204_U2866 ( .B1(DP_mult_204_n2219), .B2(DP_mult_204_n326), 
        .A(DP_mult_204_n327), .ZN(DP_mult_204_n325) );
  XNOR2_X1 DP_mult_204_U2865 ( .A(DP_mult_204_n437), .B(DP_mult_204_n311), 
        .ZN(DP_sw0_coeff_ret0[13]) );
  XNOR2_X1 DP_mult_204_U2864 ( .A(DP_sw0_13_), .B(DP_mult_204_n1935), .ZN(
        DP_mult_204_n1742) );
  XNOR2_X1 DP_mult_204_U2863 ( .A(DP_sw0_17_), .B(DP_mult_204_n1935), .ZN(
        DP_mult_204_n1738) );
  XNOR2_X1 DP_mult_204_U2862 ( .A(DP_sw0_11_), .B(DP_mult_204_n2348), .ZN(
        DP_mult_204_n1744) );
  XNOR2_X1 DP_mult_204_U2861 ( .A(DP_sw0_19_), .B(DP_mult_204_n1935), .ZN(
        DP_mult_204_n1736) );
  XNOR2_X1 DP_mult_204_U2860 ( .A(DP_sw0_15_), .B(DP_mult_204_n2348), .ZN(
        DP_mult_204_n1740) );
  OAI22_X1 DP_mult_204_U2859 ( .A1(DP_mult_204_n2316), .A2(DP_mult_204_n1724), 
        .B1(DP_mult_204_n1723), .B2(DP_mult_204_n2341), .ZN(DP_mult_204_n1426)
         );
  XNOR2_X1 DP_mult_204_U2858 ( .A(DP_sw0_21_), .B(DP_mult_204_n1935), .ZN(
        DP_mult_204_n1734) );
  OAI22_X1 DP_mult_204_U2857 ( .A1(DP_mult_204_n2316), .A2(DP_mult_204_n1719), 
        .B1(DP_mult_204_n2340), .B2(DP_mult_204_n1718), .ZN(DP_mult_204_n1421)
         );
  OAI22_X1 DP_mult_204_U2856 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1722), 
        .B1(DP_mult_204_n1721), .B2(DP_mult_204_n2341), .ZN(DP_mult_204_n1424)
         );
  OAI22_X1 DP_mult_204_U2855 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1729), 
        .B1(DP_mult_204_n2341), .B2(DP_mult_204_n1728), .ZN(DP_mult_204_n1431)
         );
  OAI22_X1 DP_mult_204_U2854 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1728), 
        .B1(DP_mult_204_n1727), .B2(DP_mult_204_n2340), .ZN(DP_mult_204_n1430)
         );
  OAI22_X1 DP_mult_204_U2853 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1723), 
        .B1(DP_mult_204_n2341), .B2(DP_mult_204_n1722), .ZN(DP_mult_204_n1425)
         );
  OAI22_X1 DP_mult_204_U2852 ( .A1(DP_mult_204_n2316), .A2(DP_mult_204_n1725), 
        .B1(DP_mult_204_n2340), .B2(DP_mult_204_n1724), .ZN(DP_mult_204_n1427)
         );
  OAI22_X1 DP_mult_204_U2851 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1730), 
        .B1(DP_mult_204_n1729), .B2(DP_mult_204_n2340), .ZN(DP_mult_204_n1432)
         );
  OAI22_X1 DP_mult_204_U2850 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1726), 
        .B1(DP_mult_204_n1725), .B2(DP_mult_204_n2340), .ZN(DP_mult_204_n1428)
         );
  OAI22_X1 DP_mult_204_U2849 ( .A1(DP_mult_204_n2316), .A2(DP_mult_204_n1721), 
        .B1(DP_mult_204_n2340), .B2(DP_mult_204_n1720), .ZN(DP_mult_204_n1423)
         );
  OAI22_X1 DP_mult_204_U2848 ( .A1(DP_mult_204_n2316), .A2(DP_mult_204_n1720), 
        .B1(DP_mult_204_n1719), .B2(DP_mult_204_n2341), .ZN(DP_mult_204_n1422)
         );
  OAI22_X1 DP_mult_204_U2847 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1727), 
        .B1(DP_mult_204_n2341), .B2(DP_mult_204_n1726), .ZN(DP_mult_204_n1429)
         );
  OAI21_X1 DP_mult_204_U2846 ( .B1(DP_mult_204_n536), .B2(DP_mult_204_n498), 
        .A(DP_mult_204_n499), .ZN(DP_mult_204_n497) );
  OAI21_X1 DP_mult_204_U2845 ( .B1(DP_mult_204_n536), .B2(DP_mult_204_n2251), 
        .A(DP_mult_204_n2208), .ZN(DP_mult_204_n504) );
  OAI21_X1 DP_mult_204_U2844 ( .B1(DP_mult_204_n536), .B2(DP_mult_204_n516), 
        .A(DP_mult_204_n517), .ZN(DP_mult_204_n515) );
  OAI21_X1 DP_mult_204_U2843 ( .B1(DP_mult_204_n536), .B2(DP_mult_204_n476), 
        .A(DP_mult_204_n477), .ZN(DP_mult_204_n475) );
  OAI21_X1 DP_mult_204_U2842 ( .B1(DP_mult_204_n536), .B2(DP_mult_204_n2271), 
        .A(DP_mult_204_n524), .ZN(DP_mult_204_n522) );
  OAI21_X1 DP_mult_204_U2841 ( .B1(DP_mult_204_n536), .B2(DP_mult_204_n463), 
        .A(DP_mult_204_n464), .ZN(DP_mult_204_n462) );
  OAI21_X1 DP_mult_204_U2840 ( .B1(DP_mult_204_n536), .B2(DP_mult_204_n487), 
        .A(DP_mult_204_n488), .ZN(DP_mult_204_n486) );
  OAI21_X1 DP_mult_204_U2839 ( .B1(DP_mult_204_n536), .B2(DP_mult_204_n534), 
        .A(DP_mult_204_n535), .ZN(DP_mult_204_n533) );
  AOI21_X1 DP_mult_204_U2838 ( .B1(DP_mult_204_n333), .B2(DP_mult_204_n1996), 
        .A(DP_mult_204_n2240), .ZN(DP_mult_204_n327) );
  NAND2_X1 DP_mult_204_U2837 ( .A1(DP_mult_204_n356), .A2(DP_mult_204_n2238), 
        .ZN(DP_mult_204_n347) );
  XNOR2_X1 DP_mult_204_U2836 ( .A(DP_sw0_11_), .B(DP_mult_204_n2346), .ZN(
        DP_mult_204_n1769) );
  XNOR2_X1 DP_mult_204_U2835 ( .A(DP_sw0_15_), .B(DP_mult_204_n2346), .ZN(
        DP_mult_204_n1765) );
  XNOR2_X1 DP_mult_204_U2834 ( .A(DP_sw0_19_), .B(DP_mult_204_n2346), .ZN(
        DP_mult_204_n1761) );
  XNOR2_X1 DP_mult_204_U2833 ( .A(DP_sw0_13_), .B(DP_mult_204_n2346), .ZN(
        DP_mult_204_n1767) );
  XNOR2_X1 DP_mult_204_U2832 ( .A(DP_sw0_21_), .B(DP_mult_204_n2346), .ZN(
        DP_mult_204_n1759) );
  OAI22_X1 DP_mult_204_U2831 ( .A1(DP_mult_204_n2317), .A2(DP_mult_204_n1733), 
        .B1(DP_mult_204_n2155), .B2(DP_mult_204_n1956), .ZN(DP_mult_204_n916)
         );
  XNOR2_X1 DP_mult_204_U2830 ( .A(DP_sw0_17_), .B(DP_mult_204_n2346), .ZN(
        DP_mult_204_n1763) );
  OAI22_X1 DP_mult_204_U2829 ( .A1(DP_mult_204_n2278), .A2(DP_mult_204_n1742), 
        .B1(DP_mult_204_n2342), .B2(DP_mult_204_n1741), .ZN(DP_mult_204_n1443)
         );
  OAI22_X1 DP_mult_204_U2828 ( .A1(DP_mult_204_n2279), .A2(DP_mult_204_n1737), 
        .B1(DP_mult_204_n1736), .B2(DP_mult_204_n2342), .ZN(DP_mult_204_n1438)
         );
  OAI22_X1 DP_mult_204_U2827 ( .A1(DP_mult_204_n2317), .A2(DP_mult_204_n1743), 
        .B1(DP_mult_204_n1742), .B2(DP_mult_204_n2342), .ZN(DP_mult_204_n1444)
         );
  OAI22_X1 DP_mult_204_U2826 ( .A1(DP_mult_204_n2278), .A2(DP_mult_204_n1734), 
        .B1(DP_mult_204_n2342), .B2(DP_mult_204_n1733), .ZN(DP_mult_204_n1435)
         );
  OAI22_X1 DP_mult_204_U2825 ( .A1(DP_mult_204_n2278), .A2(DP_mult_204_n1739), 
        .B1(DP_mult_204_n1738), .B2(DP_mult_204_n2342), .ZN(DP_mult_204_n1440)
         );
  OAI22_X1 DP_mult_204_U2824 ( .A1(DP_mult_204_n2279), .A2(DP_mult_204_n1735), 
        .B1(DP_mult_204_n1734), .B2(DP_mult_204_n2155), .ZN(DP_mult_204_n1436)
         );
  OAI22_X1 DP_mult_204_U2823 ( .A1(DP_mult_204_n2318), .A2(DP_mult_204_n1736), 
        .B1(DP_mult_204_n2342), .B2(DP_mult_204_n1735), .ZN(DP_mult_204_n1437)
         );
  OAI22_X1 DP_mult_204_U2822 ( .A1(DP_mult_204_n2279), .A2(DP_mult_204_n1740), 
        .B1(DP_mult_204_n2342), .B2(DP_mult_204_n1739), .ZN(DP_mult_204_n1441)
         );
  OAI22_X1 DP_mult_204_U2821 ( .A1(DP_mult_204_n2279), .A2(DP_mult_204_n1741), 
        .B1(DP_mult_204_n1740), .B2(DP_mult_204_n2342), .ZN(DP_mult_204_n1442)
         );
  OAI22_X1 DP_mult_204_U2820 ( .A1(DP_mult_204_n2278), .A2(DP_mult_204_n1738), 
        .B1(DP_mult_204_n1978), .B2(DP_mult_204_n1737), .ZN(DP_mult_204_n1439)
         );
  OAI22_X1 DP_mult_204_U2819 ( .A1(DP_mult_204_n1756), .A2(DP_mult_204_n1978), 
        .B1(DP_mult_204_n2278), .B2(DP_mult_204_n2349), .ZN(DP_mult_204_n1192)
         );
  INV_X1 DP_mult_204_U2818 ( .A(DP_mult_204_n2093), .ZN(DP_mult_204_n492) );
  AOI21_X1 DP_mult_204_U2817 ( .B1(DP_mult_204_n508), .B2(DP_mult_204_n489), 
        .A(DP_mult_204_n2093), .ZN(DP_mult_204_n488) );
  XNOR2_X1 DP_mult_204_U2816 ( .A(DP_sw0_13_), .B(DP_mult_204_n2134), .ZN(
        DP_mult_204_n1642) );
  XNOR2_X1 DP_mult_204_U2815 ( .A(DP_sw0_15_), .B(DP_mult_204_n2135), .ZN(
        DP_mult_204_n1640) );
  XNOR2_X1 DP_mult_204_U2814 ( .A(DP_sw0_11_), .B(DP_mult_204_n2360), .ZN(
        DP_mult_204_n1644) );
  XNOR2_X1 DP_mult_204_U2813 ( .A(DP_sw0_17_), .B(DP_mult_204_n2134), .ZN(
        DP_mult_204_n1638) );
  OAI22_X1 DP_mult_204_U2812 ( .A1(DP_mult_204_n2308), .A2(DP_mult_204_n1628), 
        .B1(DP_mult_204_n1627), .B2(DP_mult_204_n1970), .ZN(DP_mult_204_n1334)
         );
  XNOR2_X1 DP_mult_204_U2811 ( .A(DP_sw0_21_), .B(DP_mult_204_n2135), .ZN(
        DP_mult_204_n1634) );
  OAI22_X1 DP_mult_204_U2810 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1622), 
        .B1(DP_mult_204_n1621), .B2(DP_mult_204_n1969), .ZN(DP_mult_204_n1328)
         );
  OAI22_X1 DP_mult_204_U2809 ( .A1(DP_mult_204_n2070), .A2(DP_mult_204_n1627), 
        .B1(DP_mult_204_n1969), .B2(DP_mult_204_n1626), .ZN(DP_mult_204_n1333)
         );
  OAI22_X1 DP_mult_204_U2808 ( .A1(DP_mult_204_n2070), .A2(DP_mult_204_n1624), 
        .B1(DP_mult_204_n1623), .B2(DP_mult_204_n1969), .ZN(DP_mult_204_n1330)
         );
  OAI22_X1 DP_mult_204_U2807 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1619), 
        .B1(DP_mult_204_n1969), .B2(DP_mult_204_n1618), .ZN(DP_mult_204_n1325)
         );
  XNOR2_X1 DP_mult_204_U2806 ( .A(DP_sw0_19_), .B(DP_mult_204_n2360), .ZN(
        DP_mult_204_n1636) );
  OAI22_X1 DP_mult_204_U2805 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1621), 
        .B1(DP_mult_204_n1969), .B2(DP_mult_204_n1620), .ZN(DP_mult_204_n1327)
         );
  OAI22_X1 DP_mult_204_U2804 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1625), 
        .B1(DP_mult_204_n1970), .B2(DP_mult_204_n1624), .ZN(DP_mult_204_n1331)
         );
  OAI22_X1 DP_mult_204_U2803 ( .A1(DP_mult_204_n1967), .A2(DP_mult_204_n1629), 
        .B1(DP_mult_204_n1970), .B2(DP_mult_204_n1628), .ZN(DP_mult_204_n1335)
         );
  OAI22_X1 DP_mult_204_U2802 ( .A1(DP_mult_204_n1967), .A2(DP_mult_204_n1630), 
        .B1(DP_mult_204_n1629), .B2(DP_mult_204_n2333), .ZN(DP_mult_204_n1336)
         );
  OAI22_X1 DP_mult_204_U2801 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1623), 
        .B1(DP_mult_204_n1970), .B2(DP_mult_204_n1622), .ZN(DP_mult_204_n1329)
         );
  OAI22_X1 DP_mult_204_U2800 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1626), 
        .B1(DP_mult_204_n1625), .B2(DP_mult_204_n1969), .ZN(DP_mult_204_n1332)
         );
  OAI22_X1 DP_mult_204_U2799 ( .A1(DP_mult_204_n1967), .A2(DP_mult_204_n1620), 
        .B1(DP_mult_204_n1619), .B2(DP_mult_204_n1969), .ZN(DP_mult_204_n1326)
         );
  OAI21_X1 DP_mult_204_U2798 ( .B1(DP_mult_204_n572), .B2(DP_mult_204_n2046), 
        .A(DP_mult_204_n570), .ZN(DP_mult_204_n568) );
  XNOR2_X1 DP_mult_204_U2797 ( .A(DP_mult_204_n430), .B(DP_mult_204_n310), 
        .ZN(DP_sw0_coeff_ret0[14]) );
  XNOR2_X1 DP_mult_204_U2796 ( .A(DP_sw0_13_), .B(DP_mult_204_n2355), .ZN(
        DP_mult_204_n1667) );
  XNOR2_X1 DP_mult_204_U2795 ( .A(DP_sw0_21_), .B(DP_mult_204_n2357), .ZN(
        DP_mult_204_n1659) );
  XNOR2_X1 DP_mult_204_U2794 ( .A(DP_sw0_15_), .B(DP_mult_204_n2355), .ZN(
        DP_mult_204_n1665) );
  XNOR2_X1 DP_mult_204_U2793 ( .A(DP_sw0_19_), .B(DP_mult_204_n2357), .ZN(
        DP_mult_204_n1661) );
  XNOR2_X1 DP_mult_204_U2792 ( .A(DP_sw0_17_), .B(DP_mult_204_n2355), .ZN(
        DP_mult_204_n1663) );
  OAI22_X1 DP_mult_204_U2791 ( .A1(DP_mult_204_n1656), .A2(DP_mult_204_n2334), 
        .B1(DP_mult_204_n2206), .B2(DP_mult_204_n2210), .ZN(DP_mult_204_n1188)
         );
  XNOR2_X1 DP_mult_204_U2790 ( .A(DP_sw0_11_), .B(DP_mult_204_n2355), .ZN(
        DP_mult_204_n1669) );
  OAI22_X1 DP_mult_204_U2789 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1643), 
        .B1(DP_mult_204_n1642), .B2(DP_mult_204_n2334), .ZN(DP_mult_204_n1348)
         );
  OAI22_X1 DP_mult_204_U2788 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1641), 
        .B1(DP_mult_204_n1640), .B2(DP_mult_204_n2334), .ZN(DP_mult_204_n1346)
         );
  OAI22_X1 DP_mult_204_U2787 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1642), 
        .B1(DP_mult_204_n2334), .B2(DP_mult_204_n1641), .ZN(DP_mult_204_n1347)
         );
  OAI22_X1 DP_mult_204_U2786 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1633), 
        .B1(DP_mult_204_n1632), .B2(DP_mult_204_n2334), .ZN(DP_mult_204_n772)
         );
  OAI22_X1 DP_mult_204_U2785 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1638), 
        .B1(DP_mult_204_n2334), .B2(DP_mult_204_n1637), .ZN(DP_mult_204_n1343)
         );
  OAI22_X1 DP_mult_204_U2784 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1640), 
        .B1(DP_mult_204_n2042), .B2(DP_mult_204_n1639), .ZN(DP_mult_204_n1345)
         );
  OAI22_X1 DP_mult_204_U2783 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1639), 
        .B1(DP_mult_204_n1638), .B2(DP_mult_204_n2334), .ZN(DP_mult_204_n1344)
         );
  OAI22_X1 DP_mult_204_U2782 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1635), 
        .B1(DP_mult_204_n1634), .B2(DP_mult_204_n2118), .ZN(DP_mult_204_n1340)
         );
  OAI22_X1 DP_mult_204_U2781 ( .A1(DP_mult_204_n2140), .A2(DP_mult_204_n1634), 
        .B1(DP_mult_204_n2042), .B2(DP_mult_204_n1633), .ZN(DP_mult_204_n1339)
         );
  OAI22_X1 DP_mult_204_U2780 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1636), 
        .B1(DP_mult_204_n2042), .B2(DP_mult_204_n1635), .ZN(DP_mult_204_n1341)
         );
  OAI22_X1 DP_mult_204_U2779 ( .A1(DP_mult_204_n2206), .A2(DP_mult_204_n1637), 
        .B1(DP_mult_204_n1636), .B2(DP_mult_204_n2118), .ZN(DP_mult_204_n1342)
         );
  XNOR2_X1 DP_mult_204_U2778 ( .A(DP_mult_204_n419), .B(DP_mult_204_n309), 
        .ZN(DP_sw0_coeff_ret0[15]) );
  XNOR2_X1 DP_mult_204_U2777 ( .A(DP_sw0_15_), .B(DP_mult_204_n2377), .ZN(
        DP_mult_204_n1515) );
  XNOR2_X1 DP_mult_204_U2776 ( .A(DP_sw0_13_), .B(DP_mult_204_n2377), .ZN(
        DP_mult_204_n1517) );
  XNOR2_X1 DP_mult_204_U2775 ( .A(DP_sw0_19_), .B(DP_mult_204_n2378), .ZN(
        DP_mult_204_n1511) );
  XNOR2_X1 DP_mult_204_U2774 ( .A(DP_sw0_17_), .B(DP_mult_204_n2377), .ZN(
        DP_mult_204_n1513) );
  XNOR2_X1 DP_mult_204_U2773 ( .A(DP_sw0_21_), .B(DP_mult_204_n2379), .ZN(
        DP_mult_204_n1509) );
  XNOR2_X1 DP_mult_204_U2772 ( .A(DP_sw0_11_), .B(DP_mult_204_n2379), .ZN(
        DP_mult_204_n1519) );
  OAI22_X1 DP_mult_204_U2771 ( .A1(DP_mult_204_n2289), .A2(DP_mult_204_n1493), 
        .B1(DP_mult_204_n1492), .B2(DP_mult_204_n2321), .ZN(DP_mult_204_n1204)
         );
  OAI22_X1 DP_mult_204_U2770 ( .A1(DP_mult_204_n1506), .A2(DP_mult_204_n2321), 
        .B1(DP_mult_204_n2005), .B2(DP_mult_204_n2289), .ZN(DP_mult_204_n1182)
         );
  OAI22_X1 DP_mult_204_U2769 ( .A1(DP_mult_204_n2255), .A2(DP_mult_204_n1489), 
        .B1(DP_mult_204_n1488), .B2(DP_mult_204_n2321), .ZN(DP_mult_204_n1200)
         );
  OAI22_X1 DP_mult_204_U2768 ( .A1(DP_mult_204_n2254), .A2(DP_mult_204_n1492), 
        .B1(DP_mult_204_n2322), .B2(DP_mult_204_n1491), .ZN(DP_mult_204_n1203)
         );
  OAI22_X1 DP_mult_204_U2767 ( .A1(DP_mult_204_n2255), .A2(DP_mult_204_n1486), 
        .B1(DP_mult_204_n2321), .B2(DP_mult_204_n1485), .ZN(DP_mult_204_n1197)
         );
  OAI22_X1 DP_mult_204_U2766 ( .A1(DP_mult_204_n2254), .A2(DP_mult_204_n1490), 
        .B1(DP_mult_204_n2322), .B2(DP_mult_204_n1489), .ZN(DP_mult_204_n1201)
         );
  OAI22_X1 DP_mult_204_U2765 ( .A1(DP_mult_204_n2255), .A2(DP_mult_204_n1487), 
        .B1(DP_mult_204_n1486), .B2(DP_mult_204_n2321), .ZN(DP_mult_204_n1198)
         );
  OAI22_X1 DP_mult_204_U2764 ( .A1(DP_mult_204_n2254), .A2(DP_mult_204_n1488), 
        .B1(DP_mult_204_n2322), .B2(DP_mult_204_n1487), .ZN(DP_mult_204_n1199)
         );
  OAI22_X1 DP_mult_204_U2763 ( .A1(DP_mult_204_n2254), .A2(DP_mult_204_n1491), 
        .B1(DP_mult_204_n1490), .B2(DP_mult_204_n2322), .ZN(DP_mult_204_n1202)
         );
  OAI22_X1 DP_mult_204_U2762 ( .A1(DP_mult_204_n2255), .A2(DP_mult_204_n1485), 
        .B1(DP_mult_204_n1484), .B2(DP_mult_204_n2321), .ZN(DP_mult_204_n1196)
         );
  NAND2_X1 DP_mult_204_U2761 ( .A1(DP_mult_204_n717), .A2(DP_mult_204_n726), 
        .ZN(DP_mult_204_n418) );
  OAI22_X1 DP_mult_204_U2760 ( .A1(DP_mult_204_n2254), .A2(DP_mult_204_n1484), 
        .B1(DP_mult_204_n2322), .B2(DP_mult_204_n1483), .ZN(DP_mult_204_n1195)
         );
  OAI22_X1 DP_mult_204_U2759 ( .A1(DP_mult_204_n2255), .A2(DP_mult_204_n1483), 
        .B1(DP_mult_204_n1482), .B2(DP_mult_204_n2321), .ZN(DP_mult_204_n676)
         );
  NAND2_X1 DP_mult_204_U2758 ( .A1(DP_mult_204_n345), .A2(DP_mult_204_n2239), 
        .ZN(DP_mult_204_n336) );
  NAND2_X1 DP_mult_204_U2757 ( .A1(DP_mult_204_n422), .A2(DP_mult_204_n2235), 
        .ZN(DP_mult_204_n411) );
  AOI21_X1 DP_mult_204_U2756 ( .B1(DP_mult_204_n423), .B2(DP_mult_204_n2235), 
        .A(DP_mult_204_n416), .ZN(DP_mult_204_n412) );
  INV_X1 DP_mult_204_U2755 ( .A(DP_mult_204_n345), .ZN(DP_mult_204_n343) );
  NAND2_X1 DP_mult_204_U2754 ( .A1(DP_mult_204_n2235), .A2(DP_mult_204_n418), 
        .ZN(DP_mult_204_n309) );
  INV_X1 DP_mult_204_U2753 ( .A(DP_mult_204_n325), .ZN(DP_sw0_coeff_ret0[23])
         );
  NOR2_X1 DP_mult_204_U2752 ( .A1(DP_mult_204_n505), .A2(DP_mult_204_n452), 
        .ZN(DP_mult_204_n450) );
  XNOR2_X1 DP_mult_204_U2751 ( .A(DP_sw0_17_), .B(DP_mult_204_n2362), .ZN(
        DP_mult_204_n1613) );
  XNOR2_X1 DP_mult_204_U2750 ( .A(DP_sw0_15_), .B(DP_mult_204_n2362), .ZN(
        DP_mult_204_n1615) );
  XNOR2_X1 DP_mult_204_U2749 ( .A(DP_sw0_13_), .B(DP_mult_204_n2363), .ZN(
        DP_mult_204_n1617) );
  XNOR2_X1 DP_mult_204_U2748 ( .A(DP_sw0_21_), .B(DP_mult_204_n2362), .ZN(
        DP_mult_204_n1609) );
  XNOR2_X1 DP_mult_204_U2747 ( .A(DP_sw0_11_), .B(DP_mult_204_n2362), .ZN(
        DP_mult_204_n1619) );
  XNOR2_X1 DP_mult_204_U2746 ( .A(DP_sw0_19_), .B(DP_mult_204_n2364), .ZN(
        DP_mult_204_n1611) );
  OAI22_X1 DP_mult_204_U2745 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1599), 
        .B1(DP_mult_204_n1598), .B2(DP_mult_204_n2332), .ZN(DP_mult_204_n1306)
         );
  OAI22_X1 DP_mult_204_U2744 ( .A1(DP_mult_204_n2307), .A2(DP_mult_204_n1595), 
        .B1(DP_mult_204_n1594), .B2(DP_mult_204_n2331), .ZN(DP_mult_204_n1302)
         );
  OAI22_X1 DP_mult_204_U2743 ( .A1(DP_mult_204_n1977), .A2(DP_mult_204_n1597), 
        .B1(DP_mult_204_n1596), .B2(DP_mult_204_n2331), .ZN(DP_mult_204_n1304)
         );
  OAI22_X1 DP_mult_204_U2742 ( .A1(DP_mult_204_n2307), .A2(DP_mult_204_n1605), 
        .B1(DP_mult_204_n1604), .B2(DP_mult_204_n2332), .ZN(DP_mult_204_n1312)
         );
  OAI22_X1 DP_mult_204_U2741 ( .A1(DP_mult_204_n1977), .A2(DP_mult_204_n1598), 
        .B1(DP_mult_204_n2331), .B2(DP_mult_204_n1597), .ZN(DP_mult_204_n1305)
         );
  OAI22_X1 DP_mult_204_U2740 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1596), 
        .B1(DP_mult_204_n2332), .B2(DP_mult_204_n1595), .ZN(DP_mult_204_n1303)
         );
  OAI22_X1 DP_mult_204_U2739 ( .A1(DP_mult_204_n2306), .A2(DP_mult_204_n1594), 
        .B1(DP_mult_204_n2332), .B2(DP_mult_204_n1593), .ZN(DP_mult_204_n1301)
         );
  OAI22_X1 DP_mult_204_U2738 ( .A1(DP_mult_204_n2306), .A2(DP_mult_204_n1601), 
        .B1(DP_mult_204_n1600), .B2(DP_mult_204_n2332), .ZN(DP_mult_204_n1308)
         );
  OAI22_X1 DP_mult_204_U2737 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1604), 
        .B1(DP_mult_204_n2331), .B2(DP_mult_204_n1603), .ZN(DP_mult_204_n1311)
         );
  OAI22_X1 DP_mult_204_U2736 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1600), 
        .B1(DP_mult_204_n2331), .B2(DP_mult_204_n1599), .ZN(DP_mult_204_n1307)
         );
  OAI22_X1 DP_mult_204_U2735 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1603), 
        .B1(DP_mult_204_n1602), .B2(DP_mult_204_n2331), .ZN(DP_mult_204_n1310)
         );
  OAI22_X1 DP_mult_204_U2734 ( .A1(DP_mult_204_n2306), .A2(DP_mult_204_n1602), 
        .B1(DP_mult_204_n2331), .B2(DP_mult_204_n1601), .ZN(DP_mult_204_n1309)
         );
  XNOR2_X1 DP_mult_204_U2733 ( .A(DP_mult_204_n410), .B(DP_mult_204_n308), 
        .ZN(DP_sw0_coeff_ret0[16]) );
  OAI22_X1 DP_mult_204_U2732 ( .A1(DP_mult_204_n2312), .A2(DP_mult_204_n1668), 
        .B1(DP_mult_204_n1667), .B2(DP_mult_204_n2335), .ZN(DP_mult_204_n1372)
         );
  OAI22_X1 DP_mult_204_U2731 ( .A1(DP_mult_204_n2312), .A2(DP_mult_204_n1659), 
        .B1(DP_mult_204_n2335), .B2(DP_mult_204_n1658), .ZN(DP_mult_204_n1363)
         );
  OAI22_X1 DP_mult_204_U2730 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1658), 
        .B1(DP_mult_204_n1657), .B2(DP_mult_204_n2066), .ZN(DP_mult_204_n802)
         );
  OAI22_X1 DP_mult_204_U2729 ( .A1(DP_mult_204_n2312), .A2(DP_mult_204_n1662), 
        .B1(DP_mult_204_n1661), .B2(DP_mult_204_n2066), .ZN(DP_mult_204_n1366)
         );
  OAI22_X1 DP_mult_204_U2728 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1665), 
        .B1(DP_mult_204_n2335), .B2(DP_mult_204_n1664), .ZN(DP_mult_204_n1369)
         );
  OAI22_X1 DP_mult_204_U2727 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1667), 
        .B1(DP_mult_204_n2335), .B2(DP_mult_204_n1666), .ZN(DP_mult_204_n1371)
         );
  OAI22_X1 DP_mult_204_U2726 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1664), 
        .B1(DP_mult_204_n1663), .B2(DP_mult_204_n2066), .ZN(DP_mult_204_n1368)
         );
  OAI22_X1 DP_mult_204_U2725 ( .A1(DP_mult_204_n1681), .A2(DP_mult_204_n2066), 
        .B1(DP_mult_204_n2311), .B2(DP_mult_204_n2207), .ZN(DP_mult_204_n1189)
         );
  OAI22_X1 DP_mult_204_U2724 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1663), 
        .B1(DP_mult_204_n2335), .B2(DP_mult_204_n1662), .ZN(DP_mult_204_n1367)
         );
  OAI22_X1 DP_mult_204_U2723 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1660), 
        .B1(DP_mult_204_n1659), .B2(DP_mult_204_n2066), .ZN(DP_mult_204_n1364)
         );
  OAI22_X1 DP_mult_204_U2722 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1661), 
        .B1(DP_mult_204_n2069), .B2(DP_mult_204_n1660), .ZN(DP_mult_204_n1365)
         );
  XNOR2_X1 DP_mult_204_U2721 ( .A(DP_mult_204_n397), .B(DP_mult_204_n307), 
        .ZN(DP_sw0_coeff_ret0[17]) );
  XNOR2_X1 DP_mult_204_U2720 ( .A(DP_sw0_11_), .B(DP_mult_204_n2373), .ZN(
        DP_mult_204_n1544) );
  XNOR2_X1 DP_mult_204_U2719 ( .A(DP_sw0_15_), .B(DP_mult_204_n2374), .ZN(
        DP_mult_204_n1540) );
  XNOR2_X1 DP_mult_204_U2718 ( .A(DP_sw0_13_), .B(DP_mult_204_n2374), .ZN(
        DP_mult_204_n1542) );
  XNOR2_X1 DP_mult_204_U2717 ( .A(DP_sw0_17_), .B(DP_mult_204_n2374), .ZN(
        DP_mult_204_n1538) );
  OAI22_X1 DP_mult_204_U2716 ( .A1(DP_mult_204_n2067), .A2(DP_mult_204_n1527), 
        .B1(DP_mult_204_n2324), .B2(DP_mult_204_n1526), .ZN(DP_mult_204_n1237)
         );
  OAI22_X1 DP_mult_204_U2715 ( .A1(DP_mult_204_n2300), .A2(DP_mult_204_n1530), 
        .B1(DP_mult_204_n1529), .B2(DP_mult_204_n2325), .ZN(DP_mult_204_n1240)
         );
  OAI22_X1 DP_mult_204_U2714 ( .A1(DP_mult_204_n2068), .A2(DP_mult_204_n1526), 
        .B1(DP_mult_204_n1525), .B2(DP_mult_204_n2325), .ZN(DP_mult_204_n1236)
         );
  OAI22_X1 DP_mult_204_U2713 ( .A1(DP_mult_204_n2068), .A2(DP_mult_204_n1524), 
        .B1(DP_mult_204_n1523), .B2(DP_mult_204_n2324), .ZN(DP_mult_204_n1234)
         );
  OAI22_X1 DP_mult_204_U2712 ( .A1(DP_mult_204_n2067), .A2(DP_mult_204_n1529), 
        .B1(DP_mult_204_n2324), .B2(DP_mult_204_n1528), .ZN(DP_mult_204_n1239)
         );
  OAI22_X1 DP_mult_204_U2711 ( .A1(DP_mult_204_n2067), .A2(DP_mult_204_n1523), 
        .B1(DP_mult_204_n2324), .B2(DP_mult_204_n1522), .ZN(DP_mult_204_n1233)
         );
  OAI22_X1 DP_mult_204_U2710 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1525), 
        .B1(DP_mult_204_n2325), .B2(DP_mult_204_n1524), .ZN(DP_mult_204_n1235)
         );
  OAI22_X1 DP_mult_204_U2709 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1520), 
        .B1(DP_mult_204_n1519), .B2(DP_mult_204_n2324), .ZN(DP_mult_204_n1230)
         );
  XNOR2_X1 DP_mult_204_U2708 ( .A(DP_sw0_21_), .B(DP_mult_204_n2374), .ZN(
        DP_mult_204_n1534) );
  OAI22_X1 DP_mult_204_U2707 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1519), 
        .B1(DP_mult_204_n2324), .B2(DP_mult_204_n1518), .ZN(DP_mult_204_n1229)
         );
  XNOR2_X1 DP_mult_204_U2706 ( .A(DP_sw0_19_), .B(DP_mult_204_n2374), .ZN(
        DP_mult_204_n1536) );
  OAI22_X1 DP_mult_204_U2705 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1521), 
        .B1(DP_mult_204_n2325), .B2(DP_mult_204_n1520), .ZN(DP_mult_204_n1231)
         );
  OAI22_X1 DP_mult_204_U2704 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1522), 
        .B1(DP_mult_204_n1521), .B2(DP_mult_204_n2325), .ZN(DP_mult_204_n1232)
         );
  XNOR2_X1 DP_mult_204_U2703 ( .A(DP_mult_204_n388), .B(DP_mult_204_n306), 
        .ZN(DP_sw0_coeff_ret0[18]) );
  OAI22_X1 DP_mult_204_U2702 ( .A1(DP_mult_204_n2305), .A2(DP_mult_204_n1576), 
        .B1(DP_mult_204_n1575), .B2(DP_mult_204_n2328), .ZN(DP_mult_204_n1284)
         );
  OAI22_X1 DP_mult_204_U2701 ( .A1(DP_mult_204_n2305), .A2(DP_mult_204_n1574), 
        .B1(DP_mult_204_n1573), .B2(DP_mult_204_n2328), .ZN(DP_mult_204_n1282)
         );
  OAI22_X1 DP_mult_204_U2700 ( .A1(DP_mult_204_n2305), .A2(DP_mult_204_n1572), 
        .B1(DP_mult_204_n1571), .B2(DP_mult_204_n2328), .ZN(DP_mult_204_n1280)
         );
  OAI22_X1 DP_mult_204_U2699 ( .A1(DP_mult_204_n2305), .A2(DP_mult_204_n1577), 
        .B1(DP_mult_204_n2329), .B2(DP_mult_204_n1576), .ZN(DP_mult_204_n1285)
         );
  OAI22_X1 DP_mult_204_U2698 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1578), 
        .B1(DP_mult_204_n1577), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n1286)
         );
  OAI22_X1 DP_mult_204_U2697 ( .A1(DP_mult_204_n2305), .A2(DP_mult_204_n1569), 
        .B1(DP_mult_204_n2328), .B2(DP_mult_204_n1568), .ZN(DP_mult_204_n1277)
         );
  OAI22_X1 DP_mult_204_U2696 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1573), 
        .B1(DP_mult_204_n2328), .B2(DP_mult_204_n1572), .ZN(DP_mult_204_n1281)
         );
  OAI22_X1 DP_mult_204_U2695 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1575), 
        .B1(DP_mult_204_n2328), .B2(DP_mult_204_n1574), .ZN(DP_mult_204_n1283)
         );
  OAI22_X1 DP_mult_204_U2694 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1570), 
        .B1(DP_mult_204_n1569), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n1278)
         );
  OAI22_X1 DP_mult_204_U2693 ( .A1(DP_mult_204_n2305), .A2(DP_mult_204_n1579), 
        .B1(DP_mult_204_n2329), .B2(DP_mult_204_n1578), .ZN(DP_mult_204_n1287)
         );
  OAI22_X1 DP_mult_204_U2692 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1571), 
        .B1(DP_mult_204_n2329), .B2(DP_mult_204_n1570), .ZN(DP_mult_204_n1279)
         );
  OAI22_X1 DP_mult_204_U2691 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1580), 
        .B1(DP_mult_204_n1579), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n1288)
         );
  NOR2_X1 DP_mult_204_U2690 ( .A1(DP_mult_204_n897), .A2(DP_mult_204_n918), 
        .ZN(DP_mult_204_n534) );
  XNOR2_X1 DP_mult_204_U2689 ( .A(DP_mult_204_n379), .B(DP_mult_204_n305), 
        .ZN(DP_sw0_coeff_ret0[19]) );
  XNOR2_X1 DP_mult_204_U2688 ( .A(DP_sw0_13_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1692) );
  XNOR2_X1 DP_mult_204_U2687 ( .A(DP_sw0_11_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1694) );
  XNOR2_X1 DP_mult_204_U2686 ( .A(DP_sw0_21_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1684) );
  XNOR2_X1 DP_mult_204_U2685 ( .A(DP_sw0_15_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1690) );
  XNOR2_X1 DP_mult_204_U2684 ( .A(DP_sw0_19_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1686) );
  XNOR2_X1 DP_mult_204_U2683 ( .A(DP_sw0_17_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1688) );
  OAI22_X1 DP_mult_204_U2682 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1680), 
        .B1(DP_mult_204_n1679), .B2(DP_mult_204_n2066), .ZN(DP_mult_204_n1384)
         );
  OAI22_X1 DP_mult_204_U2681 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1678), 
        .B1(DP_mult_204_n1677), .B2(DP_mult_204_n2066), .ZN(DP_mult_204_n1382)
         );
  NAND2_X1 DP_mult_204_U2680 ( .A1(DP_mult_204_n761), .A2(DP_mult_204_n774), 
        .ZN(DP_mult_204_n461) );
  XNOR2_X1 DP_mult_204_U2679 ( .A(DP_mult_204_n370), .B(DP_mult_204_n304), 
        .ZN(DP_sw0_coeff_ret0[20]) );
  OAI22_X1 DP_mult_204_U2678 ( .A1(DP_mult_204_n2279), .A2(DP_mult_204_n1755), 
        .B1(DP_mult_204_n1754), .B2(DP_mult_204_n1978), .ZN(DP_mult_204_n1456)
         );
  INV_X1 DP_mult_204_U2677 ( .A(DP_mult_204_n2136), .ZN(DP_mult_204_n917) );
  OAI22_X1 DP_mult_204_U2676 ( .A1(DP_mult_204_n2278), .A2(DP_mult_204_n1753), 
        .B1(DP_mult_204_n1752), .B2(DP_mult_204_n1978), .ZN(DP_mult_204_n1454)
         );
  NAND2_X1 DP_mult_204_U2675 ( .A1(DP_mult_204_n805), .A2(DP_mult_204_n820), 
        .ZN(DP_mult_204_n496) );
  XNOR2_X1 DP_mult_204_U2674 ( .A(DP_mult_204_n353), .B(DP_mult_204_n303), 
        .ZN(DP_sw0_coeff_ret0[21]) );
  OAI22_X1 DP_mult_204_U2673 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1554), 
        .B1(DP_mult_204_n2326), .B2(DP_mult_204_n1553), .ZN(DP_mult_204_n1263)
         );
  OAI22_X1 DP_mult_204_U2672 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1550), 
        .B1(DP_mult_204_n2326), .B2(DP_mult_204_n1549), .ZN(DP_mult_204_n1259)
         );
  OAI22_X1 DP_mult_204_U2671 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1547), 
        .B1(DP_mult_204_n1546), .B2(DP_mult_204_n2327), .ZN(DP_mult_204_n1256)
         );
  OAI22_X1 DP_mult_204_U2670 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1555), 
        .B1(DP_mult_204_n1554), .B2(DP_mult_204_n2327), .ZN(DP_mult_204_n1264)
         );
  OAI22_X1 DP_mult_204_U2669 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1545), 
        .B1(DP_mult_204_n1544), .B2(DP_mult_204_n2326), .ZN(DP_mult_204_n1254)
         );
  OAI22_X1 DP_mult_204_U2668 ( .A1(DP_mult_204_n1548), .A2(DP_mult_204_n2221), 
        .B1(DP_mult_204_n2327), .B2(DP_mult_204_n1547), .ZN(DP_mult_204_n1257)
         );
  OAI22_X1 DP_mult_204_U2667 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1549), 
        .B1(DP_mult_204_n1548), .B2(DP_mult_204_n2327), .ZN(DP_mult_204_n1258)
         );
  OAI22_X1 DP_mult_204_U2666 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1552), 
        .B1(DP_mult_204_n2326), .B2(DP_mult_204_n1551), .ZN(DP_mult_204_n1261)
         );
  OAI22_X1 DP_mult_204_U2665 ( .A1(DP_mult_204_n2010), .A2(DP_mult_204_n1546), 
        .B1(DP_mult_204_n2326), .B2(DP_mult_204_n1545), .ZN(DP_mult_204_n1255)
         );
  OAI22_X1 DP_mult_204_U2664 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1544), 
        .B1(DP_mult_204_n2327), .B2(DP_mult_204_n1543), .ZN(DP_mult_204_n1253)
         );
  XNOR2_X1 DP_mult_204_U2663 ( .A(DP_mult_204_n342), .B(DP_mult_204_n302), 
        .ZN(DP_sw0_coeff_ret0[22]) );
  OAI22_X1 DP_mult_204_U2662 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1568), 
        .B1(DP_mult_204_n1567), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n1276)
         );
  OAI22_X1 DP_mult_204_U2661 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1558), 
        .B1(DP_mult_204_n1557), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n706)
         );
  OAI22_X1 DP_mult_204_U2660 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1562), 
        .B1(DP_mult_204_n1561), .B2(DP_mult_204_n2328), .ZN(DP_mult_204_n1270)
         );
  OAI22_X1 DP_mult_204_U2659 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1564), 
        .B1(DP_mult_204_n1563), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n1272)
         );
  OAI22_X1 DP_mult_204_U2658 ( .A1(DP_mult_204_n2305), .A2(DP_mult_204_n1565), 
        .B1(DP_mult_204_n2328), .B2(DP_mult_204_n1564), .ZN(DP_mult_204_n1273)
         );
  OAI22_X1 DP_mult_204_U2657 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1559), 
        .B1(DP_mult_204_n2329), .B2(DP_mult_204_n1558), .ZN(DP_mult_204_n1267)
         );
  OAI22_X1 DP_mult_204_U2656 ( .A1(DP_mult_204_n1581), .A2(DP_mult_204_n2329), 
        .B1(DP_mult_204_n2304), .B2(DP_mult_204_n2372), .ZN(DP_mult_204_n1185)
         );
  OAI22_X1 DP_mult_204_U2655 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1566), 
        .B1(DP_mult_204_n1565), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n1274)
         );
  OAI22_X1 DP_mult_204_U2654 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1561), 
        .B1(DP_mult_204_n2329), .B2(DP_mult_204_n1560), .ZN(DP_mult_204_n1269)
         );
  OAI22_X1 DP_mult_204_U2653 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1567), 
        .B1(DP_mult_204_n2329), .B2(DP_mult_204_n1566), .ZN(DP_mult_204_n1275)
         );
  OAI22_X1 DP_mult_204_U2652 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1560), 
        .B1(DP_mult_204_n1559), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n1268)
         );
  OAI22_X1 DP_mult_204_U2651 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1563), 
        .B1(DP_mult_204_n2329), .B2(DP_mult_204_n1562), .ZN(DP_mult_204_n1271)
         );
  NOR2_X1 DP_mult_204_U2650 ( .A1(DP_mult_204_n420), .A2(DP_mult_204_n347), 
        .ZN(DP_mult_204_n345) );
  OAI21_X1 DP_mult_204_U2649 ( .B1(DP_mult_204_n421), .B2(DP_mult_204_n347), 
        .A(DP_mult_204_n348), .ZN(DP_mult_204_n346) );
  AOI21_X1 DP_mult_204_U2648 ( .B1(DP_mult_204_n346), .B2(DP_mult_204_n2239), 
        .A(DP_mult_204_n339), .ZN(DP_mult_204_n337) );
  AOI21_X1 DP_mult_204_U2647 ( .B1(DP_mult_204_n383), .B2(DP_mult_204_n2234), 
        .A(DP_mult_204_n376), .ZN(DP_mult_204_n372) );
  NAND2_X1 DP_mult_204_U2646 ( .A1(DP_mult_204_n382), .A2(DP_mult_204_n2234), 
        .ZN(DP_mult_204_n371) );
  INV_X1 DP_mult_204_U2645 ( .A(DP_mult_204_n346), .ZN(DP_mult_204_n344) );
  NAND2_X1 DP_mult_204_U2644 ( .A1(DP_mult_204_n2234), .A2(DP_mult_204_n378), 
        .ZN(DP_mult_204_n305) );
  INV_X1 DP_mult_204_U2643 ( .A(DP_coeffs_fb_int[4]), .ZN(DP_mult_204_n2375)
         );
  NAND2_X1 DP_mult_204_U2642 ( .A1(DP_mult_204_n2065), .A2(DP_mult_204_n489), 
        .ZN(DP_mult_204_n452) );
  OAI21_X1 DP_mult_204_U2641 ( .B1(DP_mult_204_n506), .B2(DP_mult_204_n452), 
        .A(DP_mult_204_n453), .ZN(DP_mult_204_n451) );
  NAND2_X1 DP_mult_204_U2640 ( .A1(DP_mult_204_n1808), .A2(DP_mult_204_n1958), 
        .ZN(DP_mult_204_n293) );
  OAI22_X1 DP_mult_204_U2639 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1541), 
        .B1(DP_mult_204_n1540), .B2(DP_mult_204_n2327), .ZN(DP_mult_204_n1250)
         );
  OAI22_X1 DP_mult_204_U2638 ( .A1(DP_mult_204_n1556), .A2(DP_mult_204_n2327), 
        .B1(DP_mult_204_n2302), .B2(DP_mult_204_n1938), .ZN(DP_mult_204_n1184)
         );
  OAI22_X1 DP_mult_204_U2637 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1539), 
        .B1(DP_mult_204_n1538), .B2(DP_mult_204_n2326), .ZN(DP_mult_204_n1248)
         );
  OAI22_X1 DP_mult_204_U2636 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1533), 
        .B1(DP_mult_204_n1532), .B2(DP_mult_204_n2327), .ZN(DP_mult_204_n692)
         );
  OAI22_X1 DP_mult_204_U2635 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1543), 
        .B1(DP_mult_204_n1542), .B2(DP_mult_204_n2326), .ZN(DP_mult_204_n1252)
         );
  OAI22_X1 DP_mult_204_U2634 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1537), 
        .B1(DP_mult_204_n1536), .B2(DP_mult_204_n2327), .ZN(DP_mult_204_n1246)
         );
  OAI22_X1 DP_mult_204_U2633 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1535), 
        .B1(DP_mult_204_n1534), .B2(DP_mult_204_n2326), .ZN(DP_mult_204_n1244)
         );
  OAI21_X1 DP_mult_204_U2632 ( .B1(DP_mult_204_n2272), .B2(DP_mult_204_n550), 
        .A(DP_mult_204_n543), .ZN(DP_mult_204_n541) );
  OAI22_X1 DP_mult_204_U2631 ( .A1(DP_mult_204_n2185), .A2(DP_mult_204_n1697), 
        .B1(DP_mult_204_n1696), .B2(DP_mult_204_n2337), .ZN(DP_mult_204_n1400)
         );
  OAI22_X1 DP_mult_204_U2630 ( .A1(DP_mult_204_n2314), .A2(DP_mult_204_n1703), 
        .B1(DP_mult_204_n1702), .B2(DP_mult_204_n2337), .ZN(DP_mult_204_n1406)
         );
  OAI22_X1 DP_mult_204_U2629 ( .A1(DP_mult_204_n2314), .A2(DP_mult_204_n1699), 
        .B1(DP_mult_204_n1698), .B2(DP_mult_204_n2338), .ZN(DP_mult_204_n1402)
         );
  OAI22_X1 DP_mult_204_U2628 ( .A1(DP_mult_204_n2185), .A2(DP_mult_204_n1705), 
        .B1(DP_mult_204_n1704), .B2(DP_mult_204_n2337), .ZN(DP_mult_204_n1408)
         );
  OAI22_X1 DP_mult_204_U2627 ( .A1(DP_mult_204_n2185), .A2(DP_mult_204_n1700), 
        .B1(DP_mult_204_n2337), .B2(DP_mult_204_n1699), .ZN(DP_mult_204_n1403)
         );
  OAI22_X1 DP_mult_204_U2626 ( .A1(DP_mult_204_n2314), .A2(DP_mult_204_n1694), 
        .B1(DP_mult_204_n2337), .B2(DP_mult_204_n1693), .ZN(DP_mult_204_n1397)
         );
  OAI22_X1 DP_mult_204_U2625 ( .A1(DP_mult_204_n2186), .A2(DP_mult_204_n1698), 
        .B1(DP_mult_204_n2338), .B2(DP_mult_204_n1697), .ZN(DP_mult_204_n1401)
         );
  OAI22_X1 DP_mult_204_U2624 ( .A1(DP_mult_204_n2314), .A2(DP_mult_204_n1702), 
        .B1(DP_mult_204_n2337), .B2(DP_mult_204_n1701), .ZN(DP_mult_204_n1405)
         );
  OAI22_X1 DP_mult_204_U2623 ( .A1(DP_mult_204_n2185), .A2(DP_mult_204_n1696), 
        .B1(DP_mult_204_n2337), .B2(DP_mult_204_n1695), .ZN(DP_mult_204_n1399)
         );
  OAI22_X1 DP_mult_204_U2622 ( .A1(DP_mult_204_n2186), .A2(DP_mult_204_n1701), 
        .B1(DP_mult_204_n1700), .B2(DP_mult_204_n2337), .ZN(DP_mult_204_n1404)
         );
  OAI22_X1 DP_mult_204_U2621 ( .A1(DP_mult_204_n2186), .A2(DP_mult_204_n1704), 
        .B1(DP_mult_204_n2338), .B2(DP_mult_204_n1703), .ZN(DP_mult_204_n1407)
         );
  OAI22_X1 DP_mult_204_U2620 ( .A1(DP_mult_204_n2185), .A2(DP_mult_204_n1695), 
        .B1(DP_mult_204_n1694), .B2(DP_mult_204_n2337), .ZN(DP_mult_204_n1398)
         );
  OAI22_X1 DP_mult_204_U2619 ( .A1(DP_mult_204_n2315), .A2(DP_mult_204_n1712), 
        .B1(DP_mult_204_n1711), .B2(DP_mult_204_n2340), .ZN(DP_mult_204_n1414)
         );
  OAI22_X1 DP_mult_204_U2618 ( .A1(DP_mult_204_n1714), .A2(DP_mult_204_n2177), 
        .B1(DP_mult_204_n1713), .B2(DP_mult_204_n2341), .ZN(DP_mult_204_n1416)
         );
  OAI22_X1 DP_mult_204_U2617 ( .A1(DP_mult_204_n1710), .A2(DP_mult_204_n2177), 
        .B1(DP_mult_204_n1709), .B2(DP_mult_204_n2340), .ZN(DP_mult_204_n1412)
         );
  OAI22_X1 DP_mult_204_U2616 ( .A1(DP_mult_204_n2177), .A2(DP_mult_204_n1715), 
        .B1(DP_mult_204_n2341), .B2(DP_mult_204_n1714), .ZN(DP_mult_204_n1417)
         );
  OAI22_X1 DP_mult_204_U2615 ( .A1(DP_mult_204_n2315), .A2(DP_mult_204_n1709), 
        .B1(DP_mult_204_n2340), .B2(DP_mult_204_n1708), .ZN(DP_mult_204_n1411)
         );
  OAI22_X1 DP_mult_204_U2614 ( .A1(DP_mult_204_n2315), .A2(DP_mult_204_n1708), 
        .B1(DP_mult_204_n1707), .B2(DP_mult_204_n2341), .ZN(DP_mult_204_n874)
         );
  OAI22_X1 DP_mult_204_U2613 ( .A1(DP_mult_204_n2177), .A2(DP_mult_204_n1711), 
        .B1(DP_mult_204_n2340), .B2(DP_mult_204_n1710), .ZN(DP_mult_204_n1413)
         );
  OAI22_X1 DP_mult_204_U2612 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1716), 
        .B1(DP_mult_204_n1715), .B2(DP_mult_204_n2341), .ZN(DP_mult_204_n1418)
         );
  OAI22_X1 DP_mult_204_U2611 ( .A1(DP_mult_204_n2316), .A2(DP_mult_204_n1713), 
        .B1(DP_mult_204_n2340), .B2(DP_mult_204_n1712), .ZN(DP_mult_204_n1415)
         );
  OAI22_X1 DP_mult_204_U2610 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1717), 
        .B1(DP_mult_204_n2341), .B2(DP_mult_204_n1716), .ZN(DP_mult_204_n1419)
         );
  OAI22_X1 DP_mult_204_U2609 ( .A1(DP_mult_204_n1731), .A2(DP_mult_204_n2341), 
        .B1(DP_mult_204_n2316), .B2(DP_mult_204_n1975), .ZN(DP_mult_204_n1191)
         );
  OAI22_X1 DP_mult_204_U2608 ( .A1(DP_mult_204_n2178), .A2(DP_mult_204_n1718), 
        .B1(DP_mult_204_n1717), .B2(DP_mult_204_n2341), .ZN(DP_mult_204_n1420)
         );
  NAND2_X1 DP_mult_204_U2607 ( .A1(DP_mult_204_n1811), .A2(DP_mult_204_n2061), 
        .ZN(DP_mult_204_n287) );
  OAI22_X1 DP_mult_204_U2606 ( .A1(DP_mult_204_n2308), .A2(DP_mult_204_n1616), 
        .B1(DP_mult_204_n1615), .B2(DP_mult_204_n2333), .ZN(DP_mult_204_n1322)
         );
  OAI22_X1 DP_mult_204_U2605 ( .A1(DP_mult_204_n2070), .A2(DP_mult_204_n1608), 
        .B1(DP_mult_204_n1607), .B2(DP_mult_204_n1969), .ZN(DP_mult_204_n746)
         );
  OAI22_X1 DP_mult_204_U2604 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1618), 
        .B1(DP_mult_204_n1617), .B2(DP_mult_204_n2333), .ZN(DP_mult_204_n1324)
         );
  OAI22_X1 DP_mult_204_U2603 ( .A1(DP_mult_204_n2308), .A2(DP_mult_204_n1614), 
        .B1(DP_mult_204_n1613), .B2(DP_mult_204_n1970), .ZN(DP_mult_204_n1320)
         );
  OAI22_X1 DP_mult_204_U2602 ( .A1(DP_mult_204_n1631), .A2(DP_mult_204_n1970), 
        .B1(DP_mult_204_n2257), .B2(DP_mult_204_n1931), .ZN(DP_mult_204_n1187)
         );
  OAI22_X1 DP_mult_204_U2601 ( .A1(DP_mult_204_n1967), .A2(DP_mult_204_n1610), 
        .B1(DP_mult_204_n1609), .B2(DP_mult_204_n1970), .ZN(DP_mult_204_n1316)
         );
  OAI22_X1 DP_mult_204_U2600 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1612), 
        .B1(DP_mult_204_n1611), .B2(DP_mult_204_n2333), .ZN(DP_mult_204_n1318)
         );
  AOI21_X1 DP_mult_204_U2599 ( .B1(DP_mult_204_n589), .B2(DP_mult_204_n2227), 
        .A(DP_mult_204_n2224), .ZN(DP_mult_204_n583) );
  NAND2_X1 DP_mult_204_U2598 ( .A1(DP_mult_204_n588), .A2(DP_mult_204_n2227), 
        .ZN(DP_mult_204_n582) );
  OAI22_X1 DP_mult_204_U2597 ( .A1(DP_mult_204_n2298), .A2(DP_mult_204_n1504), 
        .B1(DP_mult_204_n2321), .B2(DP_mult_204_n1503), .ZN(DP_mult_204_n1215)
         );
  OAI22_X1 DP_mult_204_U2596 ( .A1(DP_mult_204_n2289), .A2(DP_mult_204_n1503), 
        .B1(DP_mult_204_n1502), .B2(DP_mult_204_n2321), .ZN(DP_mult_204_n1214)
         );
  OAI22_X1 DP_mult_204_U2595 ( .A1(DP_mult_204_n2289), .A2(DP_mult_204_n1498), 
        .B1(DP_mult_204_n2322), .B2(DP_mult_204_n1497), .ZN(DP_mult_204_n1209)
         );
  OAI22_X1 DP_mult_204_U2594 ( .A1(DP_mult_204_n2289), .A2(DP_mult_204_n1499), 
        .B1(DP_mult_204_n1498), .B2(DP_mult_204_n2322), .ZN(DP_mult_204_n1210)
         );
  OAI22_X1 DP_mult_204_U2593 ( .A1(DP_mult_204_n2298), .A2(DP_mult_204_n1501), 
        .B1(DP_mult_204_n1500), .B2(DP_mult_204_n2322), .ZN(DP_mult_204_n1212)
         );
  OAI22_X1 DP_mult_204_U2592 ( .A1(DP_mult_204_n2298), .A2(DP_mult_204_n1502), 
        .B1(DP_mult_204_n2321), .B2(DP_mult_204_n1501), .ZN(DP_mult_204_n1213)
         );
  OAI22_X1 DP_mult_204_U2591 ( .A1(DP_mult_204_n2298), .A2(DP_mult_204_n1500), 
        .B1(DP_mult_204_n2321), .B2(DP_mult_204_n1499), .ZN(DP_mult_204_n1211)
         );
  OAI22_X1 DP_mult_204_U2590 ( .A1(DP_mult_204_n2255), .A2(DP_mult_204_n1494), 
        .B1(DP_mult_204_n2322), .B2(DP_mult_204_n1493), .ZN(DP_mult_204_n1205)
         );
  OAI22_X1 DP_mult_204_U2589 ( .A1(DP_mult_204_n2289), .A2(DP_mult_204_n1495), 
        .B1(DP_mult_204_n1494), .B2(DP_mult_204_n2321), .ZN(DP_mult_204_n1206)
         );
  OR2_X1 DP_mult_204_U2588 ( .A1(DP_mult_204_n1215), .A2(DP_mult_204_n1237), 
        .ZN(DP_mult_204_n938) );
  OAI22_X1 DP_mult_204_U2587 ( .A1(DP_mult_204_n2255), .A2(DP_mult_204_n1496), 
        .B1(DP_mult_204_n2322), .B2(DP_mult_204_n1495), .ZN(DP_mult_204_n1207)
         );
  XNOR2_X1 DP_mult_204_U2586 ( .A(DP_mult_204_n1237), .B(DP_mult_204_n2253), 
        .ZN(DP_mult_204_n939) );
  OAI22_X1 DP_mult_204_U2585 ( .A1(DP_mult_204_n2254), .A2(DP_mult_204_n1497), 
        .B1(DP_mult_204_n1496), .B2(DP_mult_204_n2322), .ZN(DP_mult_204_n1208)
         );
  AOI21_X1 DP_mult_204_U2584 ( .B1(DP_mult_204_n1932), .B2(DP_mult_204_n553), 
        .A(DP_mult_204_n541), .ZN(DP_mult_204_n539) );
  OAI22_X1 DP_mult_204_U2583 ( .A1(DP_mult_204_n2140), .A2(DP_mult_204_n1655), 
        .B1(DP_mult_204_n1654), .B2(DP_mult_204_n2118), .ZN(DP_mult_204_n1360)
         );
  XNOR2_X1 DP_mult_204_U2582 ( .A(DP_mult_204_n475), .B(DP_mult_204_n314), 
        .ZN(DP_sw0_coeff_ret0[10]) );
  INV_X1 DP_mult_204_U2581 ( .A(DP_coeffs_fb_int[22]), .ZN(DP_mult_204_n2347)
         );
  OAI21_X1 DP_mult_204_U2580 ( .B1(DP_mult_204_n631), .B2(DP_mult_204_n634), 
        .A(DP_mult_204_n632), .ZN(DP_mult_204_n630) );
  OAI21_X1 DP_mult_204_U2579 ( .B1(DP_mult_204_n638), .B2(DP_mult_204_n636), 
        .A(DP_mult_204_n637), .ZN(DP_mult_204_n635) );
  NAND2_X1 DP_mult_204_U2578 ( .A1(DP_mult_204_n1812), .A2(DP_mult_204_n2181), 
        .ZN(DP_mult_204_n285) );
  OAI22_X1 DP_mult_204_U2577 ( .A1(DP_mult_204_n2141), .A2(DP_mult_204_n1653), 
        .B1(DP_mult_204_n1652), .B2(DP_mult_204_n2042), .ZN(DP_mult_204_n1358)
         );
  OAI21_X1 DP_mult_204_U2576 ( .B1(DP_mult_204_n558), .B2(DP_mult_204_n564), 
        .A(DP_mult_204_n559), .ZN(DP_mult_204_n553) );
  NAND2_X1 DP_mult_204_U2575 ( .A1(DP_mult_204_n540), .A2(DP_mult_204_n552), 
        .ZN(DP_mult_204_n538) );
  INV_X1 DP_mult_204_U2574 ( .A(DP_mult_204_n552), .ZN(DP_mult_204_n554) );
  AOI21_X1 DP_mult_204_U2573 ( .B1(DP_mult_204_n565), .B2(DP_mult_204_n2002), 
        .A(DP_mult_204_n2249), .ZN(DP_mult_204_n551) );
  NAND2_X1 DP_mult_204_U2572 ( .A1(DP_mult_204_n1807), .A2(DP_mult_204_n2323), 
        .ZN(DP_mult_204_n295) );
  OAI22_X1 DP_mult_204_U2571 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1516), 
        .B1(DP_mult_204_n1515), .B2(DP_mult_204_n2324), .ZN(DP_mult_204_n1226)
         );
  OAI22_X1 DP_mult_204_U2570 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1517), 
        .B1(DP_mult_204_n2324), .B2(DP_mult_204_n1516), .ZN(DP_mult_204_n1227)
         );
  OAI22_X1 DP_mult_204_U2569 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1512), 
        .B1(DP_mult_204_n1511), .B2(DP_mult_204_n2325), .ZN(DP_mult_204_n1222)
         );
  OAI22_X1 DP_mult_204_U2568 ( .A1(DP_mult_204_n1531), .A2(DP_mult_204_n2325), 
        .B1(DP_mult_204_n2180), .B2(DP_mult_204_n2034), .ZN(DP_mult_204_n1183)
         );
  OAI22_X1 DP_mult_204_U2567 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1515), 
        .B1(DP_mult_204_n2325), .B2(DP_mult_204_n1514), .ZN(DP_mult_204_n1225)
         );
  OAI22_X1 DP_mult_204_U2566 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1509), 
        .B1(DP_mult_204_n2325), .B2(DP_mult_204_n1508), .ZN(DP_mult_204_n1219)
         );
  OAI22_X1 DP_mult_204_U2565 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1510), 
        .B1(DP_mult_204_n1509), .B2(DP_mult_204_n2324), .ZN(DP_mult_204_n1220)
         );
  OAI22_X1 DP_mult_204_U2564 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1514), 
        .B1(DP_mult_204_n1513), .B2(DP_mult_204_n2324), .ZN(DP_mult_204_n1224)
         );
  OAI22_X1 DP_mult_204_U2563 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1511), 
        .B1(DP_mult_204_n2324), .B2(DP_mult_204_n1510), .ZN(DP_mult_204_n1221)
         );
  OAI22_X1 DP_mult_204_U2562 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1518), 
        .B1(DP_mult_204_n1517), .B2(DP_mult_204_n2324), .ZN(DP_mult_204_n1228)
         );
  OAI22_X1 DP_mult_204_U2561 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1513), 
        .B1(DP_mult_204_n2325), .B2(DP_mult_204_n1512), .ZN(DP_mult_204_n1223)
         );
  OAI22_X1 DP_mult_204_U2560 ( .A1(DP_mult_204_n2180), .A2(DP_mult_204_n1508), 
        .B1(DP_mult_204_n1507), .B2(DP_mult_204_n2324), .ZN(DP_mult_204_n682)
         );
  AOI21_X1 DP_mult_204_U2559 ( .B1(DP_mult_204_n401), .B2(DP_mult_204_n2230), 
        .A(DP_mult_204_n394), .ZN(DP_mult_204_n390) );
  OAI21_X1 DP_mult_204_U2558 ( .B1(DP_mult_204_n390), .B2(DP_mult_204_n384), 
        .A(DP_mult_204_n387), .ZN(DP_mult_204_n383) );
  INV_X1 DP_mult_204_U2557 ( .A(DP_mult_204_n401), .ZN(DP_mult_204_n399) );
  NAND2_X1 DP_mult_204_U2556 ( .A1(DP_mult_204_n877), .A2(DP_mult_204_n896), 
        .ZN(DP_mult_204_n532) );
  INV_X1 DP_mult_204_U2555 ( .A(DP_mult_204_n2288), .ZN(DP_mult_204_n508) );
  INV_X1 DP_mult_204_U2554 ( .A(DP_coeffs_fb_int[20]), .ZN(DP_mult_204_n2349)
         );
  OAI21_X1 DP_mult_204_U2553 ( .B1(DP_mult_204_n495), .B2(DP_mult_204_n503), 
        .A(DP_mult_204_n496), .ZN(DP_mult_204_n490) );
  OAI21_X1 DP_mult_204_U2552 ( .B1(DP_mult_204_n492), .B2(DP_mult_204_n467), 
        .A(DP_mult_204_n468), .ZN(DP_mult_204_n466) );
  OAI21_X1 DP_mult_204_U2551 ( .B1(DP_mult_204_n492), .B2(DP_mult_204_n480), 
        .A(DP_mult_204_n481), .ZN(DP_mult_204_n479) );
  OAI22_X1 DP_mult_204_U2550 ( .A1(DP_mult_204_n1977), .A2(DP_mult_204_n1591), 
        .B1(DP_mult_204_n1590), .B2(DP_mult_204_n2332), .ZN(DP_mult_204_n1298)
         );
  OAI22_X1 DP_mult_204_U2549 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1587), 
        .B1(DP_mult_204_n1586), .B2(DP_mult_204_n2331), .ZN(DP_mult_204_n1294)
         );
  OAI22_X1 DP_mult_204_U2548 ( .A1(DP_mult_204_n1606), .A2(DP_mult_204_n2331), 
        .B1(DP_mult_204_n2307), .B2(DP_mult_204_n2045), .ZN(DP_mult_204_n1186)
         );
  OAI22_X1 DP_mult_204_U2547 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1585), 
        .B1(DP_mult_204_n1584), .B2(DP_mult_204_n2332), .ZN(DP_mult_204_n1292)
         );
  OAI22_X1 DP_mult_204_U2546 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1583), 
        .B1(DP_mult_204_n1582), .B2(DP_mult_204_n2332), .ZN(DP_mult_204_n724)
         );
  OAI22_X1 DP_mult_204_U2545 ( .A1(DP_mult_204_n2306), .A2(DP_mult_204_n1589), 
        .B1(DP_mult_204_n1588), .B2(DP_mult_204_n2331), .ZN(DP_mult_204_n1296)
         );
  OAI22_X1 DP_mult_204_U2544 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1593), 
        .B1(DP_mult_204_n1592), .B2(DP_mult_204_n2332), .ZN(DP_mult_204_n1300)
         );
  AOI21_X1 DP_mult_204_U2543 ( .B1(DP_mult_204_n508), .B2(DP_mult_204_n465), 
        .A(DP_mult_204_n466), .ZN(DP_mult_204_n464) );
  AOI21_X1 DP_mult_204_U2542 ( .B1(DP_mult_204_n508), .B2(DP_mult_204_n668), 
        .A(DP_mult_204_n2149), .ZN(DP_mult_204_n499) );
  AOI21_X1 DP_mult_204_U2541 ( .B1(DP_mult_204_n508), .B2(DP_mult_204_n478), 
        .A(DP_mult_204_n479), .ZN(DP_mult_204_n477) );
  XNOR2_X1 DP_mult_204_U2540 ( .A(DP_mult_204_n462), .B(DP_mult_204_n313), 
        .ZN(DP_sw0_coeff_ret0[11]) );
  NAND2_X1 DP_mult_204_U2539 ( .A1(DP_mult_204_n839), .A2(DP_mult_204_n856), 
        .ZN(DP_mult_204_n514) );
  OAI21_X1 DP_mult_204_U2538 ( .B1(DP_mult_204_n2169), .B2(DP_mult_204_n2015), 
        .A(DP_mult_204_n2387), .ZN(DP_mult_204_n1386) );
  INV_X1 DP_mult_204_U2537 ( .A(DP_mult_204_n474), .ZN(DP_mult_204_n472) );
  NAND2_X1 DP_mult_204_U2536 ( .A1(DP_mult_204_n2225), .A2(DP_mult_204_n474), 
        .ZN(DP_mult_204_n314) );
  NOR2_X1 DP_mult_204_U2535 ( .A1(DP_mult_204_n534), .A2(DP_mult_204_n531), 
        .ZN(DP_mult_204_n525) );
  NAND2_X1 DP_mult_204_U2534 ( .A1(DP_mult_204_n525), .A2(DP_mult_204_n1933), 
        .ZN(DP_mult_204_n505) );
  INV_X1 DP_mult_204_U2533 ( .A(DP_mult_204_n534), .ZN(DP_mult_204_n672) );
  NAND2_X1 DP_mult_204_U2532 ( .A1(DP_mult_204_n525), .A2(DP_mult_204_n670), 
        .ZN(DP_mult_204_n516) );
  INV_X1 DP_mult_204_U2531 ( .A(DP_mult_204_n382), .ZN(DP_mult_204_n380) );
  INV_X1 DP_mult_204_U2530 ( .A(DP_mult_204_n746), .ZN(DP_mult_204_n747) );
  NAND2_X1 DP_mult_204_U2529 ( .A1(DP_mult_204_n709), .A2(DP_mult_204_n716), 
        .ZN(DP_mult_204_n409) );
  OAI21_X1 DP_mult_204_U2528 ( .B1(DP_mult_204_n421), .B2(DP_mult_204_n402), 
        .A(DP_mult_204_n405), .ZN(DP_mult_204_n401) );
  INV_X1 DP_mult_204_U2527 ( .A(DP_mult_204_n874), .ZN(DP_mult_204_n875) );
  NAND2_X1 DP_mult_204_U2526 ( .A1(DP_mult_204_n2007), .A2(DP_mult_204_n2225), 
        .ZN(DP_mult_204_n467) );
  AOI21_X1 DP_mult_204_U2525 ( .B1(DP_mult_204_n2225), .B2(DP_mult_204_n483), 
        .A(DP_mult_204_n472), .ZN(DP_mult_204_n468) );
  NAND2_X1 DP_mult_204_U2524 ( .A1(DP_mult_204_n807), .A2(DP_mult_204_n822), 
        .ZN(DP_mult_204_n2297) );
  NAND2_X1 DP_mult_204_U2523 ( .A1(DP_mult_204_n809), .A2(DP_mult_204_n2006), 
        .ZN(DP_mult_204_n2296) );
  NAND2_X1 DP_mult_204_U2522 ( .A1(DP_mult_204_n809), .A2(DP_mult_204_n807), 
        .ZN(DP_mult_204_n2295) );
  NAND3_X1 DP_mult_204_U2521 ( .A1(DP_mult_204_n2292), .A2(DP_mult_204_n2293), 
        .A3(DP_mult_204_n2294), .ZN(DP_mult_204_n822) );
  NAND2_X1 DP_mult_204_U2520 ( .A1(DP_mult_204_n844), .A2(DP_mult_204_n842), 
        .ZN(DP_mult_204_n2294) );
  NAND2_X1 DP_mult_204_U2519 ( .A1(DP_mult_204_n827), .A2(DP_mult_204_n2127), 
        .ZN(DP_mult_204_n2293) );
  NAND2_X1 DP_mult_204_U2518 ( .A1(DP_mult_204_n827), .A2(DP_mult_204_n844), 
        .ZN(DP_mult_204_n2292) );
  OAI22_X1 DP_mult_204_U2517 ( .A1(DP_mult_204_n2318), .A2(DP_mult_204_n1751), 
        .B1(DP_mult_204_n1750), .B2(DP_mult_204_n2342), .ZN(DP_mult_204_n1452)
         );
  OAI22_X1 DP_mult_204_U2516 ( .A1(DP_mult_204_n2279), .A2(DP_mult_204_n1752), 
        .B1(DP_mult_204_n2342), .B2(DP_mult_204_n1751), .ZN(DP_mult_204_n1453)
         );
  OAI22_X1 DP_mult_204_U2515 ( .A1(DP_mult_204_n2318), .A2(DP_mult_204_n1746), 
        .B1(DP_mult_204_n1978), .B2(DP_mult_204_n1745), .ZN(DP_mult_204_n1447)
         );
  OAI22_X1 DP_mult_204_U2514 ( .A1(DP_mult_204_n2318), .A2(DP_mult_204_n1748), 
        .B1(DP_mult_204_n2342), .B2(DP_mult_204_n1747), .ZN(DP_mult_204_n1449)
         );
  OAI22_X1 DP_mult_204_U2513 ( .A1(DP_mult_204_n2318), .A2(DP_mult_204_n1749), 
        .B1(DP_mult_204_n1748), .B2(DP_mult_204_n2342), .ZN(DP_mult_204_n1450)
         );
  OAI22_X1 DP_mult_204_U2512 ( .A1(DP_mult_204_n2278), .A2(DP_mult_204_n1744), 
        .B1(DP_mult_204_n1978), .B2(DP_mult_204_n1743), .ZN(DP_mult_204_n1445)
         );
  OAI22_X1 DP_mult_204_U2511 ( .A1(DP_mult_204_n2279), .A2(DP_mult_204_n1754), 
        .B1(DP_mult_204_n2342), .B2(DP_mult_204_n1753), .ZN(DP_mult_204_n1455)
         );
  OAI22_X1 DP_mult_204_U2510 ( .A1(DP_mult_204_n2278), .A2(DP_mult_204_n1750), 
        .B1(DP_mult_204_n2342), .B2(DP_mult_204_n1749), .ZN(DP_mult_204_n1451)
         );
  OAI22_X1 DP_mult_204_U2509 ( .A1(DP_mult_204_n2318), .A2(DP_mult_204_n1747), 
        .B1(DP_mult_204_n1746), .B2(DP_mult_204_n2342), .ZN(DP_mult_204_n1448)
         );
  OAI22_X1 DP_mult_204_U2508 ( .A1(DP_mult_204_n2279), .A2(DP_mult_204_n1745), 
        .B1(DP_mult_204_n1744), .B2(DP_mult_204_n2342), .ZN(DP_mult_204_n1446)
         );
  NAND2_X1 DP_mult_204_U2507 ( .A1(DP_mult_204_n1165), .A2(DP_mult_204_n1170), 
        .ZN(DP_mult_204_n632) );
  OAI21_X1 DP_mult_204_U2506 ( .B1(DP_mult_204_n513), .B2(DP_mult_204_n521), 
        .A(DP_mult_204_n514), .ZN(DP_mult_204_n512) );
  OAI22_X1 DP_mult_204_U2505 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1676), 
        .B1(DP_mult_204_n1675), .B2(DP_mult_204_n2335), .ZN(DP_mult_204_n1380)
         );
  OAI22_X1 DP_mult_204_U2504 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1674), 
        .B1(DP_mult_204_n1673), .B2(DP_mult_204_n2335), .ZN(DP_mult_204_n1378)
         );
  OAI22_X1 DP_mult_204_U2503 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1679), 
        .B1(DP_mult_204_n2069), .B2(DP_mult_204_n1678), .ZN(DP_mult_204_n1383)
         );
  OAI22_X1 DP_mult_204_U2502 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1677), 
        .B1(DP_mult_204_n2069), .B2(DP_mult_204_n1676), .ZN(DP_mult_204_n1381)
         );
  OAI22_X1 DP_mult_204_U2501 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1673), 
        .B1(DP_mult_204_n2335), .B2(DP_mult_204_n1672), .ZN(DP_mult_204_n1377)
         );
  OAI22_X1 DP_mult_204_U2500 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1675), 
        .B1(DP_mult_204_n2335), .B2(DP_mult_204_n1674), .ZN(DP_mult_204_n1379)
         );
  OAI22_X1 DP_mult_204_U2499 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1672), 
        .B1(DP_mult_204_n1671), .B2(DP_mult_204_n2335), .ZN(DP_mult_204_n1376)
         );
  OAI22_X1 DP_mult_204_U2498 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1669), 
        .B1(DP_mult_204_n2335), .B2(DP_mult_204_n1668), .ZN(DP_mult_204_n1373)
         );
  OAI22_X1 DP_mult_204_U2497 ( .A1(DP_mult_204_n2311), .A2(DP_mult_204_n1670), 
        .B1(DP_mult_204_n1669), .B2(DP_mult_204_n2335), .ZN(DP_mult_204_n1374)
         );
  OAI22_X1 DP_mult_204_U2496 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1671), 
        .B1(DP_mult_204_n2069), .B2(DP_mult_204_n1670), .ZN(DP_mult_204_n1375)
         );
  AOI21_X1 DP_mult_204_U2495 ( .B1(DP_mult_204_n2126), .B2(DP_mult_204_n670), 
        .A(DP_mult_204_n519), .ZN(DP_mult_204_n517) );
  INV_X1 DP_mult_204_U2494 ( .A(DP_mult_204_n2277), .ZN(DP_mult_204_n524) );
  XNOR2_X1 DP_mult_204_U2493 ( .A(DP_sw0_11_), .B(DP_mult_204_n2367), .ZN(
        DP_mult_204_n1594) );
  XNOR2_X1 DP_mult_204_U2492 ( .A(DP_sw0_19_), .B(DP_mult_204_n2367), .ZN(
        DP_mult_204_n1586) );
  XNOR2_X1 DP_mult_204_U2491 ( .A(DP_sw0_13_), .B(DP_mult_204_n2366), .ZN(
        DP_mult_204_n1592) );
  XNOR2_X1 DP_mult_204_U2490 ( .A(DP_sw0_15_), .B(DP_mult_204_n2366), .ZN(
        DP_mult_204_n1590) );
  XNOR2_X1 DP_mult_204_U2489 ( .A(DP_sw0_17_), .B(DP_mult_204_n2367), .ZN(
        DP_mult_204_n1588) );
  XNOR2_X1 DP_mult_204_U2488 ( .A(DP_sw0_21_), .B(DP_mult_204_n2367), .ZN(
        DP_mult_204_n1584) );
  INV_X1 DP_mult_204_U2487 ( .A(DP_mult_204_n706), .ZN(DP_mult_204_n707) );
  NAND2_X1 DP_mult_204_U2486 ( .A1(DP_mult_204_n685), .A2(DP_mult_204_n688), 
        .ZN(DP_mult_204_n369) );
  AOI21_X1 DP_mult_204_U2485 ( .B1(DP_mult_204_n359), .B2(DP_mult_204_n2238), 
        .A(DP_mult_204_n350), .ZN(DP_mult_204_n348) );
  AOI21_X1 DP_mult_204_U2484 ( .B1(DP_mult_204_n423), .B2(DP_mult_204_n356), 
        .A(DP_mult_204_n359), .ZN(DP_mult_204_n355) );
  OAI21_X1 DP_mult_204_U2483 ( .B1(DP_mult_204_n337), .B2(DP_mult_204_n334), 
        .A(DP_mult_204_n335), .ZN(DP_mult_204_n333) );
  XNOR2_X1 DP_mult_204_U2482 ( .A(DP_sw0_13_), .B(DP_mult_204_n2370), .ZN(
        DP_mult_204_n1567) );
  XNOR2_X1 DP_mult_204_U2481 ( .A(DP_sw0_11_), .B(DP_mult_204_n2369), .ZN(
        DP_mult_204_n1569) );
  XNOR2_X1 DP_mult_204_U2480 ( .A(DP_sw0_19_), .B(DP_mult_204_n2369), .ZN(
        DP_mult_204_n1561) );
  XNOR2_X1 DP_mult_204_U2479 ( .A(DP_sw0_17_), .B(DP_mult_204_n2369), .ZN(
        DP_mult_204_n1563) );
  XNOR2_X1 DP_mult_204_U2478 ( .A(DP_sw0_15_), .B(DP_mult_204_n2370), .ZN(
        DP_mult_204_n1565) );
  XNOR2_X1 DP_mult_204_U2477 ( .A(DP_sw0_21_), .B(DP_mult_204_n2369), .ZN(
        DP_mult_204_n1559) );
  NOR2_X1 DP_mult_204_U2476 ( .A1(DP_mult_204_n2163), .A2(DP_mult_204_n520), 
        .ZN(DP_mult_204_n511) );
  INV_X1 DP_mult_204_U2475 ( .A(DP_mult_204_n520), .ZN(DP_mult_204_n670) );
  AOI21_X1 DP_mult_204_U2474 ( .B1(DP_mult_204_n2233), .B2(DP_mult_204_n1985), 
        .A(DP_mult_204_n1994), .ZN(DP_mult_204_n600) );
  NAND2_X1 DP_mult_204_U2473 ( .A1(DP_mult_204_n2233), .A2(DP_mult_204_n2236), 
        .ZN(DP_mult_204_n599) );
  OAI21_X1 DP_mult_204_U2472 ( .B1(DP_mult_204_n600), .B2(DP_mult_204_n597), 
        .A(DP_mult_204_n598), .ZN(DP_mult_204_n596) );
  OAI21_X1 DP_mult_204_U2471 ( .B1(DP_mult_204_n481), .B2(DP_mult_204_n1936), 
        .A(DP_mult_204_n457), .ZN(DP_mult_204_n455) );
  OAI22_X1 DP_mult_204_U2470 ( .A1(DP_mult_204_n2140), .A2(DP_mult_204_n1651), 
        .B1(DP_mult_204_n1650), .B2(DP_mult_204_n2334), .ZN(DP_mult_204_n1356)
         );
  AOI21_X1 DP_mult_204_U2469 ( .B1(DP_mult_204_n2228), .B2(DP_mult_204_n1990), 
        .A(DP_mult_204_n2223), .ZN(DP_mult_204_n572) );
  NAND2_X1 DP_mult_204_U2468 ( .A1(DP_mult_204_n1071), .A2(DP_mult_204_n1084), 
        .ZN(DP_mult_204_n591) );
  OAI21_X1 DP_mult_204_U2467 ( .B1(DP_mult_204_n594), .B2(DP_mult_204_n582), 
        .A(DP_mult_204_n583), .ZN(DP_mult_204_n581) );
  XNOR2_X1 DP_mult_204_U2466 ( .A(DP_sw0_7_), .B(DP_mult_204_n2344), .ZN(
        DP_mult_204_n1773) );
  XNOR2_X1 DP_mult_204_U2465 ( .A(DP_sw0_3_), .B(DP_mult_204_n2344), .ZN(
        DP_mult_204_n1777) );
  XNOR2_X1 DP_mult_204_U2464 ( .A(DP_sw0_5_), .B(DP_mult_204_n2344), .ZN(
        DP_mult_204_n1775) );
  XNOR2_X1 DP_mult_204_U2463 ( .A(DP_sw0_9_), .B(DP_mult_204_n2344), .ZN(
        DP_mult_204_n1771) );
  XNOR2_X1 DP_mult_204_U2462 ( .A(DP_sw0_23_), .B(DP_mult_204_n2344), .ZN(
        DP_mult_204_n1757) );
  XNOR2_X1 DP_mult_204_U2461 ( .A(DP_sw0_1_), .B(DP_mult_204_n2344), .ZN(
        DP_mult_204_n1779) );
  OAI22_X1 DP_mult_204_U2460 ( .A1(DP_mult_204_n2319), .A2(DP_mult_204_n1762), 
        .B1(DP_mult_204_n1761), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1463)
         );
  OAI22_X1 DP_mult_204_U2459 ( .A1(DP_mult_204_n2320), .A2(DP_mult_204_n1758), 
        .B1(DP_mult_204_n1757), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1459)
         );
  OAI22_X1 DP_mult_204_U2458 ( .A1(DP_mult_204_n2320), .A2(DP_mult_204_n1763), 
        .B1(DP_mult_204_n1762), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1464)
         );
  OAI22_X1 DP_mult_204_U2457 ( .A1(DP_mult_204_n2121), .A2(DP_mult_204_n1765), 
        .B1(DP_mult_204_n1764), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1466)
         );
  OAI22_X1 DP_mult_204_U2456 ( .A1(DP_mult_204_n2319), .A2(DP_mult_204_n1766), 
        .B1(DP_mult_204_n1765), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1467)
         );
  OAI22_X1 DP_mult_204_U2455 ( .A1(DP_mult_204_n2121), .A2(DP_mult_204_n1760), 
        .B1(DP_mult_204_n1759), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1461)
         );
  OAI22_X1 DP_mult_204_U2454 ( .A1(DP_mult_204_n2320), .A2(DP_mult_204_n1767), 
        .B1(DP_mult_204_n1766), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1468)
         );
  OAI22_X1 DP_mult_204_U2453 ( .A1(DP_mult_204_n2319), .A2(DP_mult_204_n1761), 
        .B1(DP_mult_204_n1760), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1462)
         );
  OAI22_X1 DP_mult_204_U2452 ( .A1(DP_mult_204_n2120), .A2(DP_mult_204_n1764), 
        .B1(DP_mult_204_n1763), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1465)
         );
  OAI22_X1 DP_mult_204_U2451 ( .A1(DP_mult_204_n2120), .A2(DP_mult_204_n1768), 
        .B1(DP_mult_204_n1767), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1469)
         );
  OAI22_X1 DP_mult_204_U2450 ( .A1(DP_mult_204_n1781), .A2(DP_mult_204_n251), 
        .B1(DP_mult_204_n2120), .B2(DP_mult_204_n2028), .ZN(DP_mult_204_n1193)
         );
  OAI22_X1 DP_mult_204_U2449 ( .A1(DP_mult_204_n2121), .A2(DP_mult_204_n1759), 
        .B1(DP_mult_204_n1758), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1460)
         );
  NAND2_X1 DP_mult_204_U2448 ( .A1(DP_mult_204_n941), .A2(DP_mult_204_n962), 
        .ZN(DP_mult_204_n550) );
  NOR2_X1 DP_mult_204_U2447 ( .A1(DP_mult_204_n542), .A2(DP_mult_204_n547), 
        .ZN(DP_mult_204_n540) );
  NOR2_X1 DP_mult_204_U2446 ( .A1(DP_mult_204_n554), .A2(DP_mult_204_n2156), 
        .ZN(DP_mult_204_n545) );
  OAI21_X1 DP_mult_204_U2445 ( .B1(DP_mult_204_n555), .B2(DP_mult_204_n2156), 
        .A(DP_mult_204_n550), .ZN(DP_mult_204_n546) );
  XNOR2_X1 DP_mult_204_U2444 ( .A(DP_mult_204_n2382), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1505) );
  INV_X1 DP_mult_204_U2443 ( .A(DP_mult_204_n297), .ZN(DP_mult_204_n2299) );
  NAND2_X1 DP_mult_204_U2442 ( .A1(DP_mult_204_n1806), .A2(DP_mult_204_n2011), 
        .ZN(DP_mult_204_n297) );
  AOI21_X1 DP_mult_204_U2441 ( .B1(DP_mult_204_n526), .B2(DP_mult_204_n511), 
        .A(DP_mult_204_n512), .ZN(DP_mult_204_n506) );
  NAND2_X1 DP_mult_204_U2440 ( .A1(DP_mult_204_n2290), .A2(DP_mult_204_n2291), 
        .ZN(DP_mult_204_n1216) );
  OR2_X1 DP_mult_204_U2439 ( .A1(DP_mult_204_n1504), .A2(DP_mult_204_n2322), 
        .ZN(DP_mult_204_n2291) );
  OR2_X1 DP_mult_204_U2438 ( .A1(DP_mult_204_n2289), .A2(DP_mult_204_n1505), 
        .ZN(DP_mult_204_n2290) );
  AOI21_X1 DP_mult_204_U2437 ( .B1(DP_mult_204_n2277), .B2(DP_mult_204_n2004), 
        .A(DP_mult_204_n2179), .ZN(DP_mult_204_n2288) );
  NOR2_X1 DP_mult_204_U2436 ( .A1(DP_mult_204_n456), .A2(DP_mult_204_n480), 
        .ZN(DP_mult_204_n454) );
  NOR2_X1 DP_mult_204_U2435 ( .A1(DP_mult_204_n2147), .A2(DP_mult_204_n480), 
        .ZN(DP_mult_204_n478) );
  NAND2_X1 DP_mult_204_U2434 ( .A1(DP_mult_204_n507), .A2(DP_mult_204_n489), 
        .ZN(DP_mult_204_n487) );
  NOR2_X1 DP_mult_204_U2433 ( .A1(DP_mult_204_n2287), .A2(DP_mult_204_n455), 
        .ZN(DP_mult_204_n453) );
  AND2_X1 DP_mult_204_U2432 ( .A1(DP_mult_204_n454), .A2(DP_mult_204_n490), 
        .ZN(DP_mult_204_n2287) );
  NAND3_X1 DP_mult_204_U2431 ( .A1(DP_mult_204_n2284), .A2(DP_mult_204_n2285), 
        .A3(DP_mult_204_n2286), .ZN(DP_mult_204_n812) );
  NAND2_X1 DP_mult_204_U2430 ( .A1(DP_mult_204_n830), .A2(DP_mult_204_n1386), 
        .ZN(DP_mult_204_n2286) );
  NAND2_X1 DP_mult_204_U2429 ( .A1(DP_mult_204_n834), .A2(DP_mult_204_n1386), 
        .ZN(DP_mult_204_n2285) );
  NAND2_X1 DP_mult_204_U2428 ( .A1(DP_mult_204_n830), .A2(DP_mult_204_n2043), 
        .ZN(DP_mult_204_n2284) );
  INV_X1 DP_mult_204_U2427 ( .A(DP_mult_204_n772), .ZN(DP_mult_204_n773) );
  NOR2_X1 DP_mult_204_U2426 ( .A1(DP_mult_204_n749), .A2(DP_mult_204_n760), 
        .ZN(DP_mult_204_n438) );
  NAND2_X1 DP_mult_204_U2425 ( .A1(DP_mult_204_n749), .A2(DP_mult_204_n760), 
        .ZN(DP_mult_204_n439) );
  NAND2_X1 DP_mult_204_U2424 ( .A1(DP_mult_204_n400), .A2(DP_mult_204_n2230), 
        .ZN(DP_mult_204_n389) );
  INV_X1 DP_mult_204_U2423 ( .A(DP_mult_204_n400), .ZN(DP_mult_204_n398) );
  INV_X1 DP_mult_204_U2422 ( .A(DP_mult_204_n2130), .ZN(DP_mult_204_n2317) );
  OAI22_X1 DP_mult_204_U2421 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1615), 
        .B1(DP_mult_204_n1969), .B2(DP_mult_204_n1614), .ZN(DP_mult_204_n1321)
         );
  OAI22_X1 DP_mult_204_U2420 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1611), 
        .B1(DP_mult_204_n1969), .B2(DP_mult_204_n1610), .ZN(DP_mult_204_n1317)
         );
  OAI22_X1 DP_mult_204_U2419 ( .A1(DP_mult_204_n1967), .A2(DP_mult_204_n1609), 
        .B1(DP_mult_204_n1970), .B2(DP_mult_204_n1608), .ZN(DP_mult_204_n1315)
         );
  OAI22_X1 DP_mult_204_U2418 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1617), 
        .B1(DP_mult_204_n1970), .B2(DP_mult_204_n1616), .ZN(DP_mult_204_n1323)
         );
  OAI22_X1 DP_mult_204_U2417 ( .A1(DP_mult_204_n2257), .A2(DP_mult_204_n1613), 
        .B1(DP_mult_204_n1970), .B2(DP_mult_204_n1612), .ZN(DP_mult_204_n1319)
         );
  NAND2_X1 DP_mult_204_U2416 ( .A1(DP_mult_204_n983), .A2(DP_mult_204_n1002), 
        .ZN(DP_mult_204_n564) );
  OAI22_X1 DP_mult_204_U2415 ( .A1(DP_mult_204_n2309), .A2(DP_mult_204_n1646), 
        .B1(DP_mult_204_n2334), .B2(DP_mult_204_n1645), .ZN(DP_mult_204_n1351)
         );
  NOR2_X1 DP_mult_204_U2414 ( .A1(DP_mult_204_n857), .A2(DP_mult_204_n876), 
        .ZN(DP_mult_204_n520) );
  OAI21_X1 DP_mult_204_U2413 ( .B1(DP_mult_204_n1973), .B2(DP_mult_204_n2145), 
        .A(DP_mult_204_n2389), .ZN(DP_mult_204_n1338) );
  OAI21_X1 DP_mult_204_U2412 ( .B1(DP_mult_204_n620), .B2(DP_mult_204_n610), 
        .A(DP_mult_204_n611), .ZN(DP_mult_204_n609) );
  NAND2_X1 DP_mult_204_U2411 ( .A1(DP_mult_204_n2225), .A2(DP_mult_204_n2226), 
        .ZN(DP_mult_204_n456) );
  NAND3_X1 DP_mult_204_U2410 ( .A1(DP_mult_204_n2281), .A2(DP_mult_204_n2282), 
        .A3(DP_mult_204_n2283), .ZN(DP_mult_204_n974) );
  NAND2_X1 DP_mult_204_U2409 ( .A1(DP_mult_204_n1974), .A2(DP_mult_204_n1393), 
        .ZN(DP_mult_204_n2283) );
  NAND2_X1 DP_mult_204_U2408 ( .A1(DP_mult_204_n1988), .A2(DP_mult_204_n1393), 
        .ZN(DP_mult_204_n2282) );
  NAND2_X1 DP_mult_204_U2407 ( .A1(DP_mult_204_n1974), .A2(DP_mult_204_n1988), 
        .ZN(DP_mult_204_n2281) );
  NOR2_X1 DP_mult_204_U2406 ( .A1(DP_mult_204_n1085), .A2(DP_mult_204_n1098), 
        .ZN(DP_mult_204_n592) );
  NAND2_X1 DP_mult_204_U2405 ( .A1(DP_mult_204_n1085), .A2(DP_mult_204_n1098), 
        .ZN(DP_mult_204_n593) );
  OAI22_X1 DP_mult_204_U2404 ( .A1(DP_mult_204_n2307), .A2(DP_mult_204_n1592), 
        .B1(DP_mult_204_n2332), .B2(DP_mult_204_n1591), .ZN(DP_mult_204_n1299)
         );
  OAI22_X1 DP_mult_204_U2403 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1586), 
        .B1(DP_mult_204_n2332), .B2(DP_mult_204_n1585), .ZN(DP_mult_204_n1293)
         );
  OAI22_X1 DP_mult_204_U2402 ( .A1(DP_mult_204_n2306), .A2(DP_mult_204_n1590), 
        .B1(DP_mult_204_n2332), .B2(DP_mult_204_n1589), .ZN(DP_mult_204_n1297)
         );
  OAI22_X1 DP_mult_204_U2401 ( .A1(DP_mult_204_n2306), .A2(DP_mult_204_n1588), 
        .B1(DP_mult_204_n2332), .B2(DP_mult_204_n1587), .ZN(DP_mult_204_n1295)
         );
  OAI22_X1 DP_mult_204_U2400 ( .A1(DP_mult_204_n2104), .A2(DP_mult_204_n1584), 
        .B1(DP_mult_204_n2331), .B2(DP_mult_204_n1583), .ZN(DP_mult_204_n1291)
         );
  XNOR2_X1 DP_mult_204_U2399 ( .A(DP_mult_204_n809), .B(DP_mult_204_n807), 
        .ZN(DP_mult_204_n2280) );
  XNOR2_X1 DP_mult_204_U2398 ( .A(DP_mult_204_n2280), .B(DP_mult_204_n822), 
        .ZN(DP_mult_204_n805) );
  OAI21_X1 DP_mult_204_U2397 ( .B1(DP_mult_204_n590), .B2(DP_mult_204_n593), 
        .A(DP_mult_204_n591), .ZN(DP_mult_204_n589) );
  NAND2_X1 DP_mult_204_U2396 ( .A1(DP_mult_204_n919), .A2(DP_mult_204_n940), 
        .ZN(DP_mult_204_n543) );
  INV_X1 DP_mult_204_U2395 ( .A(DP_mult_204_n505), .ZN(DP_mult_204_n507) );
  INV_X1 DP_mult_204_U2394 ( .A(DP_mult_204_n2129), .ZN(DP_mult_204_n2318) );
  INV_X1 DP_mult_204_U2393 ( .A(DP_mult_204_n2130), .ZN(DP_mult_204_n2278) );
  INV_X1 DP_mult_204_U2392 ( .A(DP_mult_204_n1987), .ZN(DP_mult_204_n2312) );
  OAI21_X1 DP_mult_204_U2391 ( .B1(DP_mult_204_n531), .B2(DP_mult_204_n535), 
        .A(DP_mult_204_n532), .ZN(DP_mult_204_n526) );
  NOR2_X1 DP_mult_204_U2390 ( .A1(DP_mult_204_n2321), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1217) );
  OAI21_X1 DP_mult_204_U2389 ( .B1(DP_mult_204_n2220), .B2(DP_mult_204_n535), 
        .A(DP_mult_204_n532), .ZN(DP_mult_204_n2277) );
  NAND3_X1 DP_mult_204_U2388 ( .A1(DP_mult_204_n2274), .A2(DP_mult_204_n2275), 
        .A3(DP_mult_204_n2276), .ZN(DP_mult_204_n972) );
  NAND2_X1 DP_mult_204_U2387 ( .A1(DP_mult_204_n996), .A2(DP_mult_204_n1217), 
        .ZN(DP_mult_204_n2276) );
  NAND2_X1 DP_mult_204_U2386 ( .A1(DP_mult_204_n994), .A2(DP_mult_204_n1217), 
        .ZN(DP_mult_204_n2275) );
  NAND2_X1 DP_mult_204_U2385 ( .A1(DP_mult_204_n994), .A2(DP_mult_204_n996), 
        .ZN(DP_mult_204_n2274) );
  XNOR2_X1 DP_mult_204_U2384 ( .A(DP_mult_204_n830), .B(DP_mult_204_n1386), 
        .ZN(DP_mult_204_n2273) );
  XNOR2_X1 DP_mult_204_U2383 ( .A(DP_mult_204_n2205), .B(DP_mult_204_n2273), 
        .ZN(DP_mult_204_n813) );
  NAND2_X1 DP_mult_204_U2382 ( .A1(DP_mult_204_n507), .A2(DP_mult_204_n668), 
        .ZN(DP_mult_204_n498) );
  NAND2_X1 DP_mult_204_U2381 ( .A1(DP_mult_204_n465), .A2(DP_mult_204_n507), 
        .ZN(DP_mult_204_n463) );
  NAND2_X1 DP_mult_204_U2380 ( .A1(DP_mult_204_n478), .A2(DP_mult_204_n507), 
        .ZN(DP_mult_204_n476) );
  XNOR2_X1 DP_mult_204_U2379 ( .A(DP_mult_204_n497), .B(DP_mult_204_n316), 
        .ZN(DP_sw0_coeff_ret0[8]) );
  NOR2_X1 DP_mult_204_U2378 ( .A1(DP_mult_204_n940), .A2(DP_mult_204_n919), 
        .ZN(DP_mult_204_n542) );
  NOR2_X1 DP_mult_204_U2377 ( .A1(DP_mult_204_n919), .A2(DP_mult_204_n940), 
        .ZN(DP_mult_204_n2272) );
  INV_X1 DP_mult_204_U2376 ( .A(DP_mult_204_n1957), .ZN(DP_mult_204_n555) );
  OAI22_X1 DP_mult_204_U2375 ( .A1(DP_mult_204_n2141), .A2(DP_mult_204_n1654), 
        .B1(DP_mult_204_n2042), .B2(DP_mult_204_n1653), .ZN(DP_mult_204_n1359)
         );
  INV_X1 DP_mult_204_U2374 ( .A(DP_mult_204_n2243), .ZN(DP_mult_204_n2337) );
  OR2_X1 DP_mult_204_U2373 ( .A1(DP_mult_204_n2220), .A2(DP_mult_204_n534), 
        .ZN(DP_mult_204_n2271) );
  NAND3_X1 DP_mult_204_U2372 ( .A1(DP_mult_204_n2268), .A2(DP_mult_204_n2269), 
        .A3(DP_mult_204_n2270), .ZN(DP_mult_204_n842) );
  NAND2_X1 DP_mult_204_U2371 ( .A1(DP_mult_204_n849), .A2(DP_mult_204_n864), 
        .ZN(DP_mult_204_n2270) );
  NAND2_X1 DP_mult_204_U2370 ( .A1(DP_mult_204_n862), .A2(DP_mult_204_n864), 
        .ZN(DP_mult_204_n2269) );
  NAND2_X1 DP_mult_204_U2369 ( .A1(DP_mult_204_n862), .A2(DP_mult_204_n849), 
        .ZN(DP_mult_204_n2268) );
  XOR2_X1 DP_mult_204_U2368 ( .A(DP_mult_204_n862), .B(DP_mult_204_n2267), .Z(
        DP_mult_204_n843) );
  XOR2_X1 DP_mult_204_U2367 ( .A(DP_mult_204_n849), .B(DP_mult_204_n864), .Z(
        DP_mult_204_n2267) );
  INV_X1 DP_mult_204_U2366 ( .A(DP_mult_204_n521), .ZN(DP_mult_204_n519) );
  NAND2_X1 DP_mult_204_U2365 ( .A1(DP_mult_204_n670), .A2(DP_mult_204_n2201), 
        .ZN(DP_mult_204_n319) );
  NOR2_X1 DP_mult_204_U2364 ( .A1(DP_mult_204_n1171), .A2(DP_mult_204_n1174), 
        .ZN(DP_mult_204_n633) );
  NAND2_X1 DP_mult_204_U2363 ( .A1(DP_mult_204_n1171), .A2(DP_mult_204_n1174), 
        .ZN(DP_mult_204_n634) );
  NOR2_X1 DP_mult_204_U2362 ( .A1(DP_mult_204_n597), .A2(DP_mult_204_n599), 
        .ZN(DP_mult_204_n595) );
  INV_X1 DP_mult_204_U2361 ( .A(DP_mult_204_n802), .ZN(DP_mult_204_n803) );
  AOI21_X1 DP_mult_204_U2360 ( .B1(DP_mult_204_n2226), .B2(DP_mult_204_n472), 
        .A(DP_mult_204_n459), .ZN(DP_mult_204_n457) );
  NAND2_X1 DP_mult_204_U2359 ( .A1(DP_mult_204_n2226), .A2(DP_mult_204_n461), 
        .ZN(DP_mult_204_n313) );
  OAI22_X1 DP_mult_204_U2358 ( .A1(DP_mult_204_n2140), .A2(DP_mult_204_n1650), 
        .B1(DP_mult_204_n2042), .B2(DP_mult_204_n1649), .ZN(DP_mult_204_n1355)
         );
  NAND2_X1 DP_mult_204_U2357 ( .A1(DP_mult_204_n2266), .A2(DP_mult_204_n2012), 
        .ZN(DP_mult_204_n322) );
  OR2_X1 DP_mult_204_U2356 ( .A1(DP_mult_204_n940), .A2(DP_mult_204_n2086), 
        .ZN(DP_mult_204_n2266) );
  OAI21_X1 DP_mult_204_U2355 ( .B1(DP_mult_204_n2082), .B2(DP_mult_204_n2008), 
        .A(DP_mult_204_n2391), .ZN(DP_mult_204_n1290) );
  INV_X1 DP_mult_204_U2354 ( .A(DP_mult_204_n1937), .ZN(DP_mult_204_n2340) );
  OAI21_X1 DP_mult_204_U2353 ( .B1(DP_mult_204_n2018), .B2(DP_mult_204_n2080), 
        .A(DP_mult_204_n1976), .ZN(DP_mult_204_n1410) );
  NOR2_X1 DP_mult_204_U2352 ( .A1(DP_mult_204_n420), .A2(DP_mult_204_n402), 
        .ZN(DP_mult_204_n400) );
  INV_X1 DP_mult_204_U2351 ( .A(DP_mult_204_n383), .ZN(DP_mult_204_n381) );
  NAND2_X1 DP_mult_204_U2350 ( .A1(DP_mult_204_n963), .A2(DP_mult_204_n982), 
        .ZN(DP_mult_204_n559) );
  OR2_X1 DP_mult_204_U2349 ( .A1(DP_mult_204_n941), .A2(DP_mult_204_n962), 
        .ZN(DP_mult_204_n2265) );
  NAND3_X1 DP_mult_204_U2348 ( .A1(DP_mult_204_n2262), .A2(DP_mult_204_n2263), 
        .A3(DP_mult_204_n2264), .ZN(DP_mult_204_n988) );
  NAND2_X1 DP_mult_204_U2347 ( .A1(DP_mult_204_n997), .A2(DP_mult_204_n1012), 
        .ZN(DP_mult_204_n2264) );
  NAND2_X1 DP_mult_204_U2346 ( .A1(DP_mult_204_n999), .A2(DP_mult_204_n2162), 
        .ZN(DP_mult_204_n2263) );
  NAND2_X1 DP_mult_204_U2345 ( .A1(DP_mult_204_n999), .A2(DP_mult_204_n997), 
        .ZN(DP_mult_204_n2262) );
  XOR2_X1 DP_mult_204_U2344 ( .A(DP_mult_204_n2261), .B(DP_mult_204_n1012), 
        .Z(DP_mult_204_n989) );
  XOR2_X1 DP_mult_204_U2343 ( .A(DP_mult_204_n999), .B(DP_mult_204_n997), .Z(
        DP_mult_204_n2261) );
  NAND3_X1 DP_mult_204_U2342 ( .A1(DP_mult_204_n2258), .A2(DP_mult_204_n2259), 
        .A3(DP_mult_204_n2260), .ZN(DP_mult_204_n1012) );
  NAND2_X1 DP_mult_204_U2341 ( .A1(DP_mult_204_n1439), .A2(DP_mult_204_n1032), 
        .ZN(DP_mult_204_n2260) );
  NAND2_X1 DP_mult_204_U2340 ( .A1(DP_mult_204_n1036), .A2(DP_mult_204_n1032), 
        .ZN(DP_mult_204_n2259) );
  NAND2_X1 DP_mult_204_U2339 ( .A1(DP_mult_204_n1036), .A2(DP_mult_204_n1439), 
        .ZN(DP_mult_204_n2258) );
  NAND2_X1 DP_mult_204_U2338 ( .A1(DP_mult_204_n821), .A2(DP_mult_204_n838), 
        .ZN(DP_mult_204_n503) );
  NOR2_X1 DP_mult_204_U2337 ( .A1(DP_mult_204_n821), .A2(DP_mult_204_n838), 
        .ZN(DP_mult_204_n502) );
  NAND2_X1 DP_mult_204_U2336 ( .A1(DP_mult_204_n668), .A2(DP_mult_204_n503), 
        .ZN(DP_mult_204_n317) );
  OR2_X1 DP_mult_204_U2335 ( .A1(DP_mult_204_n877), .A2(DP_mult_204_n896), 
        .ZN(DP_mult_204_n2256) );
  INV_X1 DP_mult_204_U2334 ( .A(DP_mult_204_n2299), .ZN(DP_mult_204_n2254) );
  INV_X1 DP_mult_204_U2333 ( .A(DP_mult_204_n2299), .ZN(DP_mult_204_n2255) );
  OAI22_X1 DP_mult_204_U2332 ( .A1(DP_mult_204_n2298), .A2(DP_mult_204_n1504), 
        .B1(DP_mult_204_n2322), .B2(DP_mult_204_n1503), .ZN(DP_mult_204_n2253)
         );
  OAI21_X1 DP_mult_204_U2331 ( .B1(DP_mult_204_n2014), .B2(DP_mult_204_n2244), 
        .A(DP_mult_204_n2392), .ZN(DP_mult_204_n1266) );
  OAI22_X1 DP_mult_204_U2330 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1540), 
        .B1(DP_mult_204_n2326), .B2(DP_mult_204_n1539), .ZN(DP_mult_204_n1249)
         );
  OAI22_X1 DP_mult_204_U2329 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1538), 
        .B1(DP_mult_204_n2327), .B2(DP_mult_204_n1537), .ZN(DP_mult_204_n1247)
         );
  OAI22_X1 DP_mult_204_U2328 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1542), 
        .B1(DP_mult_204_n2326), .B2(DP_mult_204_n1541), .ZN(DP_mult_204_n1251)
         );
  OAI22_X1 DP_mult_204_U2327 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1534), 
        .B1(DP_mult_204_n2326), .B2(DP_mult_204_n1533), .ZN(DP_mult_204_n1243)
         );
  OAI22_X1 DP_mult_204_U2326 ( .A1(DP_mult_204_n2302), .A2(DP_mult_204_n1536), 
        .B1(DP_mult_204_n2327), .B2(DP_mult_204_n1535), .ZN(DP_mult_204_n1245)
         );
  NOR2_X1 DP_mult_204_U2325 ( .A1(DP_mult_204_n389), .A2(DP_mult_204_n384), 
        .ZN(DP_mult_204_n382) );
  INV_X1 DP_mult_204_U2324 ( .A(DP_mult_204_n507), .ZN(DP_mult_204_n2251) );
  OAI21_X1 DP_mult_204_U2323 ( .B1(DP_mult_204_n2129), .B2(DP_mult_204_n2060), 
        .A(DP_mult_204_n2386), .ZN(DP_mult_204_n1434) );
  NOR2_X1 DP_mult_204_U2322 ( .A1(DP_mult_204_n983), .A2(DP_mult_204_n1002), 
        .ZN(DP_mult_204_n563) );
  INV_X1 DP_mult_204_U2321 ( .A(DP_mult_204_n2170), .ZN(DP_mult_204_n2313) );
  NAND2_X1 DP_mult_204_U2320 ( .A1(DP_mult_204_n694), .A2(DP_mult_204_n689), 
        .ZN(DP_mult_204_n378) );
  NAND2_X1 DP_mult_204_U2319 ( .A1(DP_mult_204_n422), .A2(DP_mult_204_n356), 
        .ZN(DP_mult_204_n354) );
  NAND2_X1 DP_mult_204_U2318 ( .A1(DP_mult_204_n332), .A2(DP_mult_204_n1996), 
        .ZN(DP_mult_204_n326) );
  INV_X1 DP_mult_204_U2317 ( .A(DP_mult_204_n2365), .ZN(DP_mult_204_n2362) );
  NAND2_X1 DP_mult_204_U2316 ( .A1(DP_mult_204_n857), .A2(DP_mult_204_n876), 
        .ZN(DP_mult_204_n521) );
  INV_X1 DP_mult_204_U2315 ( .A(DP_mult_204_n555), .ZN(DP_mult_204_n2249) );
  OAI21_X1 DP_mult_204_U2314 ( .B1(DP_mult_204_n566), .B2(DP_mult_204_n538), 
        .A(DP_mult_204_n539), .ZN(DP_mult_204_n2247) );
  AOI21_X1 DP_mult_204_U2313 ( .B1(DP_mult_204_n2247), .B2(DP_mult_204_n450), 
        .A(DP_mult_204_n451), .ZN(DP_mult_204_n301) );
  INV_X1 DP_mult_204_U2312 ( .A(DP_coeffs_fb_int[18]), .ZN(DP_mult_204_n2352)
         );
  INV_X1 DP_mult_204_U2311 ( .A(DP_mult_204_n293), .ZN(DP_mult_204_n2303) );
  OAI21_X1 DP_mult_204_U2310 ( .B1(DP_mult_204_n2303), .B2(DP_mult_204_n2071), 
        .A(DP_mult_204_n2393), .ZN(DP_mult_204_n1242) );
  XNOR2_X1 DP_mult_204_U2309 ( .A(DP_mult_204_n1935), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1733) );
  XNOR2_X1 DP_mult_204_U2308 ( .A(DP_mult_204_n2354), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1683) );
  XNOR2_X1 DP_mult_204_U2307 ( .A(DP_mult_204_n2357), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1658) );
  XNOR2_X1 DP_mult_204_U2306 ( .A(DP_mult_204_n2351), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1708) );
  XNOR2_X1 DP_mult_204_U2305 ( .A(DP_mult_204_n2346), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1758) );
  XNOR2_X1 DP_mult_204_U2304 ( .A(DP_mult_204_n2360), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1633) );
  XNOR2_X1 DP_mult_204_U2303 ( .A(DP_mult_204_n2364), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1608) );
  XNOR2_X1 DP_mult_204_U2302 ( .A(DP_mult_204_n2370), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1558) );
  XNOR2_X1 DP_mult_204_U2301 ( .A(DP_mult_204_n2366), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1583) );
  XNOR2_X1 DP_mult_204_U2300 ( .A(DP_mult_204_n2374), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1533) );
  XNOR2_X1 DP_mult_204_U2299 ( .A(DP_mult_204_n2378), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1508) );
  XNOR2_X1 DP_mult_204_U2298 ( .A(DP_mult_204_n2382), .B(DP_sw0_22_), .ZN(
        DP_mult_204_n1483) );
  XNOR2_X1 DP_mult_204_U2297 ( .A(DP_sw0_23_), .B(DP_mult_204_n2381), .ZN(
        DP_mult_204_n1482) );
  NAND2_X1 DP_mult_204_U2296 ( .A1(DP_mult_204_n2217), .A2(DP_mult_204_n496), 
        .ZN(DP_mult_204_n316) );
  NAND2_X1 DP_mult_204_U2295 ( .A1(DP_mult_204_n2204), .A2(DP_mult_204_n514), 
        .ZN(DP_mult_204_n318) );
  XNOR2_X1 DP_mult_204_U2294 ( .A(DP_mult_204_n515), .B(DP_mult_204_n318), 
        .ZN(DP_sw0_coeff_ret0[6]) );
  XNOR2_X1 DP_mult_204_U2293 ( .A(DP_mult_204_n522), .B(DP_mult_204_n319), 
        .ZN(DP_sw0_coeff_ret0[5]) );
  XNOR2_X1 DP_mult_204_U2292 ( .A(DP_mult_204_n504), .B(DP_mult_204_n317), 
        .ZN(DP_sw0_coeff_ret0[7]) );
  NAND2_X1 DP_mult_204_U2291 ( .A1(DP_mult_204_n2007), .A2(DP_mult_204_n481), 
        .ZN(DP_mult_204_n315) );
  XNOR2_X1 DP_mult_204_U2290 ( .A(DP_mult_204_n486), .B(DP_mult_204_n315), 
        .ZN(DP_sw0_coeff_ret0[9]) );
  XNOR2_X1 DP_mult_204_U2289 ( .A(DP_mult_204_n2356), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1680) );
  INV_X1 DP_mult_204_U2288 ( .A(DP_mult_204_n285), .ZN(DP_mult_204_n2310) );
  NAND2_X1 DP_mult_204_U2287 ( .A1(DP_mult_204_n2256), .A2(DP_mult_204_n532), 
        .ZN(DP_mult_204_n320) );
  XNOR2_X1 DP_mult_204_U2286 ( .A(DP_mult_204_n533), .B(DP_mult_204_n320), 
        .ZN(DP_sw0_coeff_ret0[4]) );
  INV_X1 DP_mult_204_U2285 ( .A(DP_mult_204_n1757), .ZN(DP_mult_204_n2385) );
  OAI21_X1 DP_mult_204_U2284 ( .B1(DP_coeffs_fb_int[23]), .B2(
        DP_mult_204_n2242), .A(DP_mult_204_n2385), .ZN(DP_mult_204_n1458) );
  AOI21_X1 DP_mult_204_U2283 ( .B1(DP_mult_204_n565), .B2(DP_mult_204_n545), 
        .A(DP_mult_204_n546), .ZN(DP_mult_204_n544) );
  XOR2_X1 DP_mult_204_U2282 ( .A(DP_mult_204_n544), .B(DP_mult_204_n322), .Z(
        DP_sw0_coeff_ret0[2]) );
  INV_X1 DP_mult_204_U2281 ( .A(DP_coeffs_fb_int[8]), .ZN(DP_mult_204_n2368)
         );
  INV_X1 DP_mult_204_U2280 ( .A(DP_coeffs_fb_int[6]), .ZN(DP_mult_204_n2372)
         );
  INV_X1 DP_mult_204_U2279 ( .A(DP_coeffs_fb_int[14]), .ZN(DP_mult_204_n2358)
         );
  INV_X1 DP_mult_204_U2278 ( .A(DP_coeffs_fb_int[0]), .ZN(DP_mult_204_n2383)
         );
  INV_X1 DP_mult_204_U2277 ( .A(DP_coeffs_fb_int[10]), .ZN(DP_mult_204_n2365)
         );
  INV_X1 DP_mult_204_U2276 ( .A(DP_coeffs_fb_int[12]), .ZN(DP_mult_204_n2361)
         );
  XNOR2_X1 DP_mult_204_U2275 ( .A(DP_sw0_11_), .B(DP_mult_204_n2382), .ZN(
        DP_mult_204_n1494) );
  XNOR2_X1 DP_mult_204_U2274 ( .A(DP_sw0_21_), .B(DP_mult_204_n2381), .ZN(
        DP_mult_204_n1484) );
  XNOR2_X1 DP_mult_204_U2273 ( .A(DP_sw0_19_), .B(DP_mult_204_n2382), .ZN(
        DP_mult_204_n1486) );
  XNOR2_X1 DP_mult_204_U2272 ( .A(DP_sw0_15_), .B(DP_mult_204_n2381), .ZN(
        DP_mult_204_n1490) );
  XNOR2_X1 DP_mult_204_U2271 ( .A(DP_sw0_17_), .B(DP_mult_204_n2381), .ZN(
        DP_mult_204_n1488) );
  XNOR2_X1 DP_mult_204_U2270 ( .A(DP_sw0_13_), .B(DP_mult_204_n2381), .ZN(
        DP_mult_204_n1492) );
  XNOR2_X1 DP_mult_204_U2269 ( .A(DP_mult_204_n2370), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1580) );
  XNOR2_X1 DP_mult_204_U2268 ( .A(DP_sw0_9_), .B(DP_mult_204_n2382), .ZN(
        DP_mult_204_n1496) );
  XNOR2_X1 DP_mult_204_U2267 ( .A(DP_sw0_5_), .B(DP_mult_204_n2356), .ZN(
        DP_mult_204_n1675) );
  XNOR2_X1 DP_mult_204_U2266 ( .A(DP_sw0_9_), .B(DP_mult_204_n2355), .ZN(
        DP_mult_204_n1671) );
  XNOR2_X1 DP_mult_204_U2265 ( .A(DP_sw0_5_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1700) );
  XNOR2_X1 DP_mult_204_U2264 ( .A(DP_sw0_9_), .B(DP_mult_204_n2348), .ZN(
        DP_mult_204_n1746) );
  XNOR2_X1 DP_mult_204_U2263 ( .A(DP_sw0_9_), .B(DP_mult_204_n2350), .ZN(
        DP_mult_204_n1721) );
  XNOR2_X1 DP_mult_204_U2262 ( .A(DP_sw0_9_), .B(DP_mult_204_n2378), .ZN(
        DP_mult_204_n1521) );
  XNOR2_X1 DP_mult_204_U2261 ( .A(DP_sw0_5_), .B(DP_mult_204_n2351), .ZN(
        DP_mult_204_n1725) );
  XNOR2_X1 DP_mult_204_U2260 ( .A(DP_sw0_7_), .B(DP_mult_204_n2348), .ZN(
        DP_mult_204_n1748) );
  XNOR2_X1 DP_mult_204_U2259 ( .A(DP_sw0_7_), .B(DP_mult_204_n2355), .ZN(
        DP_mult_204_n1673) );
  XNOR2_X1 DP_mult_204_U2258 ( .A(DP_sw0_7_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1698) );
  XNOR2_X1 DP_mult_204_U2257 ( .A(DP_sw0_5_), .B(DP_mult_204_n2362), .ZN(
        DP_mult_204_n1625) );
  XNOR2_X1 DP_mult_204_U2256 ( .A(DP_sw0_5_), .B(DP_mult_204_n2348), .ZN(
        DP_mult_204_n1750) );
  XNOR2_X1 DP_mult_204_U2255 ( .A(DP_sw0_5_), .B(DP_mult_204_n2381), .ZN(
        DP_mult_204_n1500) );
  XNOR2_X1 DP_mult_204_U2254 ( .A(DP_sw0_5_), .B(DP_mult_204_n2366), .ZN(
        DP_mult_204_n1600) );
  XNOR2_X1 DP_mult_204_U2253 ( .A(DP_sw0_7_), .B(DP_mult_204_n2381), .ZN(
        DP_mult_204_n1498) );
  XNOR2_X1 DP_mult_204_U2252 ( .A(DP_sw0_7_), .B(DP_mult_204_n2373), .ZN(
        DP_mult_204_n1548) );
  XNOR2_X1 DP_mult_204_U2251 ( .A(DP_sw0_7_), .B(DP_mult_204_n2350), .ZN(
        DP_mult_204_n1723) );
  XNOR2_X1 DP_mult_204_U2250 ( .A(DP_sw0_9_), .B(DP_mult_204_n2373), .ZN(
        DP_mult_204_n1546) );
  XNOR2_X1 DP_mult_204_U2249 ( .A(DP_sw0_5_), .B(DP_mult_204_n2377), .ZN(
        DP_mult_204_n1525) );
  XNOR2_X1 DP_mult_204_U2248 ( .A(DP_sw0_9_), .B(DP_mult_204_n2364), .ZN(
        DP_mult_204_n1621) );
  XNOR2_X1 DP_mult_204_U2247 ( .A(DP_sw0_7_), .B(DP_mult_204_n2376), .ZN(
        DP_mult_204_n1523) );
  XNOR2_X1 DP_mult_204_U2246 ( .A(DP_sw0_7_), .B(DP_mult_204_n2363), .ZN(
        DP_mult_204_n1623) );
  XNOR2_X1 DP_mult_204_U2245 ( .A(DP_sw0_7_), .B(DP_mult_204_n2370), .ZN(
        DP_mult_204_n1573) );
  XNOR2_X1 DP_mult_204_U2244 ( .A(DP_sw0_9_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1696) );
  XNOR2_X1 DP_mult_204_U2243 ( .A(DP_sw0_5_), .B(DP_mult_204_n2134), .ZN(
        DP_mult_204_n1650) );
  XNOR2_X1 DP_mult_204_U2242 ( .A(DP_sw0_9_), .B(DP_mult_204_n2371), .ZN(
        DP_mult_204_n1571) );
  XNOR2_X1 DP_mult_204_U2241 ( .A(DP_sw0_9_), .B(DP_mult_204_n2367), .ZN(
        DP_mult_204_n1596) );
  XNOR2_X1 DP_mult_204_U2240 ( .A(DP_sw0_5_), .B(DP_mult_204_n2370), .ZN(
        DP_mult_204_n1575) );
  XNOR2_X1 DP_mult_204_U2239 ( .A(DP_sw0_5_), .B(DP_mult_204_n2373), .ZN(
        DP_mult_204_n1550) );
  XNOR2_X1 DP_mult_204_U2238 ( .A(DP_sw0_7_), .B(DP_mult_204_n2366), .ZN(
        DP_mult_204_n1598) );
  XNOR2_X1 DP_mult_204_U2237 ( .A(DP_sw0_1_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1704) );
  XNOR2_X1 DP_mult_204_U2236 ( .A(DP_sw0_1_), .B(DP_mult_204_n2356), .ZN(
        DP_mult_204_n1679) );
  XNOR2_X1 DP_mult_204_U2235 ( .A(DP_sw0_1_), .B(DP_mult_204_n2350), .ZN(
        DP_mult_204_n1729) );
  XNOR2_X1 DP_mult_204_U2234 ( .A(DP_sw0_1_), .B(DP_mult_204_n2135), .ZN(
        DP_mult_204_n1654) );
  XNOR2_X1 DP_mult_204_U2233 ( .A(DP_sw0_1_), .B(DP_mult_204_n2363), .ZN(
        DP_mult_204_n1629) );
  XNOR2_X1 DP_mult_204_U2232 ( .A(DP_sw0_1_), .B(DP_mult_204_n2348), .ZN(
        DP_mult_204_n1754) );
  XNOR2_X1 DP_mult_204_U2231 ( .A(DP_sw0_1_), .B(DP_mult_204_n2370), .ZN(
        DP_mult_204_n1579) );
  XNOR2_X1 DP_mult_204_U2230 ( .A(DP_sw0_1_), .B(DP_mult_204_n2379), .ZN(
        DP_mult_204_n1529) );
  XNOR2_X1 DP_mult_204_U2229 ( .A(DP_sw0_1_), .B(DP_mult_204_n2373), .ZN(
        DP_mult_204_n1554) );
  XNOR2_X1 DP_mult_204_U2228 ( .A(DP_sw0_1_), .B(DP_mult_204_n2367), .ZN(
        DP_mult_204_n1604) );
  XNOR2_X1 DP_mult_204_U2227 ( .A(DP_sw0_3_), .B(DP_mult_204_n2355), .ZN(
        DP_mult_204_n1677) );
  XNOR2_X1 DP_mult_204_U2226 ( .A(DP_sw0_3_), .B(DP_mult_204_n2351), .ZN(
        DP_mult_204_n1727) );
  XNOR2_X1 DP_mult_204_U2225 ( .A(DP_sw0_3_), .B(DP_mult_204_n2348), .ZN(
        DP_mult_204_n1752) );
  XNOR2_X1 DP_mult_204_U2224 ( .A(DP_sw0_3_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1702) );
  XNOR2_X1 DP_mult_204_U2223 ( .A(DP_sw0_3_), .B(DP_mult_204_n2381), .ZN(
        DP_mult_204_n1502) );
  XNOR2_X1 DP_mult_204_U2222 ( .A(DP_sw0_3_), .B(DP_mult_204_n2367), .ZN(
        DP_mult_204_n1602) );
  XNOR2_X1 DP_mult_204_U2221 ( .A(DP_sw0_3_), .B(DP_mult_204_n2373), .ZN(
        DP_mult_204_n1552) );
  XNOR2_X1 DP_mult_204_U2220 ( .A(DP_sw0_3_), .B(DP_mult_204_n2376), .ZN(
        DP_mult_204_n1527) );
  XNOR2_X1 DP_mult_204_U2219 ( .A(DP_sw0_3_), .B(DP_mult_204_n2371), .ZN(
        DP_mult_204_n1577) );
  XNOR2_X1 DP_mult_204_U2218 ( .A(DP_sw0_3_), .B(DP_mult_204_n2364), .ZN(
        DP_mult_204_n1627) );
  XNOR2_X1 DP_mult_204_U2217 ( .A(DP_mult_204_n2354), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1705) );
  XNOR2_X1 DP_mult_204_U2216 ( .A(DP_mult_204_n2362), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1630) );
  XNOR2_X1 DP_mult_204_U2215 ( .A(DP_sw0_9_), .B(DP_mult_204_n2135), .ZN(
        DP_mult_204_n1646) );
  XNOR2_X1 DP_mult_204_U2214 ( .A(DP_mult_204_n2350), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1730) );
  OAI22_X1 DP_mult_204_U2213 ( .A1(DP_mult_204_n2120), .A2(DP_mult_204_n1776), 
        .B1(DP_mult_204_n1775), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1477)
         );
  XNOR2_X1 DP_mult_204_U2212 ( .A(DP_mult_204_n2348), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1755) );
  OAI22_X1 DP_mult_204_U2211 ( .A1(DP_mult_204_n2121), .A2(DP_mult_204_n1778), 
        .B1(DP_mult_204_n1777), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1479)
         );
  XNOR2_X1 DP_mult_204_U2210 ( .A(DP_sw0_23_), .B(DP_mult_204_n2377), .ZN(
        DP_mult_204_n1507) );
  XNOR2_X1 DP_mult_204_U2209 ( .A(DP_sw0_23_), .B(DP_mult_204_n2374), .ZN(
        DP_mult_204_n1532) );
  XNOR2_X1 DP_mult_204_U2208 ( .A(DP_sw0_23_), .B(DP_mult_204_n2366), .ZN(
        DP_mult_204_n1582) );
  XNOR2_X1 DP_mult_204_U2207 ( .A(DP_sw0_23_), .B(DP_mult_204_n2370), .ZN(
        DP_mult_204_n1557) );
  XNOR2_X1 DP_mult_204_U2206 ( .A(DP_sw0_23_), .B(DP_mult_204_n2356), .ZN(
        DP_mult_204_n1657) );
  XNOR2_X1 DP_mult_204_U2205 ( .A(DP_sw0_23_), .B(DP_mult_204_n2364), .ZN(
        DP_mult_204_n1607) );
  XNOR2_X1 DP_mult_204_U2204 ( .A(DP_sw0_23_), .B(DP_mult_204_n2135), .ZN(
        DP_mult_204_n1632) );
  XNOR2_X1 DP_mult_204_U2203 ( .A(DP_sw0_23_), .B(DP_mult_204_n2350), .ZN(
        DP_mult_204_n1707) );
  XNOR2_X1 DP_mult_204_U2202 ( .A(DP_sw0_23_), .B(DP_mult_204_n2109), .ZN(
        DP_mult_204_n1682) );
  XNOR2_X1 DP_mult_204_U2201 ( .A(DP_sw0_23_), .B(DP_mult_204_n1935), .ZN(
        DP_mult_204_n1732) );
  XNOR2_X1 DP_mult_204_U2200 ( .A(DP_sw0_3_), .B(DP_mult_204_n2134), .ZN(
        DP_mult_204_n1652) );
  XNOR2_X1 DP_mult_204_U2199 ( .A(DP_sw0_7_), .B(DP_mult_204_n2134), .ZN(
        DP_mult_204_n1648) );
  XNOR2_X1 DP_mult_204_U2198 ( .A(DP_mult_204_n2378), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1518) );
  XNOR2_X1 DP_mult_204_U2197 ( .A(DP_mult_204_n2348), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1753) );
  XNOR2_X1 DP_mult_204_U2196 ( .A(DP_mult_204_n2351), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1726) );
  XNOR2_X1 DP_mult_204_U2195 ( .A(DP_mult_204_n2359), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1653) );
  XNOR2_X1 DP_mult_204_U2194 ( .A(DP_mult_204_n2350), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1728) );
  XNOR2_X1 DP_mult_204_U2193 ( .A(DP_mult_204_n2355), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1676) );
  XNOR2_X1 DP_mult_204_U2192 ( .A(DP_mult_204_n2353), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1701) );
  XNOR2_X1 DP_mult_204_U2191 ( .A(DP_mult_204_n2374), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1543) );
  XNOR2_X1 DP_mult_204_U2190 ( .A(DP_mult_204_n2348), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1751) );
  XNOR2_X1 DP_mult_204_U2189 ( .A(DP_mult_204_n2367), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1601) );
  XNOR2_X1 DP_mult_204_U2188 ( .A(DP_mult_204_n2355), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1678) );
  XNOR2_X1 DP_mult_204_U2187 ( .A(DP_mult_204_n2353), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1703) );
  XNOR2_X1 DP_mult_204_U2186 ( .A(DP_mult_204_n2381), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1493) );
  XNOR2_X1 DP_mult_204_U2185 ( .A(DP_mult_204_n2370), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1578) );
  XNOR2_X1 DP_mult_204_U2184 ( .A(DP_mult_204_n2367), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1593) );
  XNOR2_X1 DP_mult_204_U2183 ( .A(DP_mult_204_n2351), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1718) );
  XNOR2_X1 DP_mult_204_U2182 ( .A(DP_mult_204_n2363), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1626) );
  XNOR2_X1 DP_mult_204_U2181 ( .A(DP_mult_204_n2364), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1618) );
  XNOR2_X1 DP_mult_204_U2180 ( .A(DP_mult_204_n2381), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1501) );
  XNOR2_X1 DP_mult_204_U2179 ( .A(DP_mult_204_n1935), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1743) );
  XNOR2_X1 DP_mult_204_U2178 ( .A(DP_mult_204_n2371), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1568) );
  XNOR2_X1 DP_mult_204_U2177 ( .A(DP_mult_204_n2366), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1603) );
  XNOR2_X1 DP_mult_204_U2176 ( .A(DP_mult_204_n2379), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1528) );
  XNOR2_X1 DP_mult_204_U2175 ( .A(DP_mult_204_n2353), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1693) );
  XNOR2_X1 DP_mult_204_U2174 ( .A(DP_mult_204_n2376), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1526) );
  XNOR2_X1 DP_mult_204_U2173 ( .A(DP_mult_204_n2356), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1668) );
  XNOR2_X1 DP_mult_204_U2172 ( .A(DP_mult_204_n2373), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1553) );
  XNOR2_X1 DP_mult_204_U2171 ( .A(DP_mult_204_n2371), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1576) );
  XNOR2_X1 DP_mult_204_U2170 ( .A(DP_mult_204_n2373), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1551) );
  XNOR2_X1 DP_mult_204_U2169 ( .A(DP_mult_204_n2363), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1628) );
  XNOR2_X1 DP_mult_204_U2168 ( .A(DP_mult_204_n2374), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1535) );
  XNOR2_X1 DP_mult_204_U2167 ( .A(DP_mult_204_n2378), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1510) );
  XNOR2_X1 DP_mult_204_U2166 ( .A(DP_mult_204_n2381), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1487) );
  XNOR2_X1 DP_mult_204_U2165 ( .A(DP_mult_204_n2382), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1485) );
  XNOR2_X1 DP_mult_204_U2164 ( .A(DP_mult_204_n2350), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1720) );
  XNOR2_X1 DP_mult_204_U2163 ( .A(DP_mult_204_n2369), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1560) );
  XNOR2_X1 DP_mult_204_U2162 ( .A(DP_mult_204_n2379), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1514) );
  XNOR2_X1 DP_mult_204_U2161 ( .A(DP_mult_204_n2382), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1489) );
  XNOR2_X1 DP_mult_204_U2160 ( .A(DP_mult_204_n2377), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1512) );
  XNOR2_X1 DP_mult_204_U2159 ( .A(DP_mult_204_n2348), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1747) );
  XNOR2_X1 DP_mult_204_U2158 ( .A(DP_mult_204_n2348), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1745) );
  XNOR2_X1 DP_mult_204_U2157 ( .A(DP_mult_204_n2374), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1537) );
  XNOR2_X1 DP_mult_204_U2156 ( .A(DP_mult_204_n2370), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1566) );
  XNOR2_X1 DP_mult_204_U2155 ( .A(DP_mult_204_n2356), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1660) );
  XNOR2_X1 DP_mult_204_U2154 ( .A(DP_mult_204_n2351), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1722) );
  XNOR2_X1 DP_mult_204_U2153 ( .A(DP_mult_204_n2382), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1495) );
  XNOR2_X1 DP_mult_204_U2152 ( .A(DP_mult_204_n2374), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1541) );
  XNOR2_X1 DP_mult_204_U2151 ( .A(DP_mult_204_n2360), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1635) );
  XNOR2_X1 DP_mult_204_U2150 ( .A(DP_mult_204_n2348), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1749) );
  XNOR2_X1 DP_mult_204_U2149 ( .A(DP_mult_204_n2379), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1520) );
  XNOR2_X1 DP_mult_204_U2148 ( .A(DP_mult_204_n2382), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1491) );
  XNOR2_X1 DP_mult_204_U2147 ( .A(DP_mult_204_n2353), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1699) );
  XNOR2_X1 DP_mult_204_U2146 ( .A(DP_mult_204_n2366), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1587) );
  XNOR2_X1 DP_mult_204_U2145 ( .A(DP_mult_204_n2366), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1589) );
  XNOR2_X1 DP_mult_204_U2144 ( .A(DP_mult_204_n2350), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1716) );
  XNOR2_X1 DP_mult_204_U2143 ( .A(DP_mult_204_n2362), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1612) );
  XNOR2_X1 DP_mult_204_U2142 ( .A(DP_mult_204_n2353), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1687) );
  XNOR2_X1 DP_mult_204_U2141 ( .A(DP_mult_204_n2369), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1562) );
  XNOR2_X1 DP_mult_204_U2140 ( .A(DP_mult_204_n2371), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1564) );
  XNOR2_X1 DP_mult_204_U2139 ( .A(DP_mult_204_n2355), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1670) );
  XNOR2_X1 DP_mult_204_U2138 ( .A(DP_mult_204_n2364), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1620) );
  XNOR2_X1 DP_mult_204_U2137 ( .A(DP_mult_204_n2363), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1610) );
  XNOR2_X1 DP_mult_204_U2136 ( .A(DP_mult_204_n1935), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1739) );
  XNOR2_X1 DP_mult_204_U2135 ( .A(DP_mult_204_n2356), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1664) );
  XNOR2_X1 DP_mult_204_U2134 ( .A(DP_mult_204_n2366), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1585) );
  XNOR2_X1 DP_mult_204_U2133 ( .A(DP_mult_204_n2374), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1539) );
  XNOR2_X1 DP_mult_204_U2132 ( .A(DP_mult_204_n2360), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1639) );
  XNOR2_X1 DP_mult_204_U2131 ( .A(DP_mult_204_n2354), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1685) );
  XNOR2_X1 DP_mult_204_U2130 ( .A(DP_mult_204_n2370), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1570) );
  XNOR2_X1 DP_mult_204_U2129 ( .A(DP_mult_204_n2353), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1691) );
  XNOR2_X1 DP_mult_204_U2128 ( .A(DP_mult_204_n2377), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1516) );
  XNOR2_X1 DP_mult_204_U2127 ( .A(DP_mult_204_n2356), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1674) );
  XNOR2_X1 DP_mult_204_U2126 ( .A(DP_mult_204_n2351), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1724) );
  XNOR2_X1 DP_mult_204_U2125 ( .A(DP_mult_204_n2378), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1522) );
  XNOR2_X1 DP_mult_204_U2124 ( .A(DP_mult_204_n2373), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1547) );
  XNOR2_X1 DP_mult_204_U2123 ( .A(DP_mult_204_n2353), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1695) );
  XNOR2_X1 DP_mult_204_U2122 ( .A(DP_mult_204_n2355), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1672) );
  XNOR2_X1 DP_mult_204_U2121 ( .A(DP_mult_204_n2362), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1622) );
  XNOR2_X1 DP_mult_204_U2120 ( .A(DP_mult_204_n2351), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1712) );
  XNOR2_X1 DP_mult_204_U2119 ( .A(DP_mult_204_n2351), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1710) );
  XNOR2_X1 DP_mult_204_U2118 ( .A(DP_mult_204_n2364), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1624) );
  XNOR2_X1 DP_mult_204_U2117 ( .A(DP_mult_204_n2373), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1549) );
  XNOR2_X1 DP_mult_204_U2116 ( .A(DP_mult_204_n2348), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1737) );
  XNOR2_X1 DP_mult_204_U2115 ( .A(DP_mult_204_n2376), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1524) );
  XNOR2_X1 DP_mult_204_U2114 ( .A(DP_mult_204_n2364), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1616) );
  XNOR2_X1 DP_mult_204_U2113 ( .A(DP_mult_204_n2357), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1662) );
  XNOR2_X1 DP_mult_204_U2112 ( .A(DP_mult_204_n2354), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1689) );
  XNOR2_X1 DP_mult_204_U2111 ( .A(DP_mult_204_n1935), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1735) );
  XNOR2_X1 DP_mult_204_U2110 ( .A(DP_mult_204_n2366), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1597) );
  XNOR2_X1 DP_mult_204_U2109 ( .A(DP_mult_204_n2369), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1574) );
  XNOR2_X1 DP_mult_204_U2108 ( .A(DP_mult_204_n2353), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1697) );
  XNOR2_X1 DP_mult_204_U2107 ( .A(DP_mult_204_n2382), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1499) );
  XNOR2_X1 DP_mult_204_U2106 ( .A(DP_mult_204_n2348), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1741) );
  XNOR2_X1 DP_mult_204_U2105 ( .A(DP_mult_204_n2350), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1714) );
  XNOR2_X1 DP_mult_204_U2104 ( .A(DP_mult_204_n2367), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1599) );
  XNOR2_X1 DP_mult_204_U2103 ( .A(DP_mult_204_n2382), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1497) );
  XNOR2_X1 DP_mult_204_U2102 ( .A(DP_mult_204_n2371), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1572) );
  XNOR2_X1 DP_mult_204_U2101 ( .A(DP_mult_204_n2366), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1595) );
  XNOR2_X1 DP_mult_204_U2100 ( .A(DP_mult_204_n2359), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1641) );
  XNOR2_X1 DP_mult_204_U2099 ( .A(DP_mult_204_n2367), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1591) );
  XNOR2_X1 DP_mult_204_U2098 ( .A(DP_mult_204_n2359), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1637) );
  XNOR2_X1 DP_mult_204_U2097 ( .A(DP_mult_204_n2355), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1666) );
  XNOR2_X1 DP_mult_204_U2096 ( .A(DP_mult_204_n2373), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1545) );
  XNOR2_X1 DP_mult_204_U2095 ( .A(DP_mult_204_n2363), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1614) );
  XNOR2_X1 DP_mult_204_U2094 ( .A(DP_mult_204_n2346), .B(DP_sw0_20_), .ZN(
        DP_mult_204_n1760) );
  XNOR2_X1 DP_mult_204_U2093 ( .A(DP_mult_204_n2345), .B(DP_sw0_14_), .ZN(
        DP_mult_204_n1766) );
  XNOR2_X1 DP_mult_204_U2092 ( .A(DP_mult_204_n2346), .B(DP_sw0_16_), .ZN(
        DP_mult_204_n1764) );
  XNOR2_X1 DP_mult_204_U2091 ( .A(DP_mult_204_n2345), .B(DP_sw0_18_), .ZN(
        DP_mult_204_n1762) );
  XNOR2_X1 DP_mult_204_U2090 ( .A(DP_mult_204_n2346), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1780) );
  XNOR2_X1 DP_mult_204_U2089 ( .A(DP_mult_204_n2345), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1768) );
  XNOR2_X1 DP_mult_204_U2088 ( .A(DP_mult_204_n2359), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1651) );
  XNOR2_X1 DP_mult_204_U2087 ( .A(DP_mult_204_n2359), .B(DP_sw0_12_), .ZN(
        DP_mult_204_n1643) );
  XNOR2_X1 DP_mult_204_U2086 ( .A(DP_mult_204_n2382), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1503) );
  XNOR2_X1 DP_mult_204_U2085 ( .A(DP_mult_204_n2359), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1645) );
  XNOR2_X1 DP_mult_204_U2084 ( .A(DP_mult_204_n2359), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1649) );
  XNOR2_X1 DP_mult_204_U2083 ( .A(DP_mult_204_n2360), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1655) );
  XNOR2_X1 DP_mult_204_U2082 ( .A(DP_mult_204_n2367), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1605) );
  XNOR2_X1 DP_mult_204_U2081 ( .A(DP_mult_204_n2374), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1555) );
  XNOR2_X1 DP_mult_204_U2080 ( .A(DP_mult_204_n2345), .B(DP_sw0_4_), .ZN(
        DP_mult_204_n1776) );
  XNOR2_X1 DP_mult_204_U2079 ( .A(DP_mult_204_n2345), .B(DP_sw0_2_), .ZN(
        DP_mult_204_n1778) );
  XNOR2_X1 DP_mult_204_U2078 ( .A(DP_mult_204_n2345), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1772) );
  XNOR2_X1 DP_mult_204_U2077 ( .A(DP_mult_204_n2345), .B(DP_sw0_6_), .ZN(
        DP_mult_204_n1774) );
  XNOR2_X1 DP_mult_204_U2076 ( .A(DP_mult_204_n2345), .B(DP_sw0_10_), .ZN(
        DP_mult_204_n1770) );
  XNOR2_X1 DP_mult_204_U2075 ( .A(DP_mult_204_n2359), .B(DP_sw0_8_), .ZN(
        DP_mult_204_n1647) );
  XNOR2_X1 DP_mult_204_U2074 ( .A(DP_mult_204_n2376), .B(DP_sw0_0_), .ZN(
        DP_mult_204_n1530) );
  INV_X1 DP_mult_204_U2073 ( .A(DP_mult_204_n1482), .ZN(DP_mult_204_n2395) );
  OAI21_X1 DP_mult_204_U2072 ( .B1(DP_mult_204_n2299), .B2(DP_mult_204_n2063), 
        .A(DP_mult_204_n2395), .ZN(DP_mult_204_n1194) );
  INV_X1 DP_mult_204_U2071 ( .A(DP_mult_204_n1582), .ZN(DP_mult_204_n2391) );
  INV_X1 DP_mult_204_U2070 ( .A(DP_mult_204_n1956), .ZN(DP_mult_204_n2386) );
  INV_X1 DP_mult_204_U2069 ( .A(DP_mult_204_n724), .ZN(DP_mult_204_n725) );
  INV_X1 DP_mult_204_U2068 ( .A(DP_mult_204_n1657), .ZN(DP_mult_204_n2388) );
  NAND2_X1 DP_mult_204_U2067 ( .A1(DP_mult_204_n2345), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1781) );
  OAI22_X1 DP_mult_204_U2066 ( .A1(DP_mult_204_n2121), .A2(DP_mult_204_n1780), 
        .B1(DP_mult_204_n1779), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1481)
         );
  CLKBUF_X1 DP_mult_204_U2065 ( .A(DP_mult_204_n251), .Z(DP_mult_204_n2343) );
  XNOR2_X1 DP_mult_204_U2064 ( .A(DP_mult_204_n1036), .B(DP_mult_204_n1439), 
        .ZN(DP_mult_204_n2241) );
  XNOR2_X1 DP_mult_204_U2063 ( .A(DP_mult_204_n2241), .B(DP_mult_204_n1032), 
        .ZN(DP_mult_204_n1013) );
  INV_X1 DP_mult_204_U2062 ( .A(DP_mult_204_n1607), .ZN(DP_mult_204_n2390) );
  OAI21_X1 DP_mult_204_U2061 ( .B1(DP_mult_204_n2016), .B2(DP_mult_204_n1968), 
        .A(DP_mult_204_n2390), .ZN(DP_mult_204_n1314) );
  INV_X1 DP_mult_204_U2060 ( .A(DP_mult_204_n1557), .ZN(DP_mult_204_n2392) );
  OAI22_X1 DP_mult_204_U2059 ( .A1(DP_mult_204_n2141), .A2(DP_mult_204_n1648), 
        .B1(DP_mult_204_n2118), .B2(DP_mult_204_n1647), .ZN(DP_mult_204_n1353)
         );
  NOR2_X1 DP_mult_204_U2058 ( .A1(DP_mult_204_n2329), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1289) );
  NOR2_X1 DP_mult_204_U2057 ( .A1(DP_mult_204_n1970), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1337) );
  NOR2_X1 DP_mult_204_U2056 ( .A1(DP_mult_204_n2326), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1265) );
  OAI22_X1 DP_mult_204_U2055 ( .A1(DP_mult_204_n2140), .A2(DP_mult_204_n1645), 
        .B1(DP_mult_204_n1644), .B2(DP_mult_204_n2181), .ZN(DP_mult_204_n1350)
         );
  NOR2_X1 DP_mult_204_U2054 ( .A1(DP_mult_204_n2325), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1241) );
  OAI22_X1 DP_mult_204_U2053 ( .A1(DP_mult_204_n2320), .A2(DP_mult_204_n1771), 
        .B1(DP_mult_204_n1770), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1472)
         );
  NOR2_X1 DP_mult_204_U2052 ( .A1(DP_mult_204_n2042), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1361) );
  OAI22_X1 DP_mult_204_U2051 ( .A1(DP_mult_204_n2121), .A2(DP_mult_204_n1774), 
        .B1(DP_mult_204_n1773), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1475)
         );
  OAI21_X1 DP_mult_204_U2050 ( .B1(DP_mult_204_n1987), .B2(DP_mult_204_n2102), 
        .A(DP_mult_204_n2388), .ZN(DP_mult_204_n1362) );
  OAI22_X1 DP_mult_204_U2049 ( .A1(DP_mult_204_n2121), .A2(DP_mult_204_n1772), 
        .B1(DP_mult_204_n1771), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1473)
         );
  OAI22_X1 DP_mult_204_U2048 ( .A1(DP_mult_204_n2120), .A2(DP_mult_204_n1775), 
        .B1(DP_mult_204_n1774), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1476)
         );
  NOR2_X1 DP_mult_204_U2047 ( .A1(DP_mult_204_n2331), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1313) );
  OAI22_X1 DP_mult_204_U2046 ( .A1(DP_mult_204_n2120), .A2(DP_mult_204_n1769), 
        .B1(DP_mult_204_n1768), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1470)
         );
  OAI22_X1 DP_mult_204_U2045 ( .A1(DP_mult_204_n2141), .A2(DP_mult_204_n1649), 
        .B1(DP_mult_204_n1648), .B2(DP_mult_204_n2042), .ZN(DP_mult_204_n1354)
         );
  OAI22_X1 DP_mult_204_U2044 ( .A1(DP_mult_204_n2319), .A2(DP_mult_204_n1770), 
        .B1(DP_mult_204_n1769), .B2(DP_mult_204_n1929), .ZN(DP_mult_204_n1471)
         );
  NOR2_X1 DP_mult_204_U2043 ( .A1(DP_mult_204_n2338), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1409) );
  INV_X1 DP_mult_204_U2042 ( .A(DP_mult_204_n1532), .ZN(DP_mult_204_n2393) );
  INV_X1 DP_mult_204_U2041 ( .A(DP_mult_204_n1632), .ZN(DP_mult_204_n2389) );
  INV_X1 DP_mult_204_U2040 ( .A(DP_mult_204_n692), .ZN(DP_mult_204_n693) );
  NOR2_X1 DP_mult_204_U2039 ( .A1(DP_mult_204_n1181), .A2(DP_mult_204_n1192), 
        .ZN(DP_mult_204_n644) );
  NAND2_X1 DP_mult_204_U2038 ( .A1(DP_mult_204_n1181), .A2(DP_mult_204_n1192), 
        .ZN(DP_mult_204_n645) );
  NAND2_X1 DP_mult_204_U2037 ( .A1(DP_mult_204_n2378), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1531) );
  NAND2_X1 DP_mult_204_U2036 ( .A1(DP_mult_204_n2356), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1681) );
  NAND2_X1 DP_mult_204_U2035 ( .A1(DP_mult_204_n2363), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1631) );
  NAND2_X1 DP_mult_204_U2034 ( .A1(DP_mult_204_n2353), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1706) );
  NAND2_X1 DP_mult_204_U2033 ( .A1(DP_mult_204_n2369), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1581) );
  NAND2_X1 DP_mult_204_U2032 ( .A1(DP_mult_204_n2359), .A2(DP_mult_204_n2384), 
        .ZN(DP_mult_204_n1656) );
  NAND2_X1 DP_mult_204_U2031 ( .A1(DP_mult_204_n2367), .A2(DP_mult_204_n2384), 
        .ZN(DP_mult_204_n1606) );
  NAND2_X1 DP_mult_204_U2030 ( .A1(DP_mult_204_n2381), .A2(DP_mult_204_n2384), 
        .ZN(DP_mult_204_n1506) );
  NAND2_X1 DP_mult_204_U2029 ( .A1(DP_mult_204_n2374), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1556) );
  INV_X1 DP_mult_204_U2028 ( .A(DP_mult_204_n2034), .ZN(DP_mult_204_n2376) );
  OAI22_X1 DP_mult_204_U2027 ( .A1(DP_mult_204_n2141), .A2(DP_mult_204_n1652), 
        .B1(DP_mult_204_n2042), .B2(DP_mult_204_n1651), .ZN(DP_mult_204_n1357)
         );
  INV_X1 DP_mult_204_U2026 ( .A(DP_mult_204_n2246), .ZN(DP_mult_204_n2324) );
  INV_X1 DP_mult_204_U2025 ( .A(DP_mult_204_n2071), .ZN(DP_mult_204_n2326) );
  INV_X1 DP_mult_204_U2024 ( .A(DP_mult_204_n1943), .ZN(DP_mult_204_n2331) );
  INV_X1 DP_mult_204_U2023 ( .A(DP_mult_204_n2063), .ZN(DP_mult_204_n2321) );
  OAI22_X1 DP_mult_204_U2022 ( .A1(DP_mult_204_n2309), .A2(DP_mult_204_n1644), 
        .B1(DP_mult_204_n2334), .B2(DP_mult_204_n1643), .ZN(DP_mult_204_n1349)
         );
  OAI22_X1 DP_mult_204_U2021 ( .A1(DP_mult_204_n2320), .A2(DP_mult_204_n1773), 
        .B1(DP_mult_204_n1772), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1474)
         );
  NOR2_X1 DP_mult_204_U2020 ( .A1(DP_mult_204_n2069), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1385) );
  OAI22_X1 DP_mult_204_U2019 ( .A1(DP_mult_204_n2320), .A2(DP_mult_204_n1777), 
        .B1(DP_mult_204_n1776), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1478)
         );
  NAND2_X1 DP_mult_204_U2018 ( .A1(DP_mult_204_n2351), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1731) );
  INV_X1 DP_mult_204_U2017 ( .A(DP_mult_204_n682), .ZN(DP_mult_204_n683) );
  INV_X1 DP_mult_204_U2016 ( .A(DP_mult_204_n1507), .ZN(DP_mult_204_n2394) );
  OAI21_X1 DP_mult_204_U2015 ( .B1(DP_mult_204_n2301), .B2(DP_mult_204_n2019), 
        .A(DP_mult_204_n2394), .ZN(DP_mult_204_n1218) );
  INV_X2 DP_mult_204_U2014 ( .A(DP_mult_204_n2383), .ZN(DP_mult_204_n2382) );
  NOR2_X1 DP_mult_204_U2013 ( .A1(DP_mult_204_n2342), .A2(DP_mult_204_n1955), 
        .ZN(DP_mult_204_n1457) );
  INV_X1 DP_mult_204_U2012 ( .A(DP_mult_204_n1682), .ZN(DP_mult_204_n2387) );
  NOR2_X1 DP_mult_204_U2011 ( .A1(DP_mult_204_n2340), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1433) );
  INV_X1 DP_mult_204_U2010 ( .A(DP_mult_204_n2365), .ZN(DP_mult_204_n2363) );
  OAI22_X1 DP_mult_204_U2009 ( .A1(DP_mult_204_n2320), .A2(DP_mult_204_n1779), 
        .B1(DP_mult_204_n1778), .B2(DP_mult_204_n251), .ZN(DP_mult_204_n1480)
         );
  NAND2_X1 DP_mult_204_U2008 ( .A1(DP_mult_204_n2348), .A2(DP_mult_204_n1954), 
        .ZN(DP_mult_204_n1756) );
  AND2_X1 DP_mult_204_U2007 ( .A1(DP_mult_204_n1194), .A2(DP_mult_204_n676), 
        .ZN(DP_mult_204_n2240) );
  NAND2_X1 DP_mult_204_U2006 ( .A1(DP_mult_204_n1175), .A2(DP_mult_204_n1178), 
        .ZN(DP_mult_204_n637) );
  NAND2_X1 DP_mult_204_U2005 ( .A1(DP_mult_204_n1159), .A2(DP_mult_204_n1161), 
        .ZN(DP_mult_204_n627) );
  NOR2_X1 DP_mult_204_U2004 ( .A1(DP_mult_204_n1175), .A2(DP_mult_204_n1178), 
        .ZN(DP_mult_204_n636) );
  NAND2_X1 DP_mult_204_U2003 ( .A1(DP_mult_204_n679), .A2(DP_mult_204_n680), 
        .ZN(DP_mult_204_n341) );
  NAND2_X1 DP_mult_204_U2002 ( .A1(DP_mult_204_n681), .A2(DP_mult_204_n684), 
        .ZN(DP_mult_204_n352) );
  NOR2_X1 DP_mult_204_U2001 ( .A1(DP_mult_204_n1159), .A2(DP_mult_204_n1161), 
        .ZN(DP_mult_204_n626) );
  OR2_X1 DP_mult_204_U2000 ( .A1(DP_mult_204_n679), .A2(DP_mult_204_n680), 
        .ZN(DP_mult_204_n2239) );
  OR2_X1 DP_mult_204_U1999 ( .A1(DP_mult_204_n681), .A2(DP_mult_204_n684), 
        .ZN(DP_mult_204_n2238) );
  OAI21_X1 DP_mult_204_U1998 ( .B1(DP_mult_204_n646), .B2(DP_mult_204_n644), 
        .A(DP_mult_204_n645), .ZN(DP_mult_204_n643) );
  AOI21_X1 DP_mult_204_U1997 ( .B1(DP_mult_204_n643), .B2(DP_mult_204_n1983), 
        .A(DP_mult_204_n1992), .ZN(DP_mult_204_n638) );
  NOR2_X1 DP_mult_204_U1996 ( .A1(DP_mult_204_n678), .A2(DP_mult_204_n677), 
        .ZN(DP_mult_204_n334) );
  AOI21_X1 DP_mult_204_U1995 ( .B1(DP_mult_204_n1982), .B2(DP_mult_204_n1981), 
        .A(DP_mult_204_n1991), .ZN(DP_mult_204_n646) );
  OR2_X1 DP_mult_204_U1994 ( .A1(DP_mult_204_n685), .A2(DP_mult_204_n688), 
        .ZN(DP_mult_204_n2237) );
  INV_X1 DP_mult_204_U1993 ( .A(DP_mult_204_n341), .ZN(DP_mult_204_n339) );
  NAND2_X1 DP_mult_204_U1992 ( .A1(DP_mult_204_n678), .A2(DP_mult_204_n677), 
        .ZN(DP_mult_204_n335) );
  INV_X1 DP_mult_204_U1991 ( .A(DP_mult_204_n676), .ZN(DP_mult_204_n677) );
  NOR2_X1 DP_mult_204_U1990 ( .A1(DP_mult_204_n1165), .A2(DP_mult_204_n1170), 
        .ZN(DP_mult_204_n631) );
  NAND2_X1 DP_mult_204_U1989 ( .A1(DP_mult_204_n2238), .A2(DP_mult_204_n352), 
        .ZN(DP_mult_204_n303) );
  NAND2_X1 DP_mult_204_U1988 ( .A1(DP_mult_204_n2239), .A2(DP_mult_204_n341), 
        .ZN(DP_mult_204_n302) );
  NAND2_X1 DP_mult_204_U1987 ( .A1(DP_mult_204_n1003), .A2(DP_mult_204_n1020), 
        .ZN(DP_mult_204_n570) );
  NAND2_X1 DP_mult_204_U1986 ( .A1(DP_mult_204_n2237), .A2(DP_mult_204_n369), 
        .ZN(DP_mult_204_n304) );
  NAND2_X1 DP_mult_204_U1985 ( .A1(DP_mult_204_n1099), .A2(DP_mult_204_n1110), 
        .ZN(DP_mult_204_n598) );
  NOR2_X1 DP_mult_204_U1984 ( .A1(DP_mult_204_n590), .A2(DP_mult_204_n592), 
        .ZN(DP_mult_204_n588) );
  OR2_X1 DP_mult_204_U1983 ( .A1(DP_mult_204_n1123), .A2(DP_mult_204_n1132), 
        .ZN(DP_mult_204_n2236) );
  NAND2_X1 DP_mult_204_U1982 ( .A1(DP_mult_204_n2222), .A2(DP_mult_204_n2232), 
        .ZN(DP_mult_204_n610) );
  INV_X1 DP_mult_204_U1981 ( .A(DP_mult_204_n369), .ZN(DP_mult_204_n367) );
  NOR2_X1 DP_mult_204_U1980 ( .A1(DP_mult_204_n336), .A2(DP_mult_204_n334), 
        .ZN(DP_mult_204_n332) );
  OR2_X1 DP_mult_204_U1979 ( .A1(DP_mult_204_n717), .A2(DP_mult_204_n726), 
        .ZN(DP_mult_204_n2235) );
  OR2_X1 DP_mult_204_U1978 ( .A1(DP_mult_204_n694), .A2(DP_mult_204_n689), 
        .ZN(DP_mult_204_n2234) );
  NAND2_X1 DP_mult_204_U1977 ( .A1(DP_mult_204_n701), .A2(DP_mult_204_n708), 
        .ZN(DP_mult_204_n396) );
  AOI21_X1 DP_mult_204_U1976 ( .B1(DP_mult_204_n376), .B2(DP_mult_204_n2237), 
        .A(DP_mult_204_n367), .ZN(DP_mult_204_n365) );
  OAI21_X1 DP_mult_204_U1975 ( .B1(DP_mult_204_n364), .B2(DP_mult_204_n387), 
        .A(DP_mult_204_n365), .ZN(DP_mult_204_n363) );
  AOI21_X1 DP_mult_204_U1974 ( .B1(DP_mult_204_n362), .B2(DP_mult_204_n394), 
        .A(DP_mult_204_n363), .ZN(DP_mult_204_n361) );
  OAI21_X1 DP_mult_204_U1973 ( .B1(DP_mult_204_n405), .B2(DP_mult_204_n360), 
        .A(DP_mult_204_n361), .ZN(DP_mult_204_n359) );
  AOI21_X1 DP_mult_204_U1972 ( .B1(DP_mult_204_n2232), .B2(DP_mult_204_n1984), 
        .A(DP_mult_204_n1993), .ZN(DP_mult_204_n611) );
  NAND2_X1 DP_mult_204_U1971 ( .A1(DP_mult_204_n695), .A2(DP_mult_204_n700), 
        .ZN(DP_mult_204_n387) );
  OR2_X1 DP_mult_204_U1970 ( .A1(DP_mult_204_n1111), .A2(DP_mult_204_n1122), 
        .ZN(DP_mult_204_n2233) );
  OR2_X1 DP_mult_204_U1969 ( .A1(DP_mult_204_n1133), .A2(DP_mult_204_n1142), 
        .ZN(DP_mult_204_n2232) );
  NOR2_X1 DP_mult_204_U1968 ( .A1(DP_mult_204_n1099), .A2(DP_mult_204_n1110), 
        .ZN(DP_mult_204_n597) );
  NAND3_X1 DP_mult_204_U1967 ( .A1(DP_mult_204_n2295), .A2(DP_mult_204_n2296), 
        .A3(DP_mult_204_n2297), .ZN(DP_mult_204_n804) );
  NAND2_X1 DP_mult_204_U1966 ( .A1(DP_mult_204_n727), .A2(DP_mult_204_n736), 
        .ZN(DP_mult_204_n429) );
  NAND2_X1 DP_mult_204_U1965 ( .A1(DP_mult_204_n2234), .A2(DP_mult_204_n2237), 
        .ZN(DP_mult_204_n364) );
  NOR2_X1 DP_mult_204_U1964 ( .A1(DP_mult_204_n633), .A2(DP_mult_204_n631), 
        .ZN(DP_mult_204_n629) );
  AOI21_X1 DP_mult_204_U1963 ( .B1(DP_mult_204_n629), .B2(DP_mult_204_n635), 
        .A(DP_mult_204_n630), .ZN(DP_mult_204_n628) );
  OR2_X1 DP_mult_204_U1962 ( .A1(DP_mult_204_n709), .A2(DP_mult_204_n716), 
        .ZN(DP_mult_204_n2231) );
  OR2_X1 DP_mult_204_U1961 ( .A1(DP_mult_204_n701), .A2(DP_mult_204_n708), 
        .ZN(DP_mult_204_n2230) );
  NOR2_X1 DP_mult_204_U1960 ( .A1(DP_mult_204_n695), .A2(DP_mult_204_n700), 
        .ZN(DP_mult_204_n384) );
  OAI21_X1 DP_mult_204_U1959 ( .B1(DP_mult_204_n628), .B2(DP_mult_204_n626), 
        .A(DP_mult_204_n627), .ZN(DP_mult_204_n625) );
  AOI21_X1 DP_mult_204_U1958 ( .B1(DP_mult_204_n625), .B2(DP_mult_204_n1995), 
        .A(DP_mult_204_n1986), .ZN(DP_mult_204_n620) );
  INV_X1 DP_mult_204_U1957 ( .A(DP_mult_204_n352), .ZN(DP_mult_204_n350) );
  NOR2_X1 DP_mult_204_U1956 ( .A1(DP_mult_204_n727), .A2(DP_mult_204_n736), 
        .ZN(DP_mult_204_n428) );
  NAND2_X1 DP_mult_204_U1955 ( .A1(DP_mult_204_n2230), .A2(DP_mult_204_n396), 
        .ZN(DP_mult_204_n307) );
  INV_X1 DP_mult_204_U1954 ( .A(DP_mult_204_n384), .ZN(DP_mult_204_n657) );
  NAND2_X1 DP_mult_204_U1953 ( .A1(DP_mult_204_n657), .A2(DP_mult_204_n387), 
        .ZN(DP_mult_204_n306) );
  NAND2_X1 DP_mult_204_U1952 ( .A1(DP_mult_204_n2231), .A2(DP_mult_204_n409), 
        .ZN(DP_mult_204_n308) );
  OR2_X1 DP_mult_204_U1951 ( .A1(DP_mult_204_n1039), .A2(DP_mult_204_n1054), 
        .ZN(DP_mult_204_n2229) );
  OR2_X1 DP_mult_204_U1950 ( .A1(DP_mult_204_n1021), .A2(DP_mult_204_n1038), 
        .ZN(DP_mult_204_n2228) );
  NAND2_X1 DP_mult_204_U1949 ( .A1(DP_mult_204_n362), .A2(DP_mult_204_n2230), 
        .ZN(DP_mult_204_n360) );
  OR2_X1 DP_mult_204_U1948 ( .A1(DP_mult_204_n1055), .A2(DP_mult_204_n1070), 
        .ZN(DP_mult_204_n2227) );
  INV_X1 DP_mult_204_U1947 ( .A(DP_mult_204_n502), .ZN(DP_mult_204_n668) );
  INV_X1 DP_mult_204_U1946 ( .A(DP_mult_204_n378), .ZN(DP_mult_204_n376) );
  INV_X1 DP_mult_204_U1945 ( .A(DP_mult_204_n428), .ZN(DP_mult_204_n661) );
  NAND2_X1 DP_mult_204_U1944 ( .A1(DP_mult_204_n661), .A2(DP_mult_204_n429), 
        .ZN(DP_mult_204_n310) );
  INV_X1 DP_mult_204_U1943 ( .A(DP_mult_204_n396), .ZN(DP_mult_204_n394) );
  INV_X1 DP_mult_204_U1942 ( .A(DP_mult_204_n418), .ZN(DP_mult_204_n416) );
  NAND2_X1 DP_mult_204_U1941 ( .A1(DP_mult_204_n2235), .A2(DP_mult_204_n2231), 
        .ZN(DP_mult_204_n402) );
  NAND2_X1 DP_mult_204_U1940 ( .A1(DP_mult_204_n789), .A2(DP_mult_204_n804), 
        .ZN(DP_mult_204_n481) );
  INV_X1 DP_mult_204_U1939 ( .A(DP_mult_204_n563), .ZN(DP_mult_204_n561) );
  INV_X1 DP_mult_204_U1938 ( .A(DP_mult_204_n564), .ZN(DP_mult_204_n562) );
  AOI21_X1 DP_mult_204_U1937 ( .B1(DP_mult_204_n565), .B2(DP_mult_204_n561), 
        .A(DP_mult_204_n562), .ZN(DP_mult_204_n560) );
  NOR2_X1 DP_mult_204_U1936 ( .A1(DP_mult_204_n435), .A2(DP_mult_204_n428), 
        .ZN(DP_mult_204_n426) );
  AND2_X1 DP_mult_204_U1935 ( .A1(DP_mult_204_n1055), .A2(DP_mult_204_n1070), 
        .ZN(DP_mult_204_n2224) );
  NOR2_X1 DP_mult_204_U1934 ( .A1(DP_mult_204_n563), .A2(DP_mult_204_n558), 
        .ZN(DP_mult_204_n552) );
  NAND2_X1 DP_mult_204_U1933 ( .A1(DP_mult_204_n897), .A2(DP_mult_204_n918), 
        .ZN(DP_mult_204_n535) );
  NOR2_X1 DP_mult_204_U1932 ( .A1(DP_mult_204_n384), .A2(DP_mult_204_n364), 
        .ZN(DP_mult_204_n362) );
  AND2_X1 DP_mult_204_U1931 ( .A1(DP_mult_204_n1021), .A2(DP_mult_204_n1038), 
        .ZN(DP_mult_204_n2223) );
  INV_X1 DP_mult_204_U1930 ( .A(DP_mult_204_n409), .ZN(DP_mult_204_n407) );
  AOI21_X1 DP_mult_204_U1929 ( .B1(DP_mult_204_n2231), .B2(DP_mult_204_n416), 
        .A(DP_mult_204_n407), .ZN(DP_mult_204_n405) );
  OAI21_X1 DP_mult_204_U1928 ( .B1(DP_mult_204_n428), .B2(DP_mult_204_n436), 
        .A(DP_mult_204_n429), .ZN(DP_mult_204_n427) );
  AOI21_X1 DP_mult_204_U1927 ( .B1(DP_mult_204_n426), .B2(DP_mult_204_n445), 
        .A(DP_mult_204_n427), .ZN(DP_mult_204_n421) );
  NAND2_X1 DP_mult_204_U1926 ( .A1(DP_mult_204_n737), .A2(DP_mult_204_n748), 
        .ZN(DP_mult_204_n436) );
  NOR2_X1 DP_mult_204_U1925 ( .A1(DP_mult_204_n805), .A2(DP_mult_204_n820), 
        .ZN(DP_mult_204_n495) );
  NOR2_X1 DP_mult_204_U1924 ( .A1(DP_mult_204_n1071), .A2(DP_mult_204_n1084), 
        .ZN(DP_mult_204_n590) );
  NOR2_X1 DP_mult_204_U1923 ( .A1(DP_mult_204_n877), .A2(DP_mult_204_n896), 
        .ZN(DP_mult_204_n531) );
  NOR2_X1 DP_mult_204_U1922 ( .A1(DP_mult_204_n737), .A2(DP_mult_204_n748), 
        .ZN(DP_mult_204_n435) );
  INV_X1 DP_mult_204_U1921 ( .A(DP_mult_204_n421), .ZN(DP_mult_204_n423) );
  NAND2_X1 DP_mult_204_U1920 ( .A1(DP_mult_204_n662), .A2(DP_mult_204_n436), 
        .ZN(DP_mult_204_n311) );
  NAND2_X1 DP_mult_204_U1919 ( .A1(DP_mult_204_n426), .A2(DP_mult_204_n663), 
        .ZN(DP_mult_204_n420) );
  INV_X1 DP_mult_204_U1918 ( .A(DP_mult_204_n439), .ZN(DP_mult_204_n445) );
  INV_X1 DP_mult_204_U1917 ( .A(DP_mult_204_n2142), .ZN(DP_mult_204_n565) );
  INV_X1 DP_mult_204_U1916 ( .A(DP_mult_204_n438), .ZN(DP_mult_204_n663) );
  NOR2_X1 DP_mult_204_U1915 ( .A1(DP_mult_204_n402), .A2(DP_mult_204_n360), 
        .ZN(DP_mult_204_n356) );
  INV_X1 DP_mult_204_U1914 ( .A(DP_mult_204_n461), .ZN(DP_mult_204_n459) );
  INV_X1 DP_mult_204_U1913 ( .A(DP_mult_204_n481), .ZN(DP_mult_204_n483) );
  INV_X1 DP_mult_204_U1912 ( .A(DP_mult_204_n436), .ZN(DP_mult_204_n434) );
  AOI21_X1 DP_mult_204_U1911 ( .B1(DP_mult_204_n662), .B2(DP_mult_204_n445), 
        .A(DP_mult_204_n434), .ZN(DP_mult_204_n432) );
  NAND2_X1 DP_mult_204_U1910 ( .A1(DP_mult_204_n663), .A2(DP_mult_204_n662), 
        .ZN(DP_mult_204_n431) );
  INV_X1 DP_mult_204_U1909 ( .A(DP_mult_204_n435), .ZN(DP_mult_204_n662) );
  INV_X1 DP_mult_204_U1908 ( .A(DP_mult_204_n2247), .ZN(DP_mult_204_n536) );
  INV_X1 DP_mult_204_U1907 ( .A(DP_mult_204_n420), .ZN(DP_mult_204_n422) );
  NOR2_X1 DP_mult_204_U1906 ( .A1(DP_mult_204_n2147), .A2(DP_mult_204_n467), 
        .ZN(DP_mult_204_n465) );
  INV_X2 DP_mult_204_U1905 ( .A(DP_mult_204_n1946), .ZN(DP_mult_204_n2314) );
  OR2_X1 DP_mult_204_U1904 ( .A1(DP_mult_204_n1143), .A2(DP_mult_204_n1150), 
        .ZN(DP_mult_204_n2222) );
  INV_X1 DP_mult_204_U1903 ( .A(DP_mult_204_n2372), .ZN(DP_mult_204_n2369) );
  INV_X1 DP_mult_204_U1902 ( .A(DP_mult_204_n2256), .ZN(DP_mult_204_n2220) );
  INV_X1 DP_mult_204_U1901 ( .A(DP_mult_204_n2250), .ZN(DP_mult_204_n2330) );
  OR2_X1 DP_mult_204_U1900 ( .A1(DP_mult_204_n805), .A2(DP_mult_204_n820), 
        .ZN(DP_mult_204_n2217) );
  OR2_X2 DP_mult_204_U1899 ( .A1(DP_mult_204_n775), .A2(DP_mult_204_n788), 
        .ZN(DP_mult_204_n2225) );
  NAND2_X1 DP_mult_204_U1898 ( .A1(DP_mult_204_n2215), .A2(DP_mult_204_n2216), 
        .ZN(DP_mult_204_n1370) );
  OR2_X1 DP_mult_204_U1897 ( .A1(DP_mult_204_n1665), .A2(DP_mult_204_n2066), 
        .ZN(DP_mult_204_n2216) );
  OR2_X1 DP_mult_204_U1896 ( .A1(DP_mult_204_n2312), .A2(DP_mult_204_n1666), 
        .ZN(DP_mult_204_n2215) );
  NAND3_X1 DP_mult_204_U1895 ( .A1(DP_mult_204_n2212), .A2(DP_mult_204_n2213), 
        .A3(DP_mult_204_n2214), .ZN(DP_mult_204_n956) );
  NAND2_X1 DP_mult_204_U1894 ( .A1(DP_mult_204_n1459), .A2(DP_mult_204_n1436), 
        .ZN(DP_mult_204_n2214) );
  NAND2_X1 DP_mult_204_U1893 ( .A1(DP_mult_204_n1370), .A2(DP_mult_204_n1436), 
        .ZN(DP_mult_204_n2213) );
  NAND2_X1 DP_mult_204_U1892 ( .A1(DP_mult_204_n1370), .A2(DP_mult_204_n1459), 
        .ZN(DP_mult_204_n2212) );
  XOR2_X1 DP_mult_204_U1891 ( .A(DP_mult_204_n1370), .B(DP_mult_204_n2211), 
        .Z(DP_mult_204_n957) );
  XOR2_X1 DP_mult_204_U1890 ( .A(DP_mult_204_n1436), .B(DP_mult_204_n1459), 
        .Z(DP_mult_204_n2211) );
  BUF_X2 DP_mult_204_U1889 ( .A(DP_mult_204_n297), .Z(DP_mult_204_n2289) );
  INV_X1 DP_mult_204_U1888 ( .A(DP_coeffs_fb_int[12]), .ZN(DP_mult_204_n2210)
         );
  INV_X1 DP_mult_204_U1887 ( .A(DP_mult_204_n508), .ZN(DP_mult_204_n2208) );
  INV_X1 DP_mult_204_U1886 ( .A(DP_coeffs_fb_int[14]), .ZN(DP_mult_204_n2207)
         );
  CLKBUF_X1 DP_mult_204_U1885 ( .A(DP_mult_204_n2043), .Z(DP_mult_204_n2205)
         );
  OR2_X1 DP_mult_204_U1884 ( .A1(DP_mult_204_n2062), .A2(DP_mult_204_n856), 
        .ZN(DP_mult_204_n2204) );
  INV_X2 DP_mult_204_U1883 ( .A(DP_mult_204_n1987), .ZN(DP_mult_204_n2209) );
  NOR2_X1 DP_mult_204_U1882 ( .A1(DP_mult_204_n839), .A2(DP_mult_204_n856), 
        .ZN(DP_mult_204_n513) );
  INV_X1 DP_mult_204_U1881 ( .A(DP_coeffs_fb_int[16]), .ZN(DP_mult_204_n2203)
         );
  INV_X1 DP_mult_204_U1880 ( .A(DP_coeffs_fb_int[6]), .ZN(DP_mult_204_n2202)
         );
  INV_X1 DP_mult_204_U1879 ( .A(DP_mult_204_n519), .ZN(DP_mult_204_n2201) );
  XNOR2_X1 DP_mult_204_U1878 ( .A(DP_mult_204_n827), .B(DP_mult_204_n844), 
        .ZN(DP_mult_204_n2200) );
  XNOR2_X1 DP_mult_204_U1877 ( .A(DP_mult_204_n2200), .B(DP_mult_204_n2128), 
        .ZN(DP_mult_204_n823) );
  NAND3_X1 DP_mult_204_U1876 ( .A1(DP_mult_204_n2197), .A2(DP_mult_204_n2198), 
        .A3(DP_mult_204_n2199), .ZN(DP_mult_204_n884) );
  NAND2_X1 DP_mult_204_U1875 ( .A1(DP_mult_204_n895), .A2(DP_mult_204_n891), 
        .ZN(DP_mult_204_n2199) );
  NAND2_X1 DP_mult_204_U1874 ( .A1(DP_mult_204_n908), .A2(DP_mult_204_n891), 
        .ZN(DP_mult_204_n2198) );
  NAND2_X1 DP_mult_204_U1873 ( .A1(DP_mult_204_n908), .A2(DP_mult_204_n895), 
        .ZN(DP_mult_204_n2197) );
  XOR2_X1 DP_mult_204_U1872 ( .A(DP_mult_204_n908), .B(DP_mult_204_n2196), .Z(
        DP_mult_204_n885) );
  XOR2_X1 DP_mult_204_U1871 ( .A(DP_mult_204_n895), .B(DP_mult_204_n891), .Z(
        DP_mult_204_n2196) );
  NAND3_X1 DP_mult_204_U1870 ( .A1(DP_mult_204_n2193), .A2(DP_mult_204_n2194), 
        .A3(DP_mult_204_n2195), .ZN(DP_mult_204_n896) );
  NAND2_X1 DP_mult_204_U1869 ( .A1(DP_mult_204_n901), .A2(DP_mult_204_n899), 
        .ZN(DP_mult_204_n2195) );
  NAND2_X1 DP_mult_204_U1868 ( .A1(DP_mult_204_n920), .A2(DP_mult_204_n899), 
        .ZN(DP_mult_204_n2194) );
  NAND2_X1 DP_mult_204_U1867 ( .A1(DP_mult_204_n920), .A2(DP_mult_204_n901), 
        .ZN(DP_mult_204_n2193) );
  NAND3_X1 DP_mult_204_U1866 ( .A1(DP_mult_204_n2190), .A2(DP_mult_204_n2191), 
        .A3(DP_mult_204_n2192), .ZN(DP_mult_204_n898) );
  NAND2_X1 DP_mult_204_U1865 ( .A1(DP_mult_204_n924), .A2(DP_mult_204_n922), 
        .ZN(DP_mult_204_n2192) );
  NAND2_X1 DP_mult_204_U1864 ( .A1(DP_mult_204_n903), .A2(DP_mult_204_n922), 
        .ZN(DP_mult_204_n2191) );
  NAND2_X1 DP_mult_204_U1863 ( .A1(DP_mult_204_n903), .A2(DP_mult_204_n924), 
        .ZN(DP_mult_204_n2190) );
  XOR2_X1 DP_mult_204_U1862 ( .A(DP_mult_204_n2189), .B(DP_mult_204_n899), .Z(
        DP_mult_204_n897) );
  XOR2_X1 DP_mult_204_U1861 ( .A(DP_mult_204_n920), .B(DP_mult_204_n901), .Z(
        DP_mult_204_n2189) );
  XOR2_X1 DP_mult_204_U1860 ( .A(DP_mult_204_n2188), .B(DP_mult_204_n922), .Z(
        DP_mult_204_n899) );
  XOR2_X1 DP_mult_204_U1859 ( .A(DP_mult_204_n903), .B(DP_mult_204_n924), .Z(
        DP_mult_204_n2188) );
  NOR2_X1 DP_mult_204_U1858 ( .A1(DP_mult_204_n805), .A2(DP_mult_204_n820), 
        .ZN(DP_mult_204_n2187) );
  INV_X1 DP_mult_204_U1857 ( .A(DP_mult_204_n2299), .ZN(DP_mult_204_n2298) );
  INV_X1 DP_mult_204_U1856 ( .A(DP_mult_204_n2169), .ZN(DP_mult_204_n2186) );
  NAND3_X1 DP_mult_204_U1855 ( .A1(DP_mult_204_n2182), .A2(DP_mult_204_n2183), 
        .A3(DP_mult_204_n2184), .ZN(DP_mult_204_n1022) );
  NAND2_X1 DP_mult_204_U1854 ( .A1(DP_mult_204_n1027), .A2(DP_mult_204_n1044), 
        .ZN(DP_mult_204_n2184) );
  NAND2_X1 DP_mult_204_U1853 ( .A1(DP_mult_204_n1042), .A2(DP_mult_204_n1044), 
        .ZN(DP_mult_204_n2183) );
  NAND2_X1 DP_mult_204_U1852 ( .A1(DP_mult_204_n1042), .A2(DP_mult_204_n1972), 
        .ZN(DP_mult_204_n2182) );
  INV_X2 DP_mult_204_U1851 ( .A(DP_mult_204_n2368), .ZN(DP_mult_204_n2367) );
  NOR2_X2 DP_mult_204_U1850 ( .A1(DP_mult_204_n502), .A2(DP_mult_204_n2187), 
        .ZN(DP_mult_204_n489) );
  CLKBUF_X1 DP_mult_204_U1849 ( .A(DP_mult_204_n512), .Z(DP_mult_204_n2179) );
  INV_X1 DP_mult_204_U1848 ( .A(DP_mult_204_n2079), .ZN(DP_mult_204_n2315) );
  INV_X1 DP_mult_204_U1847 ( .A(DP_mult_204_n2079), .ZN(DP_mult_204_n2177) );
  INV_X2 DP_mult_204_U1846 ( .A(DP_mult_204_n2013), .ZN(DP_mult_204_n2304) );
  INV_X2 DP_mult_204_U1845 ( .A(DP_mult_204_n2252), .ZN(DP_mult_204_n2335) );
  XNOR2_X1 DP_mult_204_U1844 ( .A(DP_mult_204_n1415), .B(DP_mult_204_n1393), 
        .ZN(DP_mult_204_n2175) );
  XNOR2_X1 DP_mult_204_U1843 ( .A(DP_mult_204_n2175), .B(DP_mult_204_n1988), 
        .ZN(DP_mult_204_n975) );
  NAND3_X1 DP_mult_204_U1842 ( .A1(DP_mult_204_n2172), .A2(DP_mult_204_n2173), 
        .A3(DP_mult_204_n2174), .ZN(DP_mult_204_n1038) );
  NAND2_X1 DP_mult_204_U1841 ( .A1(DP_mult_204_n1056), .A2(DP_mult_204_n1043), 
        .ZN(DP_mult_204_n2174) );
  NAND2_X1 DP_mult_204_U1840 ( .A1(DP_mult_204_n1041), .A2(DP_mult_204_n1043), 
        .ZN(DP_mult_204_n2173) );
  NAND2_X1 DP_mult_204_U1839 ( .A1(DP_mult_204_n1041), .A2(DP_mult_204_n1056), 
        .ZN(DP_mult_204_n2172) );
  XOR2_X1 DP_mult_204_U1838 ( .A(DP_mult_204_n1041), .B(DP_mult_204_n2171), 
        .Z(DP_mult_204_n1039) );
  XOR2_X1 DP_mult_204_U1837 ( .A(DP_mult_204_n1056), .B(DP_mult_204_n1043), 
        .Z(DP_mult_204_n2171) );
  XNOR2_X1 DP_mult_204_U1836 ( .A(DP_mult_204_n1027), .B(DP_mult_204_n1044), 
        .ZN(DP_mult_204_n2168) );
  XNOR2_X1 DP_mult_204_U1835 ( .A(DP_mult_204_n2168), .B(DP_mult_204_n1042), 
        .ZN(DP_mult_204_n1023) );
  NAND3_X1 DP_mult_204_U1834 ( .A1(DP_mult_204_n2165), .A2(DP_mult_204_n2166), 
        .A3(DP_mult_204_n2167), .ZN(DP_mult_204_n954) );
  NAND2_X1 DP_mult_204_U1833 ( .A1(DP_mult_204_n1414), .A2(DP_mult_204_n1304), 
        .ZN(DP_mult_204_n2167) );
  NAND2_X1 DP_mult_204_U1832 ( .A1(DP_mult_204_n1282), .A2(DP_mult_204_n1304), 
        .ZN(DP_mult_204_n2166) );
  NAND2_X1 DP_mult_204_U1831 ( .A1(DP_mult_204_n1414), .A2(DP_mult_204_n1282), 
        .ZN(DP_mult_204_n2165) );
  XOR2_X1 DP_mult_204_U1830 ( .A(DP_mult_204_n2164), .B(DP_mult_204_n1282), 
        .Z(DP_mult_204_n955) );
  XOR2_X1 DP_mult_204_U1829 ( .A(DP_mult_204_n1414), .B(DP_mult_204_n1304), 
        .Z(DP_mult_204_n2164) );
  NOR2_X1 DP_mult_204_U1828 ( .A1(DP_mult_204_n856), .A2(DP_mult_204_n839), 
        .ZN(DP_mult_204_n2163) );
  NAND3_X1 DP_mult_204_U1827 ( .A1(DP_mult_204_n2258), .A2(DP_mult_204_n2259), 
        .A3(DP_mult_204_n2260), .ZN(DP_mult_204_n2162) );
  XNOR2_X1 DP_mult_204_U1826 ( .A(DP_mult_204_n996), .B(DP_mult_204_n1217), 
        .ZN(DP_mult_204_n2161) );
  XNOR2_X1 DP_mult_204_U1825 ( .A(DP_mult_204_n2058), .B(DP_mult_204_n2161), 
        .ZN(DP_mult_204_n973) );
  NOR2_X1 DP_mult_204_U1824 ( .A1(DP_mult_204_n941), .A2(DP_mult_204_n962), 
        .ZN(DP_mult_204_n547) );
  NAND3_X1 DP_mult_204_U1823 ( .A1(DP_mult_204_n2158), .A2(DP_mult_204_n2159), 
        .A3(DP_mult_204_n2160), .ZN(DP_mult_204_n940) );
  NAND2_X1 DP_mult_204_U1822 ( .A1(DP_mult_204_n964), .A2(DP_mult_204_n945), 
        .ZN(DP_mult_204_n2160) );
  NAND2_X1 DP_mult_204_U1821 ( .A1(DP_mult_204_n943), .A2(DP_mult_204_n945), 
        .ZN(DP_mult_204_n2159) );
  NAND2_X1 DP_mult_204_U1820 ( .A1(DP_mult_204_n943), .A2(DP_mult_204_n964), 
        .ZN(DP_mult_204_n2158) );
  XOR2_X1 DP_mult_204_U1819 ( .A(DP_mult_204_n943), .B(DP_mult_204_n2157), .Z(
        DP_mult_204_n941) );
  XOR2_X1 DP_mult_204_U1818 ( .A(DP_mult_204_n964), .B(DP_mult_204_n945), .Z(
        DP_mult_204_n2157) );
  BUF_X1 DP_mult_204_U1817 ( .A(DP_mult_204_n547), .Z(DP_mult_204_n2156) );
  INV_X1 DP_mult_204_U1816 ( .A(DP_mult_204_n2246), .ZN(DP_mult_204_n2323) );
  INV_X2 DP_mult_204_U1815 ( .A(DP_mult_204_n2060), .ZN(DP_mult_204_n2342) );
  XNOR2_X1 DP_mult_204_U1814 ( .A(DP_coeffs_fb_int[1]), .B(DP_mult_204_n2383), 
        .ZN(DP_mult_204_n1806) );
  OAI22_X1 DP_mult_204_U1813 ( .A1(DP_mult_204_n2209), .A2(DP_mult_204_n1658), 
        .B1(DP_mult_204_n1657), .B2(DP_mult_204_n2066), .ZN(DP_mult_204_n2154)
         );
  INV_X2 DP_mult_204_U1812 ( .A(DP_mult_204_n2372), .ZN(DP_mult_204_n2370) );
  NAND3_X1 DP_mult_204_U1811 ( .A1(DP_mult_204_n2151), .A2(DP_mult_204_n2152), 
        .A3(DP_mult_204_n2153), .ZN(DP_mult_204_n922) );
  NAND2_X1 DP_mult_204_U1810 ( .A1(DP_mult_204_n948), .A2(DP_mult_204_n929), 
        .ZN(DP_mult_204_n2153) );
  NAND2_X1 DP_mult_204_U1809 ( .A1(DP_mult_204_n946), .A2(DP_mult_204_n929), 
        .ZN(DP_mult_204_n2152) );
  NAND2_X1 DP_mult_204_U1808 ( .A1(DP_mult_204_n946), .A2(DP_mult_204_n948), 
        .ZN(DP_mult_204_n2151) );
  XOR2_X1 DP_mult_204_U1807 ( .A(DP_mult_204_n946), .B(DP_mult_204_n2150), .Z(
        DP_mult_204_n923) );
  XOR2_X1 DP_mult_204_U1806 ( .A(DP_mult_204_n948), .B(DP_mult_204_n929), .Z(
        DP_mult_204_n2150) );
  AND2_X1 DP_mult_204_U1805 ( .A1(DP_mult_204_n821), .A2(DP_mult_204_n838), 
        .ZN(DP_mult_204_n2149) );
  INV_X1 DP_mult_204_U1804 ( .A(DP_coeffs_fb_int[2]), .ZN(DP_mult_204_n2380)
         );
  XNOR2_X1 DP_mult_204_U1803 ( .A(DP_coeffs_fb_int[3]), .B(DP_mult_204_n2380), 
        .ZN(DP_mult_204_n1807) );
  INV_X1 DP_mult_204_U1802 ( .A(DP_mult_204_n2245), .ZN(DP_mult_204_n2339) );
  INV_X2 DP_mult_204_U1801 ( .A(DP_mult_204_n2352), .ZN(DP_mult_204_n2351) );
  INV_X2 DP_mult_204_U1800 ( .A(DP_mult_204_n2375), .ZN(DP_mult_204_n2374) );
  OR2_X1 DP_mult_204_U1799 ( .A1(DP_mult_204_n502), .A2(DP_mult_204_n2187), 
        .ZN(DP_mult_204_n2147) );
  AOI21_X1 DP_mult_204_U1798 ( .B1(DP_mult_204_n581), .B2(DP_mult_204_n567), 
        .A(DP_mult_204_n568), .ZN(DP_mult_204_n566) );
  NOR2_X1 DP_mult_204_U1797 ( .A1(DP_mult_204_n963), .A2(DP_mult_204_n982), 
        .ZN(DP_mult_204_n558) );
  OR2_X1 DP_mult_204_U1796 ( .A1(DP_mult_204_n982), .A2(DP_mult_204_n963), 
        .ZN(DP_mult_204_n2146) );
  INV_X1 DP_mult_204_U1795 ( .A(DP_mult_204_n2242), .ZN(DP_mult_204_n2319) );
  BUF_X2 DP_mult_204_U1794 ( .A(DP_mult_204_n285), .Z(DP_mult_204_n2206) );
  INV_X2 DP_mult_204_U1793 ( .A(DP_mult_204_n2145), .ZN(DP_mult_204_n2334) );
  INV_X1 DP_mult_204_U1792 ( .A(DP_mult_204_n2310), .ZN(DP_mult_204_n2309) );
  NAND2_X1 DP_mult_204_U1791 ( .A1(DP_mult_204_n2143), .A2(DP_mult_204_n2144), 
        .ZN(DP_mult_204_n1352) );
  OR2_X1 DP_mult_204_U1790 ( .A1(DP_mult_204_n1646), .A2(DP_mult_204_n2334), 
        .ZN(DP_mult_204_n2144) );
  OR2_X1 DP_mult_204_U1789 ( .A1(DP_mult_204_n2309), .A2(DP_mult_204_n1647), 
        .ZN(DP_mult_204_n2143) );
  AOI21_X1 DP_mult_204_U1788 ( .B1(DP_mult_204_n2023), .B2(DP_mult_204_n567), 
        .A(DP_mult_204_n2117), .ZN(DP_mult_204_n2142) );
  INV_X1 DP_mult_204_U1787 ( .A(DP_mult_204_n2310), .ZN(DP_mult_204_n2140) );
  INV_X1 DP_mult_204_U1786 ( .A(DP_mult_204_n2310), .ZN(DP_mult_204_n2141) );
  NAND3_X1 DP_mult_204_U1785 ( .A1(DP_mult_204_n2138), .A2(DP_mult_204_n2139), 
        .A3(DP_mult_204_n2137), .ZN(DP_mult_204_n834) );
  NAND2_X1 DP_mult_204_U1784 ( .A1(DP_mult_204_n1276), .A2(DP_mult_204_n1210), 
        .ZN(DP_mult_204_n2139) );
  NAND2_X1 DP_mult_204_U1783 ( .A1(DP_mult_204_n837), .A2(DP_mult_204_n1210), 
        .ZN(DP_mult_204_n2138) );
  NAND2_X1 DP_mult_204_U1782 ( .A1(DP_mult_204_n837), .A2(DP_mult_204_n1276), 
        .ZN(DP_mult_204_n2137) );
  OAI22_X1 DP_mult_204_U1781 ( .A1(DP_mult_204_n1733), .A2(DP_mult_204_n2317), 
        .B1(DP_mult_204_n1732), .B2(DP_mult_204_n2155), .ZN(DP_mult_204_n2136)
         );
  INV_X1 DP_mult_204_U1780 ( .A(DP_mult_204_n2361), .ZN(DP_mult_204_n2134) );
  INV_X1 DP_mult_204_U1779 ( .A(DP_mult_204_n2361), .ZN(DP_mult_204_n2135) );
  NAND3_X1 DP_mult_204_U1778 ( .A1(DP_mult_204_n2131), .A2(DP_mult_204_n2132), 
        .A3(DP_mult_204_n2133), .ZN(DP_mult_204_n806) );
  NAND2_X1 DP_mult_204_U1777 ( .A1(DP_mult_204_n811), .A2(DP_mult_204_n826), 
        .ZN(DP_mult_204_n2133) );
  NAND2_X1 DP_mult_204_U1776 ( .A1(DP_mult_204_n824), .A2(DP_mult_204_n826), 
        .ZN(DP_mult_204_n2132) );
  NAND2_X1 DP_mult_204_U1775 ( .A1(DP_mult_204_n824), .A2(DP_mult_204_n811), 
        .ZN(DP_mult_204_n2131) );
  AND2_X1 DP_mult_204_U1774 ( .A1(DP_mult_204_n1816), .A2(DP_mult_204_n2155), 
        .ZN(DP_mult_204_n2130) );
  AND2_X1 DP_mult_204_U1773 ( .A1(DP_mult_204_n1816), .A2(DP_mult_204_n2155), 
        .ZN(DP_mult_204_n2129) );
  NAND3_X1 DP_mult_204_U1772 ( .A1(DP_mult_204_n2268), .A2(DP_mult_204_n2269), 
        .A3(DP_mult_204_n2270), .ZN(DP_mult_204_n2127) );
  NAND3_X1 DP_mult_204_U1771 ( .A1(DP_mult_204_n2268), .A2(DP_mult_204_n2269), 
        .A3(DP_mult_204_n2270), .ZN(DP_mult_204_n2128) );
  INV_X1 DP_mult_204_U1770 ( .A(DP_mult_204_n524), .ZN(DP_mult_204_n2126) );
  XOR2_X1 DP_mult_204_U1769 ( .A(DP_mult_204_n1238), .B(DP_mult_204_n1216), 
        .Z(DP_mult_204_n961) );
  NAND3_X1 DP_mult_204_U1768 ( .A1(DP_mult_204_n2123), .A2(DP_mult_204_n2124), 
        .A3(DP_mult_204_n2125), .ZN(DP_mult_204_n790) );
  NAND2_X1 DP_mult_204_U1767 ( .A1(DP_mult_204_n795), .A2(DP_mult_204_n810), 
        .ZN(DP_mult_204_n2125) );
  NAND2_X1 DP_mult_204_U1766 ( .A1(DP_mult_204_n808), .A2(DP_mult_204_n810), 
        .ZN(DP_mult_204_n2124) );
  NAND2_X1 DP_mult_204_U1765 ( .A1(DP_mult_204_n808), .A2(DP_mult_204_n795), 
        .ZN(DP_mult_204_n2123) );
  XOR2_X1 DP_mult_204_U1764 ( .A(DP_mult_204_n808), .B(DP_mult_204_n2122), .Z(
        DP_mult_204_n791) );
  XOR2_X1 DP_mult_204_U1763 ( .A(DP_mult_204_n795), .B(DP_mult_204_n810), .Z(
        DP_mult_204_n2122) );
  INV_X1 DP_mult_204_U1762 ( .A(DP_mult_204_n2242), .ZN(DP_mult_204_n2320) );
  INV_X1 DP_mult_204_U1761 ( .A(DP_mult_204_n2242), .ZN(DP_mult_204_n2120) );
  XNOR2_X1 DP_mult_204_U1760 ( .A(DP_mult_204_n811), .B(DP_mult_204_n826), 
        .ZN(DP_mult_204_n2119) );
  XNOR2_X1 DP_mult_204_U1759 ( .A(DP_mult_204_n824), .B(DP_mult_204_n2119), 
        .ZN(DP_mult_204_n807) );
  INV_X1 DP_mult_204_U1758 ( .A(DP_mult_204_n2176), .ZN(DP_mult_204_n2252) );
  CLKBUF_X1 DP_mult_204_U1757 ( .A(DP_mult_204_n2181), .Z(DP_mult_204_n2118)
         );
  CLKBUF_X1 DP_mult_204_U1756 ( .A(DP_mult_204_n837), .Z(DP_mult_204_n2116) );
  INV_X2 DP_mult_204_U1755 ( .A(DP_mult_204_n2005), .ZN(DP_mult_204_n2381) );
  NAND2_X1 DP_mult_204_U1754 ( .A1(DP_mult_204_n2114), .A2(DP_mult_204_n2115), 
        .ZN(DP_mult_204_n1260) );
  OR2_X1 DP_mult_204_U1753 ( .A1(DP_mult_204_n1550), .A2(DP_mult_204_n2327), 
        .ZN(DP_mult_204_n2115) );
  OR2_X1 DP_mult_204_U1752 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1551), 
        .ZN(DP_mult_204_n2114) );
  NAND3_X1 DP_mult_204_U1751 ( .A1(DP_mult_204_n2111), .A2(DP_mult_204_n2112), 
        .A3(DP_mult_204_n2113), .ZN(DP_mult_204_n958) );
  NAND2_X1 DP_mult_204_U1750 ( .A1(DP_mult_204_n1182), .A2(DP_mult_204_n1348), 
        .ZN(DP_mult_204_n2113) );
  NAND2_X1 DP_mult_204_U1749 ( .A1(DP_mult_204_n1260), .A2(DP_mult_204_n1348), 
        .ZN(DP_mult_204_n2112) );
  NAND2_X1 DP_mult_204_U1748 ( .A1(DP_mult_204_n1260), .A2(DP_mult_204_n1182), 
        .ZN(DP_mult_204_n2111) );
  XOR2_X1 DP_mult_204_U1747 ( .A(DP_mult_204_n1260), .B(DP_mult_204_n2110), 
        .Z(DP_mult_204_n959) );
  XOR2_X1 DP_mult_204_U1746 ( .A(DP_mult_204_n1182), .B(DP_mult_204_n1348), 
        .Z(DP_mult_204_n2110) );
  AND2_X1 DP_mult_204_U1745 ( .A1(DP_mult_204_n1814), .A2(DP_mult_204_n2336), 
        .ZN(DP_mult_204_n2169) );
  INV_X1 DP_mult_204_U1744 ( .A(DP_mult_204_n2001), .ZN(DP_mult_204_n2344) );
  XNOR2_X1 DP_mult_204_U1743 ( .A(DP_coeffs_fb_int[23]), .B(DP_mult_204_n2347), 
        .ZN(DP_mult_204_n1817) );
  NAND3_X1 DP_mult_204_U1742 ( .A1(DP_mult_204_n2106), .A2(DP_mult_204_n2107), 
        .A3(DP_mult_204_n2108), .ZN(DP_mult_204_n808) );
  NAND2_X1 DP_mult_204_U1741 ( .A1(DP_mult_204_n813), .A2(DP_mult_204_n819), 
        .ZN(DP_mult_204_n2108) );
  NAND2_X1 DP_mult_204_U1740 ( .A1(DP_mult_204_n828), .A2(DP_mult_204_n819), 
        .ZN(DP_mult_204_n2107) );
  NAND2_X1 DP_mult_204_U1739 ( .A1(DP_mult_204_n828), .A2(DP_mult_204_n813), 
        .ZN(DP_mult_204_n2106) );
  XOR2_X1 DP_mult_204_U1738 ( .A(DP_mult_204_n828), .B(DP_mult_204_n2105), .Z(
        DP_mult_204_n809) );
  XOR2_X1 DP_mult_204_U1737 ( .A(DP_mult_204_n813), .B(DP_mult_204_n819), .Z(
        DP_mult_204_n2105) );
  OAI22_X1 DP_mult_204_U1736 ( .A1(DP_mult_204_n2068), .A2(DP_mult_204_n1528), 
        .B1(DP_mult_204_n1527), .B2(DP_mult_204_n2325), .ZN(DP_mult_204_n1238)
         );
  INV_X1 DP_mult_204_U1735 ( .A(DP_mult_204_n2207), .ZN(DP_mult_204_n2356) );
  XNOR2_X1 DP_mult_204_U1734 ( .A(DP_coeffs_fb_int[15]), .B(DP_mult_204_n2358), 
        .ZN(DP_mult_204_n1813) );
  INV_X1 DP_mult_204_U1733 ( .A(DP_mult_204_n2243), .ZN(DP_mult_204_n2336) );
  XNOR2_X1 DP_mult_204_U1732 ( .A(DP_coeffs_fb_int[7]), .B(DP_coeffs_fb_int[8]), .ZN(DP_mult_204_n2103) );
  INV_X1 DP_mult_204_U1731 ( .A(DP_mult_204_n2016), .ZN(DP_mult_204_n2308) );
  INV_X1 DP_mult_204_U1730 ( .A(DP_mult_204_n2069), .ZN(DP_mult_204_n2102) );
  BUF_X1 DP_mult_204_U1729 ( .A(DP_mult_204_n1327), .Z(DP_mult_204_n2101) );
  NAND3_X1 DP_mult_204_U1728 ( .A1(DP_mult_204_n2098), .A2(DP_mult_204_n2099), 
        .A3(DP_mult_204_n2100), .ZN(DP_mult_204_n970) );
  NAND2_X1 DP_mult_204_U1727 ( .A1(DP_mult_204_n979), .A2(DP_mult_204_n977), 
        .ZN(DP_mult_204_n2100) );
  NAND2_X1 DP_mult_204_U1726 ( .A1(DP_mult_204_n998), .A2(DP_mult_204_n977), 
        .ZN(DP_mult_204_n2099) );
  NAND2_X1 DP_mult_204_U1725 ( .A1(DP_mult_204_n998), .A2(DP_mult_204_n979), 
        .ZN(DP_mult_204_n2098) );
  NAND3_X1 DP_mult_204_U1724 ( .A1(DP_mult_204_n2095), .A2(DP_mult_204_n2096), 
        .A3(DP_mult_204_n2097), .ZN(DP_mult_204_n976) );
  NAND2_X1 DP_mult_204_U1723 ( .A1(DP_mult_204_n1437), .A2(DP_mult_204_n1327), 
        .ZN(DP_mult_204_n2097) );
  NAND2_X1 DP_mult_204_U1722 ( .A1(DP_mult_204_n1305), .A2(DP_mult_204_n1327), 
        .ZN(DP_mult_204_n2096) );
  NAND2_X1 DP_mult_204_U1721 ( .A1(DP_mult_204_n1305), .A2(DP_mult_204_n1437), 
        .ZN(DP_mult_204_n2095) );
  XOR2_X1 DP_mult_204_U1720 ( .A(DP_mult_204_n2094), .B(DP_mult_204_n977), .Z(
        DP_mult_204_n971) );
  XOR2_X1 DP_mult_204_U1719 ( .A(DP_mult_204_n998), .B(DP_mult_204_n979), .Z(
        DP_mult_204_n2094) );
  CLKBUF_X1 DP_mult_204_U1718 ( .A(DP_mult_204_n490), .Z(DP_mult_204_n2093) );
  INV_X2 DP_mult_204_U1717 ( .A(DP_mult_204_n2375), .ZN(DP_mult_204_n2373) );
  XNOR2_X1 DP_mult_204_U1716 ( .A(DP_coeffs_fb_int[13]), .B(
        DP_coeffs_fb_int[14]), .ZN(DP_mult_204_n2181) );
  INV_X1 DP_mult_204_U1715 ( .A(DP_mult_204_n451), .ZN(DP_mult_204_n2092) );
  NAND2_X1 DP_mult_204_U1714 ( .A1(DP_mult_204_n2247), .A2(DP_mult_204_n450), 
        .ZN(DP_mult_204_n2091) );
  NAND3_X1 DP_mult_204_U1713 ( .A1(DP_mult_204_n2088), .A2(DP_mult_204_n2089), 
        .A3(DP_mult_204_n2090), .ZN(DP_mult_204_n882) );
  NAND2_X1 DP_mult_204_U1712 ( .A1(DP_mult_204_n893), .A2(DP_mult_204_n889), 
        .ZN(DP_mult_204_n2090) );
  NAND2_X1 DP_mult_204_U1711 ( .A1(DP_mult_204_n906), .A2(DP_mult_204_n889), 
        .ZN(DP_mult_204_n2089) );
  NAND2_X1 DP_mult_204_U1710 ( .A1(DP_mult_204_n906), .A2(DP_mult_204_n893), 
        .ZN(DP_mult_204_n2088) );
  XOR2_X1 DP_mult_204_U1709 ( .A(DP_mult_204_n906), .B(DP_mult_204_n2087), .Z(
        DP_mult_204_n883) );
  XOR2_X1 DP_mult_204_U1708 ( .A(DP_mult_204_n893), .B(DP_mult_204_n889), .Z(
        DP_mult_204_n2087) );
  CLKBUF_X1 DP_mult_204_U1707 ( .A(DP_mult_204_n919), .Z(DP_mult_204_n2086) );
  NAND3_X1 DP_mult_204_U1706 ( .A1(DP_mult_204_n2083), .A2(DP_mult_204_n2084), 
        .A3(DP_mult_204_n2085), .ZN(DP_mult_204_n1018) );
  NAND2_X1 DP_mult_204_U1705 ( .A1(DP_mult_204_n1263), .A2(DP_mult_204_n2035), 
        .ZN(DP_mult_204_n2085) );
  NAND2_X1 DP_mult_204_U1704 ( .A1(DP_mult_204_n2035), .A2(DP_mult_204_n1351), 
        .ZN(DP_mult_204_n2084) );
  NAND2_X1 DP_mult_204_U1703 ( .A1(DP_mult_204_n1263), .A2(DP_mult_204_n1351), 
        .ZN(DP_mult_204_n2083) );
  AND2_X1 DP_mult_204_U1702 ( .A1(DP_mult_204_n1810), .A2(DP_mult_204_n2330), 
        .ZN(DP_mult_204_n2081) );
  XNOR2_X1 DP_mult_204_U1701 ( .A(DP_coeffs_fb_int[5]), .B(DP_mult_204_n2375), 
        .ZN(DP_mult_204_n1808) );
  AND2_X1 DP_mult_204_U1700 ( .A1(DP_mult_204_n1815), .A2(DP_mult_204_n2339), 
        .ZN(DP_mult_204_n2079) );
  NAND3_X1 DP_mult_204_U1699 ( .A1(DP_mult_204_n2076), .A2(DP_mult_204_n2077), 
        .A3(DP_mult_204_n2078), .ZN(DP_mult_204_n926) );
  NAND2_X1 DP_mult_204_U1698 ( .A1(DP_mult_204_n952), .A2(DP_mult_204_n933), 
        .ZN(DP_mult_204_n2078) );
  NAND2_X1 DP_mult_204_U1697 ( .A1(DP_mult_204_n937), .A2(DP_mult_204_n933), 
        .ZN(DP_mult_204_n2077) );
  NAND2_X1 DP_mult_204_U1696 ( .A1(DP_mult_204_n937), .A2(DP_mult_204_n952), 
        .ZN(DP_mult_204_n2076) );
  NAND3_X1 DP_mult_204_U1695 ( .A1(DP_mult_204_n2073), .A2(DP_mult_204_n2074), 
        .A3(DP_mult_204_n2075), .ZN(DP_mult_204_n932) );
  NAND2_X1 DP_mult_204_U1694 ( .A1(DP_mult_204_n1413), .A2(DP_mult_204_n1325), 
        .ZN(DP_mult_204_n2075) );
  NAND2_X1 DP_mult_204_U1693 ( .A1(DP_mult_204_n1435), .A2(DP_mult_204_n1325), 
        .ZN(DP_mult_204_n2074) );
  NAND2_X1 DP_mult_204_U1692 ( .A1(DP_mult_204_n1435), .A2(DP_mult_204_n1413), 
        .ZN(DP_mult_204_n2073) );
  XOR2_X1 DP_mult_204_U1691 ( .A(DP_mult_204_n2072), .B(DP_mult_204_n933), .Z(
        DP_mult_204_n927) );
  XOR2_X1 DP_mult_204_U1690 ( .A(DP_mult_204_n937), .B(DP_mult_204_n952), .Z(
        DP_mult_204_n2072) );
  INV_X2 DP_mult_204_U1689 ( .A(DP_mult_204_n2303), .ZN(DP_mult_204_n2302) );
  XOR2_X1 DP_mult_204_U1688 ( .A(DP_coeffs_fb_int[5]), .B(DP_coeffs_fb_int[6]), 
        .Z(DP_mult_204_n2071) );
  INV_X1 DP_mult_204_U1687 ( .A(DP_mult_204_n2016), .ZN(DP_mult_204_n2070) );
  INV_X1 DP_mult_204_U1686 ( .A(DP_mult_204_n2252), .ZN(DP_mult_204_n2069) );
  XOR2_X1 DP_mult_204_U1685 ( .A(DP_mult_204_n1966), .B(DP_mult_204_n1240), 
        .Z(DP_mult_204_n1001) );
  INV_X1 DP_mult_204_U1684 ( .A(DP_mult_204_n2301), .ZN(DP_mult_204_n2300) );
  INV_X1 DP_mult_204_U1683 ( .A(DP_mult_204_n2301), .ZN(DP_mult_204_n2067) );
  INV_X1 DP_mult_204_U1682 ( .A(DP_mult_204_n2301), .ZN(DP_mult_204_n2068) );
  INV_X2 DP_mult_204_U1681 ( .A(DP_mult_204_n2129), .ZN(DP_mult_204_n2279) );
  XNOR2_X1 DP_mult_204_U1680 ( .A(DP_coeffs_fb_int[7]), .B(DP_mult_204_n2202), 
        .ZN(DP_mult_204_n1809) );
  XNOR2_X1 DP_mult_204_U1679 ( .A(DP_coeffs_fb_int[13]), .B(DP_mult_204_n2361), 
        .ZN(DP_mult_204_n1812) );
  XNOR2_X1 DP_mult_204_U1678 ( .A(DP_coeffs_fb_int[11]), .B(DP_mult_204_n2365), 
        .ZN(DP_mult_204_n1811) );
  XNOR2_X1 DP_mult_204_U1677 ( .A(DP_coeffs_fb_int[16]), .B(
        DP_coeffs_fb_int[15]), .ZN(DP_mult_204_n2176) );
  INV_X2 DP_mult_204_U1676 ( .A(DP_mult_204_n2252), .ZN(DP_mult_204_n2066) );
  XOR2_X1 DP_mult_204_U1675 ( .A(DP_coeffs_fb_int[1]), .B(DP_coeffs_fb_int[2]), 
        .Z(DP_mult_204_n2063) );
  XOR2_X1 DP_mult_204_U1674 ( .A(DP_coeffs_fb_int[1]), .B(DP_coeffs_fb_int[2]), 
        .Z(DP_mult_204_n2064) );
  CLKBUF_X1 DP_mult_204_U1673 ( .A(DP_mult_204_n839), .Z(DP_mult_204_n2062) );
  XNOR2_X1 DP_mult_204_U1672 ( .A(DP_coeffs_fb_int[11]), .B(
        DP_coeffs_fb_int[12]), .ZN(DP_mult_204_n2061) );
  INV_X1 DP_mult_204_U1671 ( .A(DP_mult_204_n2103), .ZN(DP_mult_204_n2244) );
  INV_X2 DP_mult_204_U1670 ( .A(DP_mult_204_n2244), .ZN(DP_mult_204_n2328) );
  INV_X2 DP_mult_204_U1669 ( .A(DP_mult_204_n2014), .ZN(DP_mult_204_n2305) );
  XOR2_X1 DP_mult_204_U1668 ( .A(DP_coeffs_fb_int[21]), .B(
        DP_coeffs_fb_int[22]), .Z(DP_mult_204_n2060) );
  AND2_X2 DP_mult_204_U1667 ( .A1(DP_mult_204_n1807), .A2(DP_mult_204_n2323), 
        .ZN(DP_mult_204_n2301) );
  XOR2_X1 DP_mult_204_U1666 ( .A(DP_coeffs_fb_int[17]), .B(
        DP_coeffs_fb_int[18]), .Z(DP_mult_204_n2243) );
  XNOR2_X1 DP_mult_204_U1665 ( .A(DP_mult_204_n1435), .B(DP_mult_204_n1413), 
        .ZN(DP_mult_204_n2059) );
  XNOR2_X1 DP_mult_204_U1664 ( .A(DP_mult_204_n2059), .B(DP_mult_204_n1325), 
        .ZN(DP_mult_204_n933) );
  XNOR2_X1 DP_mult_204_U1663 ( .A(DP_coeffs_fb_int[21]), .B(DP_mult_204_n2349), 
        .ZN(DP_mult_204_n1816) );
  CLKBUF_X1 DP_mult_204_U1662 ( .A(DP_mult_204_n994), .Z(DP_mult_204_n2058) );
  NAND3_X1 DP_mult_204_U1661 ( .A1(DP_mult_204_n2055), .A2(DP_mult_204_n2056), 
        .A3(DP_mult_204_n2057), .ZN(DP_mult_204_n946) );
  NAND2_X1 DP_mult_204_U1660 ( .A1(DP_mult_204_n953), .A2(DP_mult_204_n959), 
        .ZN(DP_mult_204_n2057) );
  NAND2_X1 DP_mult_204_U1659 ( .A1(DP_mult_204_n972), .A2(DP_mult_204_n959), 
        .ZN(DP_mult_204_n2056) );
  NAND2_X1 DP_mult_204_U1658 ( .A1(DP_mult_204_n972), .A2(DP_mult_204_n953), 
        .ZN(DP_mult_204_n2055) );
  INV_X2 DP_mult_204_U1657 ( .A(DP_mult_204_n2045), .ZN(DP_mult_204_n2366) );
  NAND3_X1 DP_mult_204_U1656 ( .A1(DP_mult_204_n2052), .A2(DP_mult_204_n2053), 
        .A3(DP_mult_204_n2054), .ZN(DP_mult_204_n858) );
  NAND2_X1 DP_mult_204_U1655 ( .A1(DP_mult_204_n863), .A2(DP_mult_204_n882), 
        .ZN(DP_mult_204_n2054) );
  NAND2_X1 DP_mult_204_U1654 ( .A1(DP_mult_204_n880), .A2(DP_mult_204_n882), 
        .ZN(DP_mult_204_n2053) );
  NAND2_X1 DP_mult_204_U1653 ( .A1(DP_mult_204_n880), .A2(DP_mult_204_n863), 
        .ZN(DP_mult_204_n2052) );
  INV_X2 DP_mult_204_U1652 ( .A(DP_mult_204_n2207), .ZN(DP_mult_204_n2355) );
  INV_X2 DP_mult_204_U1651 ( .A(DP_mult_204_n2082), .ZN(DP_mult_204_n2306) );
  INV_X2 DP_mult_204_U1650 ( .A(DP_mult_204_n2347), .ZN(DP_mult_204_n2346) );
  INV_X2 DP_mult_204_U1649 ( .A(DP_mult_204_n2080), .ZN(DP_mult_204_n2316) );
  NAND3_X1 DP_mult_204_U1648 ( .A1(DP_mult_204_n2049), .A2(DP_mult_204_n2050), 
        .A3(DP_mult_204_n2051), .ZN(DP_mult_204_n844) );
  NAND2_X1 DP_mult_204_U1647 ( .A1(DP_mult_204_n853), .A2(DP_mult_204_n855), 
        .ZN(DP_mult_204_n2051) );
  NAND2_X1 DP_mult_204_U1646 ( .A1(DP_mult_204_n866), .A2(DP_mult_204_n855), 
        .ZN(DP_mult_204_n2050) );
  NAND2_X1 DP_mult_204_U1645 ( .A1(DP_mult_204_n866), .A2(DP_mult_204_n853), 
        .ZN(DP_mult_204_n2049) );
  XOR2_X1 DP_mult_204_U1644 ( .A(DP_mult_204_n866), .B(DP_mult_204_n2048), .Z(
        DP_mult_204_n845) );
  XOR2_X1 DP_mult_204_U1643 ( .A(DP_mult_204_n853), .B(DP_mult_204_n855), .Z(
        DP_mult_204_n2048) );
  XNOR2_X1 DP_mult_204_U1642 ( .A(DP_mult_204_n863), .B(DP_mult_204_n882), 
        .ZN(DP_mult_204_n2047) );
  XNOR2_X1 DP_mult_204_U1641 ( .A(DP_mult_204_n880), .B(DP_mult_204_n2047), 
        .ZN(DP_mult_204_n859) );
  INV_X2 DP_mult_204_U1640 ( .A(DP_mult_204_n1947), .ZN(DP_mult_204_n2185) );
  NOR2_X1 DP_mult_204_U1639 ( .A1(DP_mult_204_n1003), .A2(DP_mult_204_n1020), 
        .ZN(DP_mult_204_n2046) );
  INV_X1 DP_mult_204_U1638 ( .A(DP_coeffs_fb_int[8]), .ZN(DP_mult_204_n2045)
         );
  XNOR2_X1 DP_mult_204_U1637 ( .A(DP_mult_204_n953), .B(DP_mult_204_n959), 
        .ZN(DP_mult_204_n2044) );
  XNOR2_X1 DP_mult_204_U1636 ( .A(DP_mult_204_n972), .B(DP_mult_204_n2044), 
        .ZN(DP_mult_204_n947) );
  NAND3_X1 DP_mult_204_U1635 ( .A1(DP_mult_204_n2137), .A2(DP_mult_204_n2138), 
        .A3(DP_mult_204_n2139), .ZN(DP_mult_204_n2043) );
  INV_X1 DP_mult_204_U1634 ( .A(DP_mult_204_n1937), .ZN(DP_mult_204_n2341) );
  INV_X1 DP_mult_204_U1633 ( .A(DP_mult_204_n1943), .ZN(DP_mult_204_n2332) );
  XOR2_X1 DP_mult_204_U1632 ( .A(DP_sw0_1_), .B(DP_mult_204_n2005), .Z(
        DP_mult_204_n1504) );
  BUF_X4 DP_mult_204_U1631 ( .A(DP_mult_204_n295), .Z(DP_mult_204_n2180) );
  INV_X1 DP_mult_204_U1630 ( .A(DP_mult_204_n2145), .ZN(DP_mult_204_n2042) );
  XNOR2_X1 DP_mult_204_U1629 ( .A(DP_mult_204_n2040), .B(DP_mult_204_n1210), 
        .ZN(DP_mult_204_n2041) );
  XNOR2_X1 DP_mult_204_U1628 ( .A(DP_mult_204_n2116), .B(DP_mult_204_n2041), 
        .ZN(DP_mult_204_n835) );
  INV_X2 DP_mult_204_U1627 ( .A(DP_mult_204_n2244), .ZN(DP_mult_204_n2329) );
  OAI22_X1 DP_mult_204_U1626 ( .A1(DP_mult_204_n2304), .A2(DP_mult_204_n1568), 
        .B1(DP_mult_204_n1567), .B2(DP_mult_204_n2329), .ZN(DP_mult_204_n2040)
         );
  XNOR2_X1 DP_mult_204_U1625 ( .A(DP_coeffs_fb_int[13]), .B(DP_mult_204_n2358), 
        .ZN(DP_mult_204_n2145) );
  NAND3_X1 DP_mult_204_U1624 ( .A1(DP_mult_204_n2037), .A2(DP_mult_204_n2038), 
        .A3(DP_mult_204_n2039), .ZN(DP_mult_204_n830) );
  NAND2_X1 DP_mult_204_U1623 ( .A1(DP_mult_204_n1298), .A2(DP_mult_204_n1254), 
        .ZN(DP_mult_204_n2039) );
  NAND2_X1 DP_mult_204_U1622 ( .A1(DP_mult_204_n1320), .A2(DP_mult_204_n1254), 
        .ZN(DP_mult_204_n2038) );
  NAND2_X1 DP_mult_204_U1621 ( .A1(DP_mult_204_n1320), .A2(DP_mult_204_n1298), 
        .ZN(DP_mult_204_n2037) );
  XOR2_X1 DP_mult_204_U1620 ( .A(DP_mult_204_n1320), .B(DP_mult_204_n2036), 
        .Z(DP_mult_204_n831) );
  XOR2_X1 DP_mult_204_U1619 ( .A(DP_mult_204_n1298), .B(DP_mult_204_n1254), 
        .Z(DP_mult_204_n2036) );
  INV_X1 DP_mult_204_U1618 ( .A(DP_mult_204_n2061), .ZN(DP_mult_204_n2248) );
  OAI22_X1 DP_mult_204_U1617 ( .A1(DP_mult_204_n2305), .A2(DP_mult_204_n1577), 
        .B1(DP_mult_204_n2328), .B2(DP_mult_204_n1576), .ZN(DP_mult_204_n2035)
         );
  INV_X1 DP_mult_204_U1616 ( .A(DP_coeffs_fb_int[2]), .ZN(DP_mult_204_n2034)
         );
  INV_X2 DP_mult_204_U1615 ( .A(DP_mult_204_n2001), .ZN(DP_mult_204_n2345) );
  XNOR2_X1 DP_mult_204_U1614 ( .A(DP_coeffs_fb_int[17]), .B(DP_mult_204_n2203), 
        .ZN(DP_mult_204_n1814) );
  BUF_X1 DP_mult_204_U1613 ( .A(DP_mult_204_n1351), .Z(DP_mult_204_n2033) );
  NAND3_X1 DP_mult_204_U1612 ( .A1(DP_mult_204_n2030), .A2(DP_mult_204_n2031), 
        .A3(DP_mult_204_n2032), .ZN(DP_mult_204_n880) );
  NAND2_X1 DP_mult_204_U1611 ( .A1(DP_mult_204_n904), .A2(DP_mult_204_n887), 
        .ZN(DP_mult_204_n2032) );
  NAND2_X1 DP_mult_204_U1610 ( .A1(DP_mult_204_n902), .A2(DP_mult_204_n887), 
        .ZN(DP_mult_204_n2031) );
  NAND2_X1 DP_mult_204_U1609 ( .A1(DP_mult_204_n902), .A2(DP_mult_204_n904), 
        .ZN(DP_mult_204_n2030) );
  XOR2_X1 DP_mult_204_U1608 ( .A(DP_mult_204_n902), .B(DP_mult_204_n2029), .Z(
        DP_mult_204_n881) );
  XOR2_X1 DP_mult_204_U1607 ( .A(DP_mult_204_n904), .B(DP_mult_204_n887), .Z(
        DP_mult_204_n2029) );
  INV_X1 DP_mult_204_U1606 ( .A(DP_mult_204_n2345), .ZN(DP_mult_204_n2028) );
  NAND3_X1 DP_mult_204_U1605 ( .A1(DP_mult_204_n2025), .A2(DP_mult_204_n2026), 
        .A3(DP_mult_204_n2027), .ZN(DP_mult_204_n796) );
  NAND2_X1 DP_mult_204_U1604 ( .A1(DP_mult_204_n1274), .A2(DP_mult_204_n1296), 
        .ZN(DP_mult_204_n2027) );
  NAND2_X1 DP_mult_204_U1603 ( .A1(DP_mult_204_n818), .A2(DP_mult_204_n1296), 
        .ZN(DP_mult_204_n2026) );
  NAND2_X1 DP_mult_204_U1602 ( .A1(DP_mult_204_n818), .A2(DP_mult_204_n1274), 
        .ZN(DP_mult_204_n2025) );
  XOR2_X1 DP_mult_204_U1601 ( .A(DP_mult_204_n818), .B(DP_mult_204_n2024), .Z(
        DP_mult_204_n797) );
  XOR2_X1 DP_mult_204_U1600 ( .A(DP_mult_204_n1274), .B(DP_mult_204_n1296), 
        .Z(DP_mult_204_n2024) );
  XNOR2_X1 DP_mult_204_U1599 ( .A(DP_coeffs_fb_int[9]), .B(DP_mult_204_n2368), 
        .ZN(DP_mult_204_n1810) );
  INV_X2 DP_mult_204_U1598 ( .A(DP_mult_204_n2349), .ZN(DP_mult_204_n2348) );
  NAND3_X1 DP_mult_204_U1597 ( .A1(DP_mult_204_n2020), .A2(DP_mult_204_n2021), 
        .A3(DP_mult_204_n2022), .ZN(DP_mult_204_n862) );
  NAND2_X1 DP_mult_204_U1596 ( .A1(DP_mult_204_n873), .A2(DP_mult_204_n888), 
        .ZN(DP_mult_204_n2022) );
  NAND2_X1 DP_mult_204_U1595 ( .A1(DP_mult_204_n886), .A2(DP_mult_204_n888), 
        .ZN(DP_mult_204_n2021) );
  NAND2_X1 DP_mult_204_U1594 ( .A1(DP_mult_204_n886), .A2(DP_mult_204_n873), 
        .ZN(DP_mult_204_n2020) );
  XOR2_X1 DP_mult_204_U1593 ( .A(DP_coeffs_fb_int[3]), .B(DP_coeffs_fb_int[4]), 
        .Z(DP_mult_204_n2246) );
  INV_X1 DP_mult_204_U1592 ( .A(DP_mult_204_n2324), .ZN(DP_mult_204_n2019) );
  XOR2_X1 DP_mult_204_U1591 ( .A(DP_coeffs_fb_int[19]), .B(
        DP_coeffs_fb_int[20]), .Z(DP_mult_204_n2245) );
  INV_X1 DP_mult_204_U1590 ( .A(DP_mult_204_n2339), .ZN(DP_mult_204_n2018) );
  NOR2_X1 DP_mult_204_U1589 ( .A1(DP_mult_204_n2017), .A2(DP_mult_204_n596), 
        .ZN(DP_mult_204_n594) );
  AND2_X1 DP_mult_204_U1588 ( .A1(DP_mult_204_n595), .A2(DP_mult_204_n609), 
        .ZN(DP_mult_204_n2017) );
  INV_X2 DP_mult_204_U1587 ( .A(DP_mult_204_n2210), .ZN(DP_mult_204_n2359) );
  INV_X2 DP_mult_204_U1586 ( .A(DP_mult_204_n2082), .ZN(DP_mult_204_n2104) );
  AND2_X2 DP_mult_204_U1585 ( .A1(DP_mult_204_n1810), .A2(DP_mult_204_n2330), 
        .ZN(DP_mult_204_n2082) );
  INV_X1 DP_mult_204_U1584 ( .A(DP_mult_204_n2338), .ZN(DP_mult_204_n2015) );
  AND2_X1 DP_mult_204_U1583 ( .A1(DP_mult_204_n1809), .A2(DP_mult_204_n2103), 
        .ZN(DP_mult_204_n2014) );
  AND2_X1 DP_mult_204_U1582 ( .A1(DP_mult_204_n1809), .A2(DP_mult_204_n2103), 
        .ZN(DP_mult_204_n2013) );
  BUF_X1 DP_mult_204_U1581 ( .A(DP_mult_204_n543), .Z(DP_mult_204_n2012) );
  XNOR2_X1 DP_mult_204_U1580 ( .A(DP_coeffs_fb_int[1]), .B(DP_coeffs_fb_int[2]), .ZN(DP_mult_204_n2011) );
  CLKBUF_X1 DP_mult_204_U1579 ( .A(DP_mult_204_n2221), .Z(DP_mult_204_n2010)
         );
  INV_X2 DP_mult_204_U1578 ( .A(DP_mult_204_n2080), .ZN(DP_mult_204_n2178) );
  XNOR2_X1 DP_mult_204_U1577 ( .A(DP_mult_204_n1437), .B(DP_mult_204_n1305), 
        .ZN(DP_mult_204_n2009) );
  XNOR2_X1 DP_mult_204_U1576 ( .A(DP_mult_204_n2009), .B(DP_mult_204_n2101), 
        .ZN(DP_mult_204_n977) );
  XOR2_X1 DP_mult_204_U1575 ( .A(DP_coeffs_fb_int[9]), .B(DP_coeffs_fb_int[10]), .Z(DP_mult_204_n2250) );
  BUF_X1 DP_mult_204_U1574 ( .A(DP_mult_204_n301), .Z(DP_mult_204_n2218) );
  INV_X1 DP_mult_204_U1573 ( .A(DP_mult_204_n2330), .ZN(DP_mult_204_n2008) );
  OR2_X1 DP_mult_204_U1572 ( .A1(DP_mult_204_n789), .A2(DP_mult_204_n804), 
        .ZN(DP_mult_204_n2007) );
  NAND3_X1 DP_mult_204_U1571 ( .A1(DP_mult_204_n2292), .A2(DP_mult_204_n2293), 
        .A3(DP_mult_204_n2294), .ZN(DP_mult_204_n2006) );
  BUF_X1 DP_mult_204_U1570 ( .A(DP_mult_204_n454), .Z(DP_mult_204_n2065) );
  INV_X2 DP_mult_204_U1569 ( .A(DP_coeffs_fb_int[23]), .ZN(DP_mult_204_n251)
         );
  INV_X1 DP_mult_204_U1568 ( .A(DP_coeffs_fb_int[0]), .ZN(DP_mult_204_n2005)
         );
  CLKBUF_X1 DP_mult_204_U1567 ( .A(DP_mult_204_n1933), .Z(DP_mult_204_n2004)
         );
  AND2_X1 DP_mult_204_U1566 ( .A1(DP_mult_204_n2091), .A2(DP_mult_204_n2092), 
        .ZN(DP_mult_204_n2148) );
  AND2_X1 DP_mult_204_U1565 ( .A1(DP_mult_204_n2091), .A2(DP_mult_204_n2092), 
        .ZN(DP_mult_204_n2003) );
  INV_X1 DP_mult_204_U1564 ( .A(DP_mult_204_n554), .ZN(DP_mult_204_n2002) );
  INV_X1 DP_mult_204_U1563 ( .A(DP_coeffs_fb_int[22]), .ZN(DP_mult_204_n2001)
         );
  OR2_X1 DP_mult_204_U1562 ( .A1(DP_mult_204_n1003), .A2(DP_mult_204_n1020), 
        .ZN(DP_mult_204_n2000) );
  AND2_X1 DP_mult_204_U1561 ( .A1(DP_mult_204_n2228), .A2(DP_mult_204_n2229), 
        .ZN(DP_mult_204_n1999) );
  AND2_X1 DP_mult_204_U1560 ( .A1(DP_mult_204_n1999), .A2(DP_mult_204_n2000), 
        .ZN(DP_mult_204_n567) );
  AND2_X1 DP_mult_204_U1559 ( .A1(DP_mult_204_n2146), .A2(DP_mult_204_n559), 
        .ZN(DP_mult_204_n1998) );
  XNOR2_X1 DP_mult_204_U1558 ( .A(DP_mult_204_n560), .B(DP_mult_204_n1998), 
        .ZN(DP_sw0_coeff_ret0[0]) );
  AND2_X1 DP_mult_204_U1557 ( .A1(DP_mult_204_n2265), .A2(DP_mult_204_n550), 
        .ZN(DP_mult_204_n1997) );
  XNOR2_X1 DP_mult_204_U1556 ( .A(DP_mult_204_n551), .B(DP_mult_204_n1997), 
        .ZN(DP_sw0_coeff_ret0[1]) );
  OR2_X1 DP_mult_204_U1555 ( .A1(DP_mult_204_n1194), .A2(DP_mult_204_n676), 
        .ZN(DP_mult_204_n1996) );
  OR2_X1 DP_mult_204_U1554 ( .A1(DP_mult_204_n1151), .A2(DP_mult_204_n1158), 
        .ZN(DP_mult_204_n1995) );
  AND2_X1 DP_mult_204_U1553 ( .A1(DP_mult_204_n1111), .A2(DP_mult_204_n1122), 
        .ZN(DP_mult_204_n1994) );
  AND2_X1 DP_mult_204_U1552 ( .A1(DP_mult_204_n1133), .A2(DP_mult_204_n1142), 
        .ZN(DP_mult_204_n1993) );
  AND2_X1 DP_mult_204_U1551 ( .A1(DP_mult_204_n1179), .A2(DP_mult_204_n1433), 
        .ZN(DP_mult_204_n1992) );
  AND2_X1 DP_mult_204_U1550 ( .A1(DP_mult_204_n1457), .A2(DP_mult_204_n1480), 
        .ZN(DP_mult_204_n1991) );
  AND2_X1 DP_mult_204_U1549 ( .A1(DP_mult_204_n1039), .A2(DP_mult_204_n1054), 
        .ZN(DP_mult_204_n1990) );
  AND2_X1 DP_mult_204_U1548 ( .A1(DP_mult_204_n1238), .A2(DP_mult_204_n1216), 
        .ZN(DP_mult_204_n1989) );
  AND2_X1 DP_mult_204_U1547 ( .A1(DP_mult_204_n1240), .A2(DP_mult_204_n1966), 
        .ZN(DP_mult_204_n1988) );
  AND2_X1 DP_mult_204_U1546 ( .A1(DP_mult_204_n1813), .A2(DP_mult_204_n2176), 
        .ZN(DP_mult_204_n1987) );
  AND2_X1 DP_mult_204_U1545 ( .A1(DP_mult_204_n1151), .A2(DP_mult_204_n1158), 
        .ZN(DP_mult_204_n1986) );
  AND2_X1 DP_mult_204_U1544 ( .A1(DP_mult_204_n1123), .A2(DP_mult_204_n1132), 
        .ZN(DP_mult_204_n1985) );
  AND2_X1 DP_mult_204_U1543 ( .A1(DP_mult_204_n1143), .A2(DP_mult_204_n1150), 
        .ZN(DP_mult_204_n1984) );
  OR2_X1 DP_mult_204_U1542 ( .A1(DP_mult_204_n1179), .A2(DP_mult_204_n1433), 
        .ZN(DP_mult_204_n1983) );
  OR2_X1 DP_mult_204_U1541 ( .A1(DP_mult_204_n1457), .A2(DP_mult_204_n1480), 
        .ZN(DP_mult_204_n1982) );
  AND2_X1 DP_mult_204_U1540 ( .A1(DP_mult_204_n1193), .A2(DP_mult_204_n1481), 
        .ZN(DP_mult_204_n1981) );
  NOR2_X1 DP_mult_204_U1539 ( .A1(DP_mult_204_n789), .A2(DP_mult_204_n804), 
        .ZN(DP_mult_204_n480) );
  BUF_X2 DP_mult_204_U1538 ( .A(DP_mult_204_n293), .Z(DP_mult_204_n2221) );
  AND2_X1 DP_mult_204_U1537 ( .A1(DP_mult_204_n1814), .A2(DP_mult_204_n2336), 
        .ZN(DP_mult_204_n2170) );
  BUF_X2 DP_mult_204_U1536 ( .A(DP_mult_204_n301), .Z(DP_mult_204_n2219) );
  XNOR2_X1 DP_mult_204_U1535 ( .A(DP_mult_204_n873), .B(DP_mult_204_n888), 
        .ZN(DP_mult_204_n1980) );
  XNOR2_X1 DP_mult_204_U1534 ( .A(DP_mult_204_n886), .B(DP_mult_204_n1980), 
        .ZN(DP_mult_204_n863) );
  CLKBUF_X1 DP_mult_204_U1533 ( .A(DP_mult_204_n2246), .Z(DP_mult_204_n1979)
         );
  XNOR2_X1 DP_mult_204_U1532 ( .A(DP_coeffs_fb_int[21]), .B(
        DP_coeffs_fb_int[22]), .ZN(DP_mult_204_n2155) );
  CLKBUF_X1 DP_mult_204_U1531 ( .A(DP_mult_204_n2155), .Z(DP_mult_204_n1978)
         );
  INV_X1 DP_mult_204_U1530 ( .A(DP_mult_204_n2081), .ZN(DP_mult_204_n2307) );
  INV_X1 DP_mult_204_U1529 ( .A(DP_mult_204_n2081), .ZN(DP_mult_204_n1977) );
  INV_X2 DP_mult_204_U1528 ( .A(DP_mult_204_n2352), .ZN(DP_mult_204_n2350) );
  XOR2_X1 DP_mult_204_U1527 ( .A(DP_sw0_23_), .B(DP_mult_204_n2350), .Z(
        DP_mult_204_n1976) );
  INV_X1 DP_mult_204_U1526 ( .A(DP_mult_204_n2350), .ZN(DP_mult_204_n1975) );
  INV_X1 DP_mult_204_U1525 ( .A(DP_mult_204_n2309), .ZN(DP_mult_204_n1973) );
  CLKBUF_X1 DP_mult_204_U1524 ( .A(DP_mult_204_n1027), .Z(DP_mult_204_n1972)
         );
  XNOR2_X1 DP_mult_204_U1523 ( .A(DP_mult_204_n1263), .B(DP_mult_204_n1285), 
        .ZN(DP_mult_204_n1971) );
  XNOR2_X1 DP_mult_204_U1522 ( .A(DP_mult_204_n1971), .B(DP_mult_204_n2033), 
        .ZN(DP_mult_204_n1019) );
  INV_X1 DP_mult_204_U1521 ( .A(DP_mult_204_n2248), .ZN(DP_mult_204_n2333) );
  INV_X2 DP_mult_204_U1520 ( .A(DP_mult_204_n2248), .ZN(DP_mult_204_n1969) );
  INV_X2 DP_mult_204_U1519 ( .A(DP_mult_204_n2248), .ZN(DP_mult_204_n1970) );
  INV_X1 DP_mult_204_U1518 ( .A(DP_mult_204_n1969), .ZN(DP_mult_204_n1968) );
  BUF_X2 DP_mult_204_U1517 ( .A(DP_mult_204_n287), .Z(DP_mult_204_n2257) );
  AND2_X2 DP_mult_204_U1516 ( .A1(DP_mult_204_n1811), .A2(DP_mult_204_n2061), 
        .ZN(DP_mult_204_n2016) );
  INV_X1 DP_mult_204_U1515 ( .A(DP_mult_204_n2016), .ZN(DP_mult_204_n1967) );
  OAI22_X1 DP_mult_204_U1514 ( .A1(DP_mult_204_n2221), .A2(DP_mult_204_n1553), 
        .B1(DP_mult_204_n1552), .B2(DP_mult_204_n2327), .ZN(DP_mult_204_n1966)
         );
  INV_X2 DP_mult_204_U1513 ( .A(DP_mult_204_n2064), .ZN(DP_mult_204_n2322) );
  INV_X2 DP_mult_204_U1512 ( .A(DP_mult_204_n2071), .ZN(DP_mult_204_n2327) );
  NAND3_X1 DP_mult_204_U1511 ( .A1(DP_mult_204_n1963), .A2(DP_mult_204_n1964), 
        .A3(DP_mult_204_n1965), .ZN(DP_mult_204_n860) );
  NAND2_X1 DP_mult_204_U1510 ( .A1(DP_mult_204_n865), .A2(DP_mult_204_n867), 
        .ZN(DP_mult_204_n1965) );
  NAND2_X1 DP_mult_204_U1509 ( .A1(DP_mult_204_n884), .A2(DP_mult_204_n867), 
        .ZN(DP_mult_204_n1964) );
  NAND2_X1 DP_mult_204_U1508 ( .A1(DP_mult_204_n865), .A2(DP_mult_204_n884), 
        .ZN(DP_mult_204_n1963) );
  NAND3_X1 DP_mult_204_U1507 ( .A1(DP_mult_204_n1960), .A2(DP_mult_204_n1961), 
        .A3(DP_mult_204_n1962), .ZN(DP_mult_204_n866) );
  NAND2_X1 DP_mult_204_U1506 ( .A1(DP_mult_204_n1300), .A2(DP_mult_204_n892), 
        .ZN(DP_mult_204_n1962) );
  NAND2_X1 DP_mult_204_U1505 ( .A1(DP_mult_204_n894), .A2(DP_mult_204_n892), 
        .ZN(DP_mult_204_n1961) );
  NAND2_X1 DP_mult_204_U1504 ( .A1(DP_mult_204_n894), .A2(DP_mult_204_n1300), 
        .ZN(DP_mult_204_n1960) );
  XOR2_X1 DP_mult_204_U1503 ( .A(DP_mult_204_n1959), .B(DP_mult_204_n867), .Z(
        DP_mult_204_n861) );
  XOR2_X1 DP_mult_204_U1502 ( .A(DP_mult_204_n865), .B(DP_mult_204_n884), .Z(
        DP_mult_204_n1959) );
  INV_X2 DP_mult_204_U1501 ( .A(DP_mult_204_n1979), .ZN(DP_mult_204_n2325) );
  XNOR2_X1 DP_mult_204_U1500 ( .A(DP_coeffs_fb_int[5]), .B(DP_coeffs_fb_int[6]), .ZN(DP_mult_204_n1958) );
  CLKBUF_X1 DP_mult_204_U1499 ( .A(DP_mult_204_n553), .Z(DP_mult_204_n1957) );
  INV_X1 DP_mult_204_U1498 ( .A(DP_sw0_0_), .ZN(DP_mult_204_n2384) );
  INV_X1 DP_mult_204_U1497 ( .A(DP_sw0_0_), .ZN(DP_mult_204_n1954) );
  INV_X1 DP_mult_204_U1496 ( .A(DP_sw0_0_), .ZN(DP_mult_204_n1955) );
  NAND3_X1 DP_mult_204_U1495 ( .A1(DP_mult_204_n1951), .A2(DP_mult_204_n1952), 
        .A3(DP_mult_204_n1953), .ZN(DP_mult_204_n848) );
  NAND2_X1 DP_mult_204_U1494 ( .A1(DP_mult_204_n1365), .A2(DP_mult_204_n1410), 
        .ZN(DP_mult_204_n1953) );
  NAND2_X1 DP_mult_204_U1493 ( .A1(DP_mult_204_n872), .A2(DP_mult_204_n1410), 
        .ZN(DP_mult_204_n1952) );
  NAND2_X1 DP_mult_204_U1492 ( .A1(DP_mult_204_n872), .A2(DP_mult_204_n1365), 
        .ZN(DP_mult_204_n1951) );
  XOR2_X1 DP_mult_204_U1491 ( .A(DP_mult_204_n872), .B(DP_mult_204_n1950), .Z(
        DP_mult_204_n849) );
  XOR2_X1 DP_mult_204_U1490 ( .A(DP_mult_204_n1365), .B(DP_mult_204_n1410), 
        .Z(DP_mult_204_n1950) );
  XNOR2_X1 DP_mult_204_U1489 ( .A(DP_mult_204_n894), .B(DP_mult_204_n1300), 
        .ZN(DP_mult_204_n1949) );
  XNOR2_X2 DP_mult_204_U1488 ( .A(DP_mult_204_n1949), .B(DP_mult_204_n892), 
        .ZN(DP_mult_204_n867) );
  INV_X1 DP_mult_204_U1487 ( .A(DP_mult_204_n536), .ZN(DP_mult_204_n1948) );
  INV_X2 DP_mult_204_U1486 ( .A(DP_mult_204_n2034), .ZN(DP_mult_204_n2378) );
  INV_X2 DP_mult_204_U1485 ( .A(DP_mult_204_n2203), .ZN(DP_mult_204_n2353) );
  AND2_X1 DP_mult_204_U1484 ( .A1(DP_mult_204_n1814), .A2(DP_mult_204_n2336), 
        .ZN(DP_mult_204_n1946) );
  AND2_X1 DP_mult_204_U1483 ( .A1(DP_mult_204_n1814), .A2(DP_mult_204_n2336), 
        .ZN(DP_mult_204_n1947) );
  INV_X2 DP_mult_204_U1482 ( .A(DP_mult_204_n2034), .ZN(DP_mult_204_n2377) );
  NAND2_X1 DP_mult_204_U1481 ( .A1(DP_mult_204_n672), .A2(DP_mult_204_n535), 
        .ZN(DP_mult_204_n1945) );
  XNOR2_X1 DP_mult_204_U1480 ( .A(DP_mult_204_n1948), .B(DP_mult_204_n1945), 
        .ZN(DP_sw0_coeff_ret0[3]) );
  AND2_X1 DP_mult_204_U1479 ( .A1(DP_mult_204_n663), .A2(DP_mult_204_n439), 
        .ZN(DP_mult_204_n1944) );
  XNOR2_X1 DP_mult_204_U1478 ( .A(DP_mult_204_n2219), .B(DP_mult_204_n1944), 
        .ZN(DP_sw0_coeff_ret0[12]) );
  BUF_X1 DP_mult_204_U1477 ( .A(DP_mult_204_n568), .Z(DP_mult_204_n2117) );
  BUF_X1 DP_mult_204_U1476 ( .A(DP_mult_204_n2250), .Z(DP_mult_204_n1943) );
  BUF_X1 DP_mult_204_U1475 ( .A(DP_mult_204_n1732), .Z(DP_mult_204_n1956) );
  CLKBUF_X1 DP_mult_204_U1474 ( .A(DP_mult_204_n1415), .Z(DP_mult_204_n1974)
         );
  NAND3_X1 DP_mult_204_U1473 ( .A1(DP_mult_204_n1940), .A2(DP_mult_204_n1941), 
        .A3(DP_mult_204_n1942), .ZN(DP_mult_204_n1002) );
  NAND2_X1 DP_mult_204_U1472 ( .A1(DP_mult_204_n1022), .A2(DP_mult_204_n1007), 
        .ZN(DP_mult_204_n1942) );
  NAND2_X1 DP_mult_204_U1471 ( .A1(DP_mult_204_n1005), .A2(DP_mult_204_n1007), 
        .ZN(DP_mult_204_n1941) );
  NAND2_X1 DP_mult_204_U1470 ( .A1(DP_mult_204_n1005), .A2(DP_mult_204_n1022), 
        .ZN(DP_mult_204_n1940) );
  XOR2_X1 DP_mult_204_U1469 ( .A(DP_mult_204_n1005), .B(DP_mult_204_n1939), 
        .Z(DP_mult_204_n1003) );
  XOR2_X1 DP_mult_204_U1468 ( .A(DP_mult_204_n1022), .B(DP_mult_204_n1007), 
        .Z(DP_mult_204_n1939) );
  INV_X1 DP_mult_204_U1467 ( .A(DP_mult_204_n2374), .ZN(DP_mult_204_n1938) );
  BUF_X1 DP_mult_204_U1466 ( .A(DP_mult_204_n2245), .Z(DP_mult_204_n1937) );
  CLKBUF_X2 DP_mult_204_U1465 ( .A(DP_coeffs_fb_int[16]), .Z(DP_mult_204_n2109) );
  OR2_X2 DP_mult_204_U1464 ( .A1(DP_mult_204_n761), .A2(DP_mult_204_n774), 
        .ZN(DP_mult_204_n2226) );
  NAND2_X1 DP_mult_204_U1463 ( .A1(DP_mult_204_n2225), .A2(DP_mult_204_n2226), 
        .ZN(DP_mult_204_n1936) );
  INV_X2 DP_mult_204_U1462 ( .A(DP_mult_204_n2242), .ZN(DP_mult_204_n2121) );
  AND2_X2 DP_mult_204_U1461 ( .A1(DP_mult_204_n1817), .A2(DP_mult_204_n251), 
        .ZN(DP_mult_204_n2242) );
  CLKBUF_X1 DP_mult_204_U1460 ( .A(DP_mult_204_n1934), .Z(DP_mult_204_n2023)
         );
  INV_X2 DP_mult_204_U1459 ( .A(DP_mult_204_n2380), .ZN(DP_mult_204_n2379) );
  INV_X1 DP_mult_204_U1458 ( .A(DP_mult_204_n2372), .ZN(DP_mult_204_n2371) );
  OAI21_X1 DP_mult_204_U1457 ( .B1(DP_mult_204_n594), .B2(DP_mult_204_n582), 
        .A(DP_mult_204_n583), .ZN(DP_mult_204_n1934) );
  NOR2_X1 DP_mult_204_U1456 ( .A1(DP_mult_204_n2163), .A2(DP_mult_204_n520), 
        .ZN(DP_mult_204_n1933) );
  NOR2_X1 DP_mult_204_U1455 ( .A1(DP_mult_204_n542), .A2(DP_mult_204_n547), 
        .ZN(DP_mult_204_n1932) );
  INV_X2 DP_mult_204_U1454 ( .A(DP_mult_204_n2365), .ZN(DP_mult_204_n2364) );
  INV_X1 DP_mult_204_U1453 ( .A(DP_mult_204_n2364), .ZN(DP_mult_204_n1931) );
  AND2_X2 DP_mult_204_U1452 ( .A1(DP_mult_204_n1815), .A2(DP_mult_204_n2339), 
        .ZN(DP_mult_204_n2080) );
  XNOR2_X1 DP_mult_204_U1451 ( .A(DP_coeffs_fb_int[19]), .B(DP_mult_204_n2352), 
        .ZN(DP_mult_204_n1815) );
  OAI22_X1 DP_mult_204_U1450 ( .A1(DP_mult_204_n2313), .A2(DP_mult_204_n1683), 
        .B1(DP_mult_204_n1682), .B2(DP_mult_204_n2338), .ZN(DP_mult_204_n1930)
         );
  BUF_X1 DP_mult_204_U1449 ( .A(DP_coeffs_fb_int[20]), .Z(DP_mult_204_n1935)
         );
  BUF_X2 DP_mult_204_U1448 ( .A(DP_mult_204_n2343), .Z(DP_mult_204_n1929) );
  HA_X1 DP_mult_204_U798 ( .A(DP_mult_204_n1456), .B(DP_mult_204_n1479), .CO(
        DP_mult_204_n1180), .S(DP_mult_204_n1181) );
  FA_X1 DP_mult_204_U797 ( .A(DP_mult_204_n1455), .B(DP_mult_204_n1478), .CI(
        DP_mult_204_n1180), .CO(DP_mult_204_n1178), .S(DP_mult_204_n1179) );
  HA_X1 DP_mult_204_U796 ( .A(DP_mult_204_n1432), .B(DP_mult_204_n1477), .CO(
        DP_mult_204_n1176), .S(DP_mult_204_n1177) );
  FA_X1 DP_mult_204_U795 ( .A(DP_mult_204_n1191), .B(DP_mult_204_n1454), .CI(
        DP_mult_204_n1177), .CO(DP_mult_204_n1174), .S(DP_mult_204_n1175) );
  FA_X1 DP_mult_204_U794 ( .A(DP_mult_204_n1476), .B(DP_mult_204_n1431), .CI(
        DP_mult_204_n1453), .CO(DP_mult_204_n1172), .S(DP_mult_204_n1173) );
  FA_X1 DP_mult_204_U793 ( .A(DP_mult_204_n1409), .B(DP_mult_204_n1176), .CI(
        DP_mult_204_n1173), .CO(DP_mult_204_n1170), .S(DP_mult_204_n1171) );
  HA_X1 DP_mult_204_U792 ( .A(DP_mult_204_n1408), .B(DP_mult_204_n1430), .CO(
        DP_mult_204_n1168), .S(DP_mult_204_n1169) );
  FA_X1 DP_mult_204_U791 ( .A(DP_mult_204_n1452), .B(DP_mult_204_n1475), .CI(
        DP_mult_204_n1190), .CO(DP_mult_204_n1166), .S(DP_mult_204_n1167) );
  FA_X1 DP_mult_204_U790 ( .A(DP_mult_204_n1172), .B(DP_mult_204_n1169), .CI(
        DP_mult_204_n1167), .CO(DP_mult_204_n1164), .S(DP_mult_204_n1165) );
  FA_X1 DP_mult_204_U789 ( .A(DP_mult_204_n1451), .B(DP_mult_204_n1474), .CI(
        DP_mult_204_n1407), .CO(DP_mult_204_n1162), .S(DP_mult_204_n1163) );
  FA_X1 DP_mult_204_U788 ( .A(DP_mult_204_n1168), .B(DP_mult_204_n1429), .CI(
        DP_mult_204_n1166), .CO(DP_mult_204_n1160), .S(DP_mult_204_n1161) );
  FA_X1 DP_mult_204_U787 ( .A(DP_mult_204_n1163), .B(DP_mult_204_n1385), .CI(
        DP_mult_204_n1164), .CO(DP_mult_204_n1158), .S(DP_mult_204_n1159) );
  HA_X1 DP_mult_204_U786 ( .A(DP_mult_204_n1384), .B(DP_mult_204_n1406), .CO(
        DP_mult_204_n1156), .S(DP_mult_204_n1157) );
  FA_X1 DP_mult_204_U785 ( .A(DP_mult_204_n1450), .B(DP_mult_204_n1428), .CI(
        DP_mult_204_n1189), .CO(DP_mult_204_n1154), .S(DP_mult_204_n1155) );
  FA_X1 DP_mult_204_U784 ( .A(DP_mult_204_n1157), .B(DP_mult_204_n1473), .CI(
        DP_mult_204_n1162), .CO(DP_mult_204_n1152), .S(DP_mult_204_n1153) );
  FA_X1 DP_mult_204_U783 ( .A(DP_mult_204_n1160), .B(DP_mult_204_n1155), .CI(
        DP_mult_204_n1153), .CO(DP_mult_204_n1150), .S(DP_mult_204_n1151) );
  FA_X1 DP_mult_204_U782 ( .A(DP_mult_204_n1383), .B(DP_mult_204_n1472), .CI(
        DP_mult_204_n1405), .CO(DP_mult_204_n1148), .S(DP_mult_204_n1149) );
  FA_X1 DP_mult_204_U781 ( .A(DP_mult_204_n1427), .B(DP_mult_204_n1449), .CI(
        DP_mult_204_n1156), .CO(DP_mult_204_n1146), .S(DP_mult_204_n1147) );
  FA_X1 DP_mult_204_U780 ( .A(DP_mult_204_n1361), .B(DP_mult_204_n1154), .CI(
        DP_mult_204_n1149), .CO(DP_mult_204_n1144), .S(DP_mult_204_n1145) );
  FA_X1 DP_mult_204_U779 ( .A(DP_mult_204_n1152), .B(DP_mult_204_n1147), .CI(
        DP_mult_204_n1145), .CO(DP_mult_204_n1142), .S(DP_mult_204_n1143) );
  HA_X1 DP_mult_204_U778 ( .A(DP_mult_204_n1360), .B(DP_mult_204_n1382), .CO(
        DP_mult_204_n1140), .S(DP_mult_204_n1141) );
  FA_X1 DP_mult_204_U777 ( .A(DP_mult_204_n1471), .B(DP_mult_204_n1188), .CI(
        DP_mult_204_n1426), .CO(DP_mult_204_n1138), .S(DP_mult_204_n1139) );
  FA_X1 DP_mult_204_U776 ( .A(DP_mult_204_n1404), .B(DP_mult_204_n1448), .CI(
        DP_mult_204_n1141), .CO(DP_mult_204_n1136), .S(DP_mult_204_n1137) );
  FA_X1 DP_mult_204_U775 ( .A(DP_mult_204_n1146), .B(DP_mult_204_n1148), .CI(
        DP_mult_204_n1139), .CO(DP_mult_204_n1134), .S(DP_mult_204_n1135) );
  FA_X1 DP_mult_204_U774 ( .A(DP_mult_204_n1144), .B(DP_mult_204_n1137), .CI(
        DP_mult_204_n1135), .CO(DP_mult_204_n1132), .S(DP_mult_204_n1133) );
  FA_X1 DP_mult_204_U773 ( .A(DP_mult_204_n1359), .B(DP_mult_204_n1470), .CI(
        DP_mult_204_n1381), .CO(DP_mult_204_n1130), .S(DP_mult_204_n1131) );
  FA_X1 DP_mult_204_U772 ( .A(DP_mult_204_n1403), .B(DP_mult_204_n1447), .CI(
        DP_mult_204_n1425), .CO(DP_mult_204_n1128), .S(DP_mult_204_n1129) );
  FA_X1 DP_mult_204_U771 ( .A(DP_mult_204_n1337), .B(DP_mult_204_n1140), .CI(
        DP_mult_204_n1138), .CO(DP_mult_204_n1126), .S(DP_mult_204_n1127) );
  FA_X1 DP_mult_204_U770 ( .A(DP_mult_204_n1131), .B(DP_mult_204_n1129), .CI(
        DP_mult_204_n1136), .CO(DP_mult_204_n1124), .S(DP_mult_204_n1125) );
  FA_X1 DP_mult_204_U769 ( .A(DP_mult_204_n1127), .B(DP_mult_204_n1134), .CI(
        DP_mult_204_n1125), .CO(DP_mult_204_n1122), .S(DP_mult_204_n1123) );
  HA_X1 DP_mult_204_U768 ( .A(DP_mult_204_n1336), .B(DP_mult_204_n1358), .CO(
        DP_mult_204_n1120), .S(DP_mult_204_n1121) );
  FA_X1 DP_mult_204_U767 ( .A(DP_mult_204_n1380), .B(DP_mult_204_n1187), .CI(
        DP_mult_204_n1402), .CO(DP_mult_204_n1118), .S(DP_mult_204_n1119) );
  FA_X1 DP_mult_204_U766 ( .A(DP_mult_204_n1424), .B(DP_mult_204_n1469), .CI(
        DP_mult_204_n1446), .CO(DP_mult_204_n1116), .S(DP_mult_204_n1117) );
  FA_X1 DP_mult_204_U765 ( .A(DP_mult_204_n1130), .B(DP_mult_204_n1121), .CI(
        DP_mult_204_n1128), .CO(DP_mult_204_n1114), .S(DP_mult_204_n1115) );
  FA_X1 DP_mult_204_U764 ( .A(DP_mult_204_n1119), .B(DP_mult_204_n1117), .CI(
        DP_mult_204_n1126), .CO(DP_mult_204_n1112), .S(DP_mult_204_n1113) );
  FA_X1 DP_mult_204_U763 ( .A(DP_mult_204_n1124), .B(DP_mult_204_n1115), .CI(
        DP_mult_204_n1113), .CO(DP_mult_204_n1110), .S(DP_mult_204_n1111) );
  FA_X1 DP_mult_204_U762 ( .A(DP_mult_204_n1335), .B(DP_mult_204_n1468), .CI(
        DP_mult_204_n1357), .CO(DP_mult_204_n1108), .S(DP_mult_204_n1109) );
  FA_X1 DP_mult_204_U761 ( .A(DP_mult_204_n1379), .B(DP_mult_204_n1445), .CI(
        DP_mult_204_n1401), .CO(DP_mult_204_n1106), .S(DP_mult_204_n1107) );
  FA_X1 DP_mult_204_U760 ( .A(DP_mult_204_n1120), .B(DP_mult_204_n1423), .CI(
        DP_mult_204_n1118), .CO(DP_mult_204_n1104), .S(DP_mult_204_n1105) );
  FA_X1 DP_mult_204_U759 ( .A(DP_mult_204_n1313), .B(DP_mult_204_n1116), .CI(
        DP_mult_204_n1107), .CO(DP_mult_204_n1102), .S(DP_mult_204_n1103) );
  FA_X1 DP_mult_204_U758 ( .A(DP_mult_204_n1114), .B(DP_mult_204_n1109), .CI(
        DP_mult_204_n1105), .CO(DP_mult_204_n1100), .S(DP_mult_204_n1101) );
  FA_X1 DP_mult_204_U757 ( .A(DP_mult_204_n1103), .B(DP_mult_204_n1112), .CI(
        DP_mult_204_n1101), .CO(DP_mult_204_n1098), .S(DP_mult_204_n1099) );
  HA_X1 DP_mult_204_U756 ( .A(DP_mult_204_n1334), .B(DP_mult_204_n1312), .CO(
        DP_mult_204_n1096), .S(DP_mult_204_n1097) );
  FA_X1 DP_mult_204_U755 ( .A(DP_mult_204_n1186), .B(DP_mult_204_n1467), .CI(
        DP_mult_204_n1400), .CO(DP_mult_204_n1094), .S(DP_mult_204_n1095) );
  FA_X1 DP_mult_204_U754 ( .A(DP_mult_204_n1356), .B(DP_mult_204_n1444), .CI(
        DP_mult_204_n1378), .CO(DP_mult_204_n1092), .S(DP_mult_204_n1093) );
  FA_X1 DP_mult_204_U753 ( .A(DP_mult_204_n1097), .B(DP_mult_204_n1422), .CI(
        DP_mult_204_n1108), .CO(DP_mult_204_n1090), .S(DP_mult_204_n1091) );
  FA_X1 DP_mult_204_U752 ( .A(DP_mult_204_n1093), .B(DP_mult_204_n1106), .CI(
        DP_mult_204_n1095), .CO(DP_mult_204_n1088), .S(DP_mult_204_n1089) );
  FA_X1 DP_mult_204_U751 ( .A(DP_mult_204_n1102), .B(DP_mult_204_n1104), .CI(
        DP_mult_204_n1091), .CO(DP_mult_204_n1086), .S(DP_mult_204_n1087) );
  FA_X1 DP_mult_204_U750 ( .A(DP_mult_204_n1100), .B(DP_mult_204_n1089), .CI(
        DP_mult_204_n1087), .CO(DP_mult_204_n1084), .S(DP_mult_204_n1085) );
  FA_X1 DP_mult_204_U749 ( .A(DP_mult_204_n1311), .B(DP_mult_204_n1466), .CI(
        DP_mult_204_n1333), .CO(DP_mult_204_n1082), .S(DP_mult_204_n1083) );
  FA_X1 DP_mult_204_U748 ( .A(DP_mult_204_n1355), .B(DP_mult_204_n1443), .CI(
        DP_mult_204_n1377), .CO(DP_mult_204_n1080), .S(DP_mult_204_n1081) );
  FA_X1 DP_mult_204_U747 ( .A(DP_mult_204_n1399), .B(DP_mult_204_n1421), .CI(
        DP_mult_204_n1096), .CO(DP_mult_204_n1078), .S(DP_mult_204_n1079) );
  FA_X1 DP_mult_204_U746 ( .A(DP_mult_204_n1092), .B(DP_mult_204_n1094), .CI(
        DP_mult_204_n1289), .CO(DP_mult_204_n1076), .S(DP_mult_204_n1077) );
  FA_X1 DP_mult_204_U745 ( .A(DP_mult_204_n1083), .B(DP_mult_204_n1081), .CI(
        DP_mult_204_n1079), .CO(DP_mult_204_n1074), .S(DP_mult_204_n1075) );
  FA_X1 DP_mult_204_U744 ( .A(DP_mult_204_n1088), .B(DP_mult_204_n1090), .CI(
        DP_mult_204_n1077), .CO(DP_mult_204_n1072), .S(DP_mult_204_n1073) );
  FA_X1 DP_mult_204_U743 ( .A(DP_mult_204_n1086), .B(DP_mult_204_n1075), .CI(
        DP_mult_204_n1073), .CO(DP_mult_204_n1070), .S(DP_mult_204_n1071) );
  HA_X1 DP_mult_204_U742 ( .A(DP_mult_204_n1288), .B(DP_mult_204_n1310), .CO(
        DP_mult_204_n1068), .S(DP_mult_204_n1069) );
  FA_X1 DP_mult_204_U741 ( .A(DP_mult_204_n1465), .B(DP_mult_204_n1376), .CI(
        DP_mult_204_n1185), .CO(DP_mult_204_n1066), .S(DP_mult_204_n1067) );
  FA_X1 DP_mult_204_U740 ( .A(DP_mult_204_n1442), .B(DP_mult_204_n1354), .CI(
        DP_mult_204_n1332), .CO(DP_mult_204_n1064), .S(DP_mult_204_n1065) );
  FA_X1 DP_mult_204_U739 ( .A(DP_mult_204_n1398), .B(DP_mult_204_n1420), .CI(
        DP_mult_204_n1069), .CO(DP_mult_204_n1062), .S(DP_mult_204_n1063) );
  FA_X1 DP_mult_204_U738 ( .A(DP_mult_204_n1080), .B(DP_mult_204_n1082), .CI(
        DP_mult_204_n1078), .CO(DP_mult_204_n1060), .S(DP_mult_204_n1061) );
  FA_X1 DP_mult_204_U737 ( .A(DP_mult_204_n1067), .B(DP_mult_204_n1065), .CI(
        DP_mult_204_n1076), .CO(DP_mult_204_n1058), .S(DP_mult_204_n1059) );
  FA_X1 DP_mult_204_U736 ( .A(DP_mult_204_n1074), .B(DP_mult_204_n1063), .CI(
        DP_mult_204_n1061), .CO(DP_mult_204_n1056), .S(DP_mult_204_n1057) );
  FA_X1 DP_mult_204_U735 ( .A(DP_mult_204_n1072), .B(DP_mult_204_n1059), .CI(
        DP_mult_204_n1057), .CO(DP_mult_204_n1054), .S(DP_mult_204_n1055) );
  FA_X1 DP_mult_204_U734 ( .A(DP_mult_204_n1309), .B(DP_mult_204_n1287), .CI(
        DP_mult_204_n1464), .CO(DP_mult_204_n1052), .S(DP_mult_204_n1053) );
  FA_X1 DP_mult_204_U733 ( .A(DP_mult_204_n1331), .B(DP_mult_204_n1353), .CI(
        DP_mult_204_n1375), .CO(DP_mult_204_n1050), .S(DP_mult_204_n1051) );
  FA_X1 DP_mult_204_U732 ( .A(DP_mult_204_n1397), .B(DP_mult_204_n1441), .CI(
        DP_mult_204_n1419), .CO(DP_mult_204_n1048), .S(DP_mult_204_n1049) );
  FA_X1 DP_mult_204_U731 ( .A(DP_mult_204_n1064), .B(DP_mult_204_n1068), .CI(
        DP_mult_204_n1066), .CO(DP_mult_204_n1046), .S(DP_mult_204_n1047) );
  FA_X1 DP_mult_204_U730 ( .A(DP_mult_204_n1049), .B(DP_mult_204_n1265), .CI(
        DP_mult_204_n1051), .CO(DP_mult_204_n1044), .S(DP_mult_204_n1045) );
  FA_X1 DP_mult_204_U729 ( .A(DP_mult_204_n1062), .B(DP_mult_204_n1053), .CI(
        DP_mult_204_n1060), .CO(DP_mult_204_n1042), .S(DP_mult_204_n1043) );
  FA_X1 DP_mult_204_U728 ( .A(DP_mult_204_n1045), .B(DP_mult_204_n1047), .CI(
        DP_mult_204_n1058), .CO(DP_mult_204_n1040), .S(DP_mult_204_n1041) );
  HA_X1 DP_mult_204_U726 ( .A(DP_mult_204_n1264), .B(DP_mult_204_n1286), .CO(
        DP_mult_204_n1036), .S(DP_mult_204_n1037) );
  FA_X1 DP_mult_204_U725 ( .A(DP_mult_204_n1308), .B(DP_mult_204_n1374), .CI(
        DP_mult_204_n1184), .CO(DP_mult_204_n1034), .S(DP_mult_204_n1035) );
  FA_X1 DP_mult_204_U724 ( .A(DP_mult_204_n1463), .B(DP_mult_204_n1396), .CI(
        DP_mult_204_n1330), .CO(DP_mult_204_n1032), .S(DP_mult_204_n1033) );
  FA_X1 DP_mult_204_U723 ( .A(DP_mult_204_n1352), .B(DP_mult_204_n1440), .CI(
        DP_mult_204_n1418), .CO(DP_mult_204_n1030), .S(DP_mult_204_n1031) );
  FA_X1 DP_mult_204_U722 ( .A(DP_mult_204_n1052), .B(DP_mult_204_n1037), .CI(
        DP_mult_204_n1050), .CO(DP_mult_204_n1028), .S(DP_mult_204_n1029) );
  FA_X1 DP_mult_204_U721 ( .A(DP_mult_204_n1033), .B(DP_mult_204_n1048), .CI(
        DP_mult_204_n1031), .CO(DP_mult_204_n1026), .S(DP_mult_204_n1027) );
  FA_X1 DP_mult_204_U720 ( .A(DP_mult_204_n1046), .B(DP_mult_204_n1035), .CI(
        DP_mult_204_n1029), .CO(DP_mult_204_n1024), .S(DP_mult_204_n1025) );
  FA_X1 DP_mult_204_U718 ( .A(DP_mult_204_n1040), .B(DP_mult_204_n1025), .CI(
        DP_mult_204_n1023), .CO(DP_mult_204_n1020), .S(DP_mult_204_n1021) );
  FA_X1 DP_mult_204_U716 ( .A(DP_mult_204_n1307), .B(DP_mult_204_n1373), .CI(
        DP_mult_204_n1329), .CO(DP_mult_204_n1016), .S(DP_mult_204_n1017) );
  FA_X1 DP_mult_204_U715 ( .A(DP_mult_204_n1417), .B(DP_mult_204_n1462), .CI(
        DP_mult_204_n1395), .CO(DP_mult_204_n1014), .S(DP_mult_204_n1015) );
  FA_X1 DP_mult_204_U713 ( .A(DP_mult_204_n1030), .B(DP_mult_204_n1034), .CI(
        DP_mult_204_n1241), .CO(DP_mult_204_n1010), .S(DP_mult_204_n1011) );
  FA_X1 DP_mult_204_U712 ( .A(DP_mult_204_n1015), .B(DP_mult_204_n1019), .CI(
        DP_mult_204_n1017), .CO(DP_mult_204_n1008), .S(DP_mult_204_n1009) );
  FA_X1 DP_mult_204_U711 ( .A(DP_mult_204_n1013), .B(DP_mult_204_n1028), .CI(
        DP_mult_204_n1026), .CO(DP_mult_204_n1006), .S(DP_mult_204_n1007) );
  FA_X1 DP_mult_204_U710 ( .A(DP_mult_204_n1009), .B(DP_mult_204_n1011), .CI(
        DP_mult_204_n1024), .CO(DP_mult_204_n1004), .S(DP_mult_204_n1005) );
  FA_X1 DP_mult_204_U707 ( .A(DP_mult_204_n1183), .B(DP_mult_204_n1350), .CI(
        DP_mult_204_n1461), .CO(DP_mult_204_n998), .S(DP_mult_204_n999) );
  FA_X1 DP_mult_204_U706 ( .A(DP_mult_204_n1284), .B(DP_mult_204_n1372), .CI(
        DP_mult_204_n1438), .CO(DP_mult_204_n996), .S(DP_mult_204_n997) );
  FA_X1 DP_mult_204_U705 ( .A(DP_mult_204_n1328), .B(DP_mult_204_n1416), .CI(
        DP_mult_204_n1306), .CO(DP_mult_204_n994), .S(DP_mult_204_n995) );
  FA_X1 DP_mult_204_U704 ( .A(DP_mult_204_n1001), .B(DP_mult_204_n1394), .CI(
        DP_mult_204_n1018), .CO(DP_mult_204_n992), .S(DP_mult_204_n993) );
  FA_X1 DP_mult_204_U703 ( .A(DP_mult_204_n1014), .B(DP_mult_204_n1016), .CI(
        DP_mult_204_n995), .CO(DP_mult_204_n990), .S(DP_mult_204_n991) );
  FA_X1 DP_mult_204_U701 ( .A(DP_mult_204_n993), .B(DP_mult_204_n1010), .CI(
        DP_mult_204_n1008), .CO(DP_mult_204_n986), .S(DP_mult_204_n987) );
  FA_X1 DP_mult_204_U700 ( .A(DP_mult_204_n989), .B(DP_mult_204_n991), .CI(
        DP_mult_204_n1006), .CO(DP_mult_204_n984), .S(DP_mult_204_n985) );
  FA_X1 DP_mult_204_U699 ( .A(DP_mult_204_n1004), .B(DP_mult_204_n987), .CI(
        DP_mult_204_n985), .CO(DP_mult_204_n982), .S(DP_mult_204_n983) );
  FA_X1 DP_mult_204_U698 ( .A(DP_mult_204_n1239), .B(DP_mult_204_n1349), .CI(
        DP_mult_204_n1261), .CO(DP_mult_204_n980), .S(DP_mult_204_n981) );
  FA_X1 DP_mult_204_U697 ( .A(DP_mult_204_n1371), .B(DP_mult_204_n1460), .CI(
        DP_mult_204_n1283), .CO(DP_mult_204_n978), .S(DP_mult_204_n979) );
  FA_X1 DP_mult_204_U692 ( .A(DP_mult_204_n975), .B(DP_mult_204_n981), .CI(
        DP_mult_204_n992), .CO(DP_mult_204_n968), .S(DP_mult_204_n969) );
  FA_X1 DP_mult_204_U691 ( .A(DP_mult_204_n973), .B(DP_mult_204_n990), .CI(
        DP_mult_204_n988), .CO(DP_mult_204_n966), .S(DP_mult_204_n967) );
  FA_X1 DP_mult_204_U690 ( .A(DP_mult_204_n969), .B(DP_mult_204_n971), .CI(
        DP_mult_204_n986), .CO(DP_mult_204_n964), .S(DP_mult_204_n965) );
  FA_X1 DP_mult_204_U689 ( .A(DP_mult_204_n984), .B(DP_mult_204_n967), .CI(
        DP_mult_204_n965), .CO(DP_mult_204_n962), .S(DP_mult_204_n963) );
  FA_X1 DP_mult_204_U684 ( .A(DP_mult_204_n1326), .B(DP_mult_204_n1392), .CI(
        DP_mult_204_n961), .CO(DP_mult_204_n952), .S(DP_mult_204_n953) );
  FA_X1 DP_mult_204_U683 ( .A(DP_mult_204_n976), .B(DP_mult_204_n980), .CI(
        DP_mult_204_n978), .CO(DP_mult_204_n950), .S(DP_mult_204_n951) );
  FA_X1 DP_mult_204_U682 ( .A(DP_mult_204_n955), .B(DP_mult_204_n974), .CI(
        DP_mult_204_n957), .CO(DP_mult_204_n948), .S(DP_mult_204_n949) );
  FA_X1 DP_mult_204_U680 ( .A(DP_mult_204_n951), .B(DP_mult_204_n970), .CI(
        DP_mult_204_n968), .CO(DP_mult_204_n944), .S(DP_mult_204_n945) );
  FA_X1 DP_mult_204_U679 ( .A(DP_mult_204_n947), .B(DP_mult_204_n949), .CI(
        DP_mult_204_n966), .CO(DP_mult_204_n942), .S(DP_mult_204_n943) );
  FA_X1 DP_mult_204_U675 ( .A(DP_mult_204_n1259), .B(DP_mult_204_n1347), .CI(
        DP_mult_204_n1303), .CO(DP_mult_204_n936), .S(DP_mult_204_n937) );
  FA_X1 DP_mult_204_U674 ( .A(DP_mult_204_n1281), .B(DP_mult_204_n1391), .CI(
        DP_mult_204_n1369), .CO(DP_mult_204_n934), .S(DP_mult_204_n935) );
  FA_X1 DP_mult_204_U672 ( .A(DP_mult_204_n1458), .B(DP_mult_204_n1989), .CI(
        DP_mult_204_n939), .CO(DP_mult_204_n930), .S(DP_mult_204_n931) );
  FA_X1 DP_mult_204_U671 ( .A(DP_mult_204_n954), .B(DP_mult_204_n958), .CI(
        DP_mult_204_n956), .CO(DP_mult_204_n928), .S(DP_mult_204_n929) );
  FA_X1 DP_mult_204_U669 ( .A(DP_mult_204_n931), .B(DP_mult_204_n935), .CI(
        DP_mult_204_n950), .CO(DP_mult_204_n924), .S(DP_mult_204_n925) );
  FA_X1 DP_mult_204_U667 ( .A(DP_mult_204_n925), .B(DP_mult_204_n927), .CI(
        DP_mult_204_n944), .CO(DP_mult_204_n920), .S(DP_mult_204_n921) );
  FA_X1 DP_mult_204_U666 ( .A(DP_mult_204_n942), .B(DP_mult_204_n923), .CI(
        DP_mult_204_n921), .CO(DP_mult_204_n918), .S(DP_mult_204_n919) );
  FA_X1 DP_mult_204_U664 ( .A(DP_mult_204_n1302), .B(DP_mult_204_n1214), .CI(
        DP_mult_204_n917), .CO(DP_mult_204_n914), .S(DP_mult_204_n915) );
  FA_X1 DP_mult_204_U663 ( .A(DP_mult_204_n1236), .B(DP_mult_204_n1258), .CI(
        DP_mult_204_n1412), .CO(DP_mult_204_n912), .S(DP_mult_204_n913) );
  FA_X1 DP_mult_204_U662 ( .A(DP_mult_204_n1280), .B(DP_mult_204_n1346), .CI(
        DP_mult_204_n1324), .CO(DP_mult_204_n910), .S(DP_mult_204_n911) );
  FA_X1 DP_mult_204_U661 ( .A(DP_mult_204_n1368), .B(DP_mult_204_n1390), .CI(
        DP_mult_204_n938), .CO(DP_mult_204_n908), .S(DP_mult_204_n909) );
  FA_X1 DP_mult_204_U660 ( .A(DP_mult_204_n932), .B(DP_mult_204_n936), .CI(
        DP_mult_204_n934), .CO(DP_mult_204_n906), .S(DP_mult_204_n907) );
  FA_X1 DP_mult_204_U659 ( .A(DP_mult_204_n915), .B(DP_mult_204_n911), .CI(
        DP_mult_204_n913), .CO(DP_mult_204_n904), .S(DP_mult_204_n905) );
  FA_X1 DP_mult_204_U658 ( .A(DP_mult_204_n909), .B(DP_mult_204_n930), .CI(
        DP_mult_204_n928), .CO(DP_mult_204_n902), .S(DP_mult_204_n903) );
  FA_X1 DP_mult_204_U657 ( .A(DP_mult_204_n907), .B(DP_mult_204_n926), .CI(
        DP_mult_204_n905), .CO(DP_mult_204_n900), .S(DP_mult_204_n901) );
  FA_X1 DP_mult_204_U654 ( .A(DP_mult_204_n1411), .B(DP_mult_204_n1213), .CI(
        DP_mult_204_n1235), .CO(DP_mult_204_n894), .S(DP_mult_204_n895) );
  FA_X1 DP_mult_204_U653 ( .A(DP_mult_204_n1323), .B(DP_mult_204_n916), .CI(
        DP_mult_204_n1279), .CO(DP_mult_204_n892), .S(DP_mult_204_n893) );
  FA_X1 DP_mult_204_U652 ( .A(DP_mult_204_n1257), .B(DP_mult_204_n1301), .CI(
        DP_mult_204_n1345), .CO(DP_mult_204_n890), .S(DP_mult_204_n891) );
  FA_X1 DP_mult_204_U651 ( .A(DP_mult_204_n1367), .B(DP_mult_204_n1389), .CI(
        DP_mult_204_n1434), .CO(DP_mult_204_n888), .S(DP_mult_204_n889) );
  FA_X1 DP_mult_204_U650 ( .A(DP_mult_204_n910), .B(DP_mult_204_n914), .CI(
        DP_mult_204_n912), .CO(DP_mult_204_n886), .S(DP_mult_204_n887) );
  FA_X1 DP_mult_204_U646 ( .A(DP_mult_204_n883), .B(DP_mult_204_n885), .CI(
        DP_mult_204_n900), .CO(DP_mult_204_n878), .S(DP_mult_204_n879) );
  FA_X1 DP_mult_204_U645 ( .A(DP_mult_204_n898), .B(DP_mult_204_n881), .CI(
        DP_mult_204_n879), .CO(DP_mult_204_n876), .S(DP_mult_204_n877) );
  FA_X1 DP_mult_204_U643 ( .A(DP_mult_204_n1388), .B(DP_mult_204_n1278), .CI(
        DP_mult_204_n875), .CO(DP_mult_204_n872), .S(DP_mult_204_n873) );
  FA_X1 DP_mult_204_U642 ( .A(DP_mult_204_n1344), .B(DP_mult_204_n1366), .CI(
        DP_mult_204_n1212), .CO(DP_mult_204_n870), .S(DP_mult_204_n871) );
  FA_X1 DP_mult_204_U641 ( .A(DP_mult_204_n1256), .B(DP_mult_204_n1322), .CI(
        DP_mult_204_n1234), .CO(DP_mult_204_n868), .S(DP_mult_204_n869) );
  FA_X1 DP_mult_204_U639 ( .A(DP_mult_204_n869), .B(DP_mult_204_n890), .CI(
        DP_mult_204_n871), .CO(DP_mult_204_n864), .S(DP_mult_204_n865) );
  FA_X1 DP_mult_204_U635 ( .A(DP_mult_204_n878), .B(DP_mult_204_n861), .CI(
        DP_mult_204_n859), .CO(DP_mult_204_n856), .S(DP_mult_204_n857) );
  FA_X1 DP_mult_204_U634 ( .A(DP_mult_204_n1211), .B(DP_mult_204_n1233), .CI(
        DP_mult_204_n1387), .CO(DP_mult_204_n854), .S(DP_mult_204_n855) );
  FA_X1 DP_mult_204_U633 ( .A(DP_mult_204_n1255), .B(DP_mult_204_n1321), .CI(
        DP_mult_204_n874), .CO(DP_mult_204_n852), .S(DP_mult_204_n853) );
  FA_X1 DP_mult_204_U632 ( .A(DP_mult_204_n1343), .B(DP_mult_204_n1299), .CI(
        DP_mult_204_n1277), .CO(DP_mult_204_n850), .S(DP_mult_204_n851) );
  FA_X1 DP_mult_204_U630 ( .A(DP_mult_204_n868), .B(DP_mult_204_n870), .CI(
        DP_mult_204_n851), .CO(DP_mult_204_n846), .S(DP_mult_204_n847) );
  FA_X1 DP_mult_204_U627 ( .A(DP_mult_204_n845), .B(DP_mult_204_n847), .CI(
        DP_mult_204_n860), .CO(DP_mult_204_n840), .S(DP_mult_204_n841) );
  FA_X1 DP_mult_204_U626 ( .A(DP_mult_204_n858), .B(DP_mult_204_n843), .CI(
        DP_mult_204_n841), .CO(DP_mult_204_n838), .S(DP_mult_204_n839) );
  FA_X1 DP_mult_204_U623 ( .A(DP_mult_204_n1232), .B(DP_mult_204_n1364), .CI(
        DP_mult_204_n1342), .CO(DP_mult_204_n832), .S(DP_mult_204_n833) );
  FA_X1 DP_mult_204_U621 ( .A(DP_mult_204_n850), .B(DP_mult_204_n854), .CI(
        DP_mult_204_n852), .CO(DP_mult_204_n828), .S(DP_mult_204_n829) );
  FA_X1 DP_mult_204_U620 ( .A(DP_mult_204_n835), .B(DP_mult_204_n831), .CI(
        DP_mult_204_n833), .CO(DP_mult_204_n826), .S(DP_mult_204_n827) );
  FA_X1 DP_mult_204_U619 ( .A(DP_mult_204_n846), .B(DP_mult_204_n848), .CI(
        DP_mult_204_n829), .CO(DP_mult_204_n824), .S(DP_mult_204_n825) );
  FA_X1 DP_mult_204_U617 ( .A(DP_mult_204_n840), .B(DP_mult_204_n825), .CI(
        DP_mult_204_n823), .CO(DP_mult_204_n820), .S(DP_mult_204_n821) );
  FA_X1 DP_mult_204_U616 ( .A(DP_mult_204_n1209), .B(DP_mult_204_n1363), .CI(
        DP_mult_204_n1930), .CO(DP_mult_204_n818), .S(DP_mult_204_n819) );
  FA_X1 DP_mult_204_U615 ( .A(DP_mult_204_n1231), .B(DP_mult_204_n1297), .CI(
        DP_mult_204_n1275), .CO(DP_mult_204_n816), .S(DP_mult_204_n817) );
  FA_X1 DP_mult_204_U614 ( .A(DP_mult_204_n1319), .B(DP_mult_204_n1253), .CI(
        DP_mult_204_n1341), .CO(DP_mult_204_n814), .S(DP_mult_204_n815) );
  FA_X1 DP_mult_204_U612 ( .A(DP_mult_204_n815), .B(DP_mult_204_n832), .CI(
        DP_mult_204_n817), .CO(DP_mult_204_n810), .S(DP_mult_204_n811) );
  FA_X1 DP_mult_204_U607 ( .A(DP_mult_204_n1340), .B(DP_mult_204_n1252), .CI(
        DP_mult_204_n803), .CO(DP_mult_204_n800), .S(DP_mult_204_n801) );
  FA_X1 DP_mult_204_U606 ( .A(DP_mult_204_n1208), .B(DP_mult_204_n1318), .CI(
        DP_mult_204_n1230), .CO(DP_mult_204_n798), .S(DP_mult_204_n799) );
  FA_X1 DP_mult_204_U604 ( .A(DP_mult_204_n814), .B(DP_mult_204_n816), .CI(
        DP_mult_204_n799), .CO(DP_mult_204_n794), .S(DP_mult_204_n795) );
  FA_X1 DP_mult_204_U603 ( .A(DP_mult_204_n801), .B(DP_mult_204_n812), .CI(
        DP_mult_204_n797), .CO(DP_mult_204_n792), .S(DP_mult_204_n793) );
  FA_X1 DP_mult_204_U601 ( .A(DP_mult_204_n806), .B(DP_mult_204_n793), .CI(
        DP_mult_204_n791), .CO(DP_mult_204_n788), .S(DP_mult_204_n789) );
  FA_X1 DP_mult_204_U600 ( .A(DP_mult_204_n1207), .B(DP_mult_204_n2154), .CI(
        DP_mult_204_n1251), .CO(DP_mult_204_n786), .S(DP_mult_204_n787) );
  FA_X1 DP_mult_204_U599 ( .A(DP_mult_204_n1273), .B(DP_mult_204_n1317), .CI(
        DP_mult_204_n1295), .CO(DP_mult_204_n784), .S(DP_mult_204_n785) );
  FA_X1 DP_mult_204_U598 ( .A(DP_mult_204_n1339), .B(DP_mult_204_n1229), .CI(
        DP_mult_204_n1362), .CO(DP_mult_204_n782), .S(DP_mult_204_n783) );
  FA_X1 DP_mult_204_U597 ( .A(DP_mult_204_n798), .B(DP_mult_204_n800), .CI(
        DP_mult_204_n785), .CO(DP_mult_204_n780), .S(DP_mult_204_n781) );
  FA_X1 DP_mult_204_U596 ( .A(DP_mult_204_n796), .B(DP_mult_204_n787), .CI(
        DP_mult_204_n783), .CO(DP_mult_204_n778), .S(DP_mult_204_n779) );
  FA_X1 DP_mult_204_U595 ( .A(DP_mult_204_n781), .B(DP_mult_204_n794), .CI(
        DP_mult_204_n792), .CO(DP_mult_204_n776), .S(DP_mult_204_n777) );
  FA_X1 DP_mult_204_U594 ( .A(DP_mult_204_n790), .B(DP_mult_204_n779), .CI(
        DP_mult_204_n777), .CO(DP_mult_204_n774), .S(DP_mult_204_n775) );
  FA_X1 DP_mult_204_U592 ( .A(DP_mult_204_n1316), .B(DP_mult_204_n1250), .CI(
        DP_mult_204_n773), .CO(DP_mult_204_n770), .S(DP_mult_204_n771) );
  FA_X1 DP_mult_204_U591 ( .A(DP_mult_204_n1294), .B(DP_mult_204_n1206), .CI(
        DP_mult_204_n1272), .CO(DP_mult_204_n768), .S(DP_mult_204_n769) );
  FA_X1 DP_mult_204_U590 ( .A(DP_mult_204_n786), .B(DP_mult_204_n1228), .CI(
        DP_mult_204_n784), .CO(DP_mult_204_n766), .S(DP_mult_204_n767) );
  FA_X1 DP_mult_204_U589 ( .A(DP_mult_204_n771), .B(DP_mult_204_n769), .CI(
        DP_mult_204_n782), .CO(DP_mult_204_n764), .S(DP_mult_204_n765) );
  FA_X1 DP_mult_204_U588 ( .A(DP_mult_204_n767), .B(DP_mult_204_n780), .CI(
        DP_mult_204_n778), .CO(DP_mult_204_n762), .S(DP_mult_204_n763) );
  FA_X1 DP_mult_204_U587 ( .A(DP_mult_204_n776), .B(DP_mult_204_n765), .CI(
        DP_mult_204_n763), .CO(DP_mult_204_n760), .S(DP_mult_204_n761) );
  FA_X1 DP_mult_204_U586 ( .A(DP_mult_204_n772), .B(DP_mult_204_n1205), .CI(
        DP_mult_204_n1227), .CO(DP_mult_204_n758), .S(DP_mult_204_n759) );
  FA_X1 DP_mult_204_U585 ( .A(DP_mult_204_n1249), .B(DP_mult_204_n1293), .CI(
        DP_mult_204_n1315), .CO(DP_mult_204_n756), .S(DP_mult_204_n757) );
  FA_X1 DP_mult_204_U584 ( .A(DP_mult_204_n1338), .B(DP_mult_204_n1271), .CI(
        DP_mult_204_n770), .CO(DP_mult_204_n754), .S(DP_mult_204_n755) );
  FA_X1 DP_mult_204_U583 ( .A(DP_mult_204_n757), .B(DP_mult_204_n768), .CI(
        DP_mult_204_n759), .CO(DP_mult_204_n752), .S(DP_mult_204_n753) );
  FA_X1 DP_mult_204_U582 ( .A(DP_mult_204_n755), .B(DP_mult_204_n766), .CI(
        DP_mult_204_n764), .CO(DP_mult_204_n750), .S(DP_mult_204_n751) );
  FA_X1 DP_mult_204_U581 ( .A(DP_mult_204_n762), .B(DP_mult_204_n753), .CI(
        DP_mult_204_n751), .CO(DP_mult_204_n748), .S(DP_mult_204_n749) );
  FA_X1 DP_mult_204_U579 ( .A(DP_mult_204_n1292), .B(DP_mult_204_n1248), .CI(
        DP_mult_204_n747), .CO(DP_mult_204_n744), .S(DP_mult_204_n745) );
  FA_X1 DP_mult_204_U578 ( .A(DP_mult_204_n1226), .B(DP_mult_204_n1204), .CI(
        DP_mult_204_n1270), .CO(DP_mult_204_n742), .S(DP_mult_204_n743) );
  FA_X1 DP_mult_204_U577 ( .A(DP_mult_204_n756), .B(DP_mult_204_n758), .CI(
        DP_mult_204_n743), .CO(DP_mult_204_n740), .S(DP_mult_204_n741) );
  FA_X1 DP_mult_204_U576 ( .A(DP_mult_204_n754), .B(DP_mult_204_n745), .CI(
        DP_mult_204_n752), .CO(DP_mult_204_n738), .S(DP_mult_204_n739) );
  FA_X1 DP_mult_204_U575 ( .A(DP_mult_204_n750), .B(DP_mult_204_n741), .CI(
        DP_mult_204_n739), .CO(DP_mult_204_n736), .S(DP_mult_204_n737) );
  FA_X1 DP_mult_204_U574 ( .A(DP_mult_204_n746), .B(DP_mult_204_n1203), .CI(
        DP_mult_204_n1247), .CO(DP_mult_204_n734), .S(DP_mult_204_n735) );
  FA_X1 DP_mult_204_U573 ( .A(DP_mult_204_n1225), .B(DP_mult_204_n1291), .CI(
        DP_mult_204_n1269), .CO(DP_mult_204_n732), .S(DP_mult_204_n733) );
  FA_X1 DP_mult_204_U572 ( .A(DP_mult_204_n744), .B(DP_mult_204_n1314), .CI(
        DP_mult_204_n742), .CO(DP_mult_204_n730), .S(DP_mult_204_n731) );
  FA_X1 DP_mult_204_U571 ( .A(DP_mult_204_n735), .B(DP_mult_204_n733), .CI(
        DP_mult_204_n740), .CO(DP_mult_204_n728), .S(DP_mult_204_n729) );
  FA_X1 DP_mult_204_U570 ( .A(DP_mult_204_n738), .B(DP_mult_204_n731), .CI(
        DP_mult_204_n729), .CO(DP_mult_204_n726), .S(DP_mult_204_n727) );
  FA_X1 DP_mult_204_U568 ( .A(DP_mult_204_n1268), .B(DP_mult_204_n1224), .CI(
        DP_mult_204_n725), .CO(DP_mult_204_n722), .S(DP_mult_204_n723) );
  FA_X1 DP_mult_204_U567 ( .A(DP_mult_204_n1202), .B(DP_mult_204_n1246), .CI(
        DP_mult_204_n734), .CO(DP_mult_204_n720), .S(DP_mult_204_n721) );
  FA_X1 DP_mult_204_U566 ( .A(DP_mult_204_n723), .B(DP_mult_204_n732), .CI(
        DP_mult_204_n730), .CO(DP_mult_204_n718), .S(DP_mult_204_n719) );
  FA_X1 DP_mult_204_U565 ( .A(DP_mult_204_n728), .B(DP_mult_204_n721), .CI(
        DP_mult_204_n719), .CO(DP_mult_204_n716), .S(DP_mult_204_n717) );
  FA_X1 DP_mult_204_U564 ( .A(DP_mult_204_n1267), .B(DP_mult_204_n1201), .CI(
        DP_mult_204_n724), .CO(DP_mult_204_n714), .S(DP_mult_204_n715) );
  FA_X1 DP_mult_204_U563 ( .A(DP_mult_204_n1245), .B(DP_mult_204_n1223), .CI(
        DP_mult_204_n1290), .CO(DP_mult_204_n712), .S(DP_mult_204_n713) );
  FA_X1 DP_mult_204_U562 ( .A(DP_mult_204_n715), .B(DP_mult_204_n722), .CI(
        DP_mult_204_n720), .CO(DP_mult_204_n710), .S(DP_mult_204_n711) );
  FA_X1 DP_mult_204_U561 ( .A(DP_mult_204_n718), .B(DP_mult_204_n713), .CI(
        DP_mult_204_n711), .CO(DP_mult_204_n708), .S(DP_mult_204_n709) );
  FA_X1 DP_mult_204_U559 ( .A(DP_mult_204_n1222), .B(DP_mult_204_n1200), .CI(
        DP_mult_204_n707), .CO(DP_mult_204_n704), .S(DP_mult_204_n705) );
  FA_X1 DP_mult_204_U558 ( .A(DP_mult_204_n714), .B(DP_mult_204_n1244), .CI(
        DP_mult_204_n705), .CO(DP_mult_204_n702), .S(DP_mult_204_n703) );
  FA_X1 DP_mult_204_U557 ( .A(DP_mult_204_n710), .B(DP_mult_204_n712), .CI(
        DP_mult_204_n703), .CO(DP_mult_204_n700), .S(DP_mult_204_n701) );
  FA_X1 DP_mult_204_U556 ( .A(DP_mult_204_n1221), .B(DP_mult_204_n1199), .CI(
        DP_mult_204_n706), .CO(DP_mult_204_n698), .S(DP_mult_204_n699) );
  FA_X1 DP_mult_204_U555 ( .A(DP_mult_204_n1266), .B(DP_mult_204_n1243), .CI(
        DP_mult_204_n704), .CO(DP_mult_204_n696), .S(DP_mult_204_n697) );
  FA_X1 DP_mult_204_U554 ( .A(DP_mult_204_n702), .B(DP_mult_204_n699), .CI(
        DP_mult_204_n697), .CO(DP_mult_204_n694), .S(DP_mult_204_n695) );
  FA_X1 DP_mult_204_U552 ( .A(DP_mult_204_n1198), .B(DP_mult_204_n1220), .CI(
        DP_mult_204_n693), .CO(DP_mult_204_n690), .S(DP_mult_204_n691) );
  FA_X1 DP_mult_204_U551 ( .A(DP_mult_204_n691), .B(DP_mult_204_n698), .CI(
        DP_mult_204_n696), .CO(DP_mult_204_n688), .S(DP_mult_204_n689) );
  FA_X1 DP_mult_204_U550 ( .A(DP_mult_204_n1219), .B(DP_mult_204_n692), .CI(
        DP_mult_204_n1197), .CO(DP_mult_204_n686), .S(DP_mult_204_n687) );
  FA_X1 DP_mult_204_U549 ( .A(DP_mult_204_n690), .B(DP_mult_204_n1242), .CI(
        DP_mult_204_n687), .CO(DP_mult_204_n684), .S(DP_mult_204_n685) );
  FA_X1 DP_mult_204_U547 ( .A(DP_mult_204_n683), .B(DP_mult_204_n1196), .CI(
        DP_mult_204_n686), .CO(DP_mult_204_n680), .S(DP_mult_204_n681) );
  FA_X1 DP_mult_204_U546 ( .A(DP_mult_204_n1195), .B(DP_mult_204_n682), .CI(
        DP_mult_204_n1218), .CO(DP_mult_204_n678), .S(DP_mult_204_n679) );
  INV_X2 DP_mult_206_U2832 ( .A(DP_pipe00[0]), .ZN(DP_mult_206_n2327) );
  INV_X1 DP_mult_206_U2831 ( .A(DP_coeffs_ff_int[2]), .ZN(DP_mult_206_n2323)
         );
  INV_X1 DP_mult_206_U2830 ( .A(DP_mult_206_n2323), .ZN(DP_mult_206_n2321) );
  INV_X1 DP_mult_206_U2829 ( .A(DP_coeffs_ff_int[4]), .ZN(DP_mult_206_n2318)
         );
  INV_X1 DP_mult_206_U2828 ( .A(DP_coeffs_ff_int[4]), .ZN(DP_mult_206_n2317)
         );
  INV_X1 DP_mult_206_U2827 ( .A(DP_mult_206_n2317), .ZN(DP_mult_206_n2316) );
  INV_X1 DP_mult_206_U2826 ( .A(DP_coeffs_ff_int[6]), .ZN(DP_mult_206_n2313)
         );
  INV_X1 DP_mult_206_U2825 ( .A(DP_mult_206_n2313), .ZN(DP_mult_206_n2312) );
  INV_X1 DP_mult_206_U2824 ( .A(DP_coeffs_ff_int[8]), .ZN(DP_mult_206_n2310)
         );
  INV_X1 DP_mult_206_U2823 ( .A(DP_mult_206_n2310), .ZN(DP_mult_206_n2309) );
  INV_X1 DP_mult_206_U2822 ( .A(DP_coeffs_ff_int[10]), .ZN(DP_mult_206_n2306)
         );
  INV_X1 DP_mult_206_U2821 ( .A(DP_coeffs_ff_int[10]), .ZN(DP_mult_206_n2305)
         );
  INV_X1 DP_mult_206_U2820 ( .A(DP_mult_206_n2306), .ZN(DP_mult_206_n2304) );
  INV_X1 DP_mult_206_U2819 ( .A(DP_coeffs_ff_int[12]), .ZN(DP_mult_206_n2301)
         );
  INV_X1 DP_mult_206_U2818 ( .A(DP_coeffs_ff_int[12]), .ZN(DP_mult_206_n2300)
         );
  INV_X1 DP_mult_206_U2817 ( .A(DP_mult_206_n2300), .ZN(DP_mult_206_n2299) );
  INV_X1 DP_mult_206_U2816 ( .A(DP_coeffs_ff_int[14]), .ZN(DP_mult_206_n2296)
         );
  INV_X1 DP_mult_206_U2815 ( .A(DP_coeffs_ff_int[14]), .ZN(DP_mult_206_n2295)
         );
  INV_X1 DP_mult_206_U2814 ( .A(DP_mult_206_n2296), .ZN(DP_mult_206_n2294) );
  INV_X1 DP_mult_206_U2813 ( .A(DP_coeffs_ff_int[16]), .ZN(DP_mult_206_n2291)
         );
  INV_X1 DP_mult_206_U2812 ( .A(DP_coeffs_ff_int[16]), .ZN(DP_mult_206_n2290)
         );
  INV_X1 DP_mult_206_U2811 ( .A(DP_coeffs_ff_int[18]), .ZN(DP_mult_206_n2286)
         );
  INV_X1 DP_mult_206_U2810 ( .A(DP_coeffs_ff_int[18]), .ZN(DP_mult_206_n2285)
         );
  INV_X1 DP_mult_206_U2809 ( .A(DP_mult_206_n2286), .ZN(DP_mult_206_n2284) );
  INV_X1 DP_mult_206_U2808 ( .A(DP_coeffs_ff_int[20]), .ZN(DP_mult_206_n2281)
         );
  INV_X1 DP_mult_206_U2807 ( .A(DP_coeffs_ff_int[20]), .ZN(DP_mult_206_n2280)
         );
  INV_X1 DP_mult_206_U2806 ( .A(DP_mult_206_n2281), .ZN(DP_mult_206_n2279) );
  INV_X1 DP_mult_206_U2805 ( .A(DP_coeffs_ff_int[22]), .ZN(DP_mult_206_n2276)
         );
  INV_X1 DP_mult_206_U2804 ( .A(DP_coeffs_ff_int[22]), .ZN(DP_mult_206_n2275)
         );
  INV_X1 DP_mult_206_U2803 ( .A(DP_mult_206_n1949), .ZN(DP_mult_206_n2274) );
  INV_X1 DP_mult_206_U2802 ( .A(DP_mult_206_n2120), .ZN(DP_mult_206_n2247) );
  INV_X2 DP_mult_206_U2801 ( .A(DP_mult_206_n2317), .ZN(DP_mult_206_n2315) );
  INV_X2 DP_mult_206_U2800 ( .A(DP_mult_206_n2197), .ZN(DP_mult_206_n2239) );
  XNOR2_X1 DP_mult_206_U2799 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2284), .ZN(
        DP_mult_206_n1713) );
  XNOR2_X1 DP_mult_206_U2798 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2284), .ZN(
        DP_mult_206_n1711) );
  XNOR2_X1 DP_mult_206_U2797 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2284), .ZN(
        DP_mult_206_n1719) );
  XNOR2_X1 DP_mult_206_U2796 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2283), .ZN(
        DP_mult_206_n1715) );
  XNOR2_X1 DP_mult_206_U2795 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2283), .ZN(
        DP_mult_206_n1709) );
  XNOR2_X1 DP_mult_206_U2794 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2283), .ZN(
        DP_mult_206_n1717) );
  OAI22_X1 DP_mult_206_U2793 ( .A1(DP_mult_206_n2236), .A2(DP_mult_206_n1693), 
        .B1(DP_mult_206_n1692), .B2(DP_mult_206_n2261), .ZN(DP_mult_206_n1396)
         );
  OAI22_X1 DP_mult_206_U2792 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n2291), 
        .B1(DP_mult_206_n1706), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1190)
         );
  OAI22_X1 DP_mult_206_U2791 ( .A1(DP_mult_206_n2134), .A2(DP_mult_206_n1684), 
        .B1(DP_mult_206_n2261), .B2(DP_mult_206_n1683), .ZN(DP_mult_206_n1387)
         );
  OAI22_X1 DP_mult_206_U2790 ( .A1(DP_mult_206_n2135), .A2(DP_mult_206_n1688), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1687), .ZN(DP_mult_206_n1391)
         );
  OAI22_X1 DP_mult_206_U2789 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1685), 
        .B1(DP_mult_206_n1684), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1388)
         );
  OAI22_X1 DP_mult_206_U2788 ( .A1(DP_mult_206_n2135), .A2(DP_mult_206_n1692), 
        .B1(DP_mult_206_n2261), .B2(DP_mult_206_n1691), .ZN(DP_mult_206_n1395)
         );
  OAI22_X1 DP_mult_206_U2787 ( .A1(DP_mult_206_n2134), .A2(DP_mult_206_n1687), 
        .B1(DP_mult_206_n1686), .B2(DP_mult_206_n2261), .ZN(DP_mult_206_n1390)
         );
  OAI22_X1 DP_mult_206_U2786 ( .A1(DP_mult_206_n2134), .A2(DP_mult_206_n1690), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1689), .ZN(DP_mult_206_n1393)
         );
  OAI22_X1 DP_mult_206_U2785 ( .A1(DP_mult_206_n2135), .A2(DP_mult_206_n1689), 
        .B1(DP_mult_206_n1688), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1392)
         );
  OAI22_X1 DP_mult_206_U2784 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1686), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1685), .ZN(DP_mult_206_n1389)
         );
  OAI22_X1 DP_mult_206_U2783 ( .A1(DP_mult_206_n2135), .A2(DP_mult_206_n1691), 
        .B1(DP_mult_206_n1690), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1394)
         );
  NAND2_X1 DP_mult_206_U2782 ( .A1(DP_mult_206_n775), .A2(DP_mult_206_n788), 
        .ZN(DP_mult_206_n474) );
  OAI21_X1 DP_mult_206_U2781 ( .B1(DP_mult_206_n2218), .B2(DP_mult_206_n398), 
        .A(DP_mult_206_n399), .ZN(DP_mult_206_n397) );
  OAI21_X1 DP_mult_206_U2780 ( .B1(DP_mult_206_n2218), .B2(DP_mult_206_n389), 
        .A(DP_mult_206_n390), .ZN(DP_mult_206_n388) );
  OAI21_X1 DP_mult_206_U2779 ( .B1(DP_mult_206_n301), .B2(DP_mult_206_n431), 
        .A(DP_mult_206_n432), .ZN(DP_mult_206_n430) );
  OAI21_X1 DP_mult_206_U2778 ( .B1(DP_mult_206_n301), .B2(DP_mult_206_n411), 
        .A(DP_mult_206_n412), .ZN(DP_mult_206_n410) );
  OAI21_X1 DP_mult_206_U2777 ( .B1(DP_mult_206_n301), .B2(DP_mult_206_n420), 
        .A(DP_mult_206_n421), .ZN(DP_mult_206_n419) );
  OAI21_X1 DP_mult_206_U2776 ( .B1(DP_mult_206_n2218), .B2(DP_mult_206_n343), 
        .A(DP_mult_206_n344), .ZN(DP_mult_206_n342) );
  OAI21_X1 DP_mult_206_U2775 ( .B1(DP_mult_206_n301), .B2(DP_mult_206_n380), 
        .A(DP_mult_206_n381), .ZN(DP_mult_206_n379) );
  OAI21_X1 DP_mult_206_U2774 ( .B1(DP_mult_206_n2219), .B2(DP_mult_206_n371), 
        .A(DP_mult_206_n372), .ZN(DP_mult_206_n370) );
  OAI21_X1 DP_mult_206_U2773 ( .B1(DP_mult_206_n2219), .B2(DP_mult_206_n354), 
        .A(DP_mult_206_n355), .ZN(DP_mult_206_n353) );
  OAI21_X1 DP_mult_206_U2772 ( .B1(DP_mult_206_n2219), .B2(DP_mult_206_n438), 
        .A(DP_mult_206_n439), .ZN(DP_mult_206_n437) );
  INV_X1 DP_mult_206_U2771 ( .A(DP_mult_206_n2219), .ZN(DP_mult_206_n448) );
  OAI21_X1 DP_mult_206_U2770 ( .B1(DP_mult_206_n2218), .B2(DP_mult_206_n326), 
        .A(DP_mult_206_n327), .ZN(DP_mult_206_n325) );
  XNOR2_X1 DP_mult_206_U2769 ( .A(DP_mult_206_n437), .B(DP_mult_206_n311), 
        .ZN(DP_pipe0_coeff_pipe00[13]) );
  AOI21_X1 DP_mult_206_U2768 ( .B1(DP_mult_206_n333), .B2(DP_mult_206_n2186), 
        .A(DP_mult_206_n2187), .ZN(DP_mult_206_n327) );
  NAND2_X1 DP_mult_206_U2767 ( .A1(DP_mult_206_n356), .A2(DP_mult_206_n2184), 
        .ZN(DP_mult_206_n347) );
  XNOR2_X1 DP_mult_206_U2766 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2277), .ZN(
        DP_mult_206_n1742) );
  XNOR2_X1 DP_mult_206_U2765 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2277), .ZN(
        DP_mult_206_n1738) );
  XNOR2_X1 DP_mult_206_U2764 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2277), .ZN(
        DP_mult_206_n1744) );
  XNOR2_X1 DP_mult_206_U2763 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2277), .ZN(
        DP_mult_206_n1736) );
  XNOR2_X1 DP_mult_206_U2762 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2277), .ZN(
        DP_mult_206_n1740) );
  OAI22_X1 DP_mult_206_U2761 ( .A1(DP_mult_206_n1724), .A2(DP_mult_206_n2160), 
        .B1(DP_mult_206_n1723), .B2(DP_mult_206_n2264), .ZN(DP_mult_206_n1426)
         );
  XNOR2_X1 DP_mult_206_U2760 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2277), .ZN(
        DP_mult_206_n1734) );
  OAI22_X1 DP_mult_206_U2759 ( .A1(DP_mult_206_n2159), .A2(DP_mult_206_n1719), 
        .B1(DP_mult_206_n2264), .B2(DP_mult_206_n1718), .ZN(DP_mult_206_n1421)
         );
  OAI22_X1 DP_mult_206_U2758 ( .A1(DP_mult_206_n2159), .A2(DP_mult_206_n1722), 
        .B1(DP_mult_206_n1721), .B2(DP_mult_206_n2263), .ZN(DP_mult_206_n1424)
         );
  OAI22_X1 DP_mult_206_U2757 ( .A1(DP_mult_206_n2159), .A2(DP_mult_206_n1729), 
        .B1(DP_mult_206_n2263), .B2(DP_mult_206_n1728), .ZN(DP_mult_206_n1431)
         );
  OAI22_X1 DP_mult_206_U2756 ( .A1(DP_mult_206_n2237), .A2(DP_mult_206_n1728), 
        .B1(DP_mult_206_n1727), .B2(DP_mult_206_n2264), .ZN(DP_mult_206_n1430)
         );
  OAI22_X1 DP_mult_206_U2755 ( .A1(DP_mult_206_n2237), .A2(DP_mult_206_n1723), 
        .B1(DP_mult_206_n2264), .B2(DP_mult_206_n1722), .ZN(DP_mult_206_n1425)
         );
  OAI22_X1 DP_mult_206_U2754 ( .A1(DP_mult_206_n2237), .A2(DP_mult_206_n1725), 
        .B1(DP_mult_206_n2264), .B2(DP_mult_206_n1724), .ZN(DP_mult_206_n1427)
         );
  OAI22_X1 DP_mult_206_U2753 ( .A1(DP_mult_206_n2159), .A2(DP_mult_206_n1730), 
        .B1(DP_mult_206_n1729), .B2(DP_mult_206_n2264), .ZN(DP_mult_206_n1432)
         );
  OAI22_X1 DP_mult_206_U2752 ( .A1(DP_mult_206_n2159), .A2(DP_mult_206_n1726), 
        .B1(DP_mult_206_n1725), .B2(DP_mult_206_n2263), .ZN(DP_mult_206_n1428)
         );
  OAI22_X1 DP_mult_206_U2751 ( .A1(DP_mult_206_n2160), .A2(DP_mult_206_n1721), 
        .B1(DP_mult_206_n2264), .B2(DP_mult_206_n1720), .ZN(DP_mult_206_n1423)
         );
  OAI22_X1 DP_mult_206_U2750 ( .A1(DP_mult_206_n2160), .A2(DP_mult_206_n1720), 
        .B1(DP_mult_206_n1719), .B2(DP_mult_206_n2263), .ZN(DP_mult_206_n1422)
         );
  OAI22_X1 DP_mult_206_U2749 ( .A1(DP_mult_206_n2237), .A2(DP_mult_206_n1727), 
        .B1(DP_mult_206_n2263), .B2(DP_mult_206_n1726), .ZN(DP_mult_206_n1429)
         );
  OAI21_X1 DP_mult_206_U2748 ( .B1(DP_mult_206_n536), .B2(DP_mult_206_n498), 
        .A(DP_mult_206_n499), .ZN(DP_mult_206_n497) );
  OAI21_X1 DP_mult_206_U2747 ( .B1(DP_mult_206_n536), .B2(DP_mult_206_n2090), 
        .A(DP_mult_206_n2212), .ZN(DP_mult_206_n504) );
  OAI21_X1 DP_mult_206_U2746 ( .B1(DP_mult_206_n536), .B2(DP_mult_206_n516), 
        .A(DP_mult_206_n517), .ZN(DP_mult_206_n515) );
  OAI21_X1 DP_mult_206_U2745 ( .B1(DP_mult_206_n536), .B2(DP_mult_206_n476), 
        .A(DP_mult_206_n477), .ZN(DP_mult_206_n475) );
  OAI21_X1 DP_mult_206_U2744 ( .B1(DP_mult_206_n536), .B2(DP_mult_206_n523), 
        .A(DP_mult_206_n524), .ZN(DP_mult_206_n522) );
  OAI21_X1 DP_mult_206_U2743 ( .B1(DP_mult_206_n536), .B2(DP_mult_206_n463), 
        .A(DP_mult_206_n464), .ZN(DP_mult_206_n462) );
  OAI21_X1 DP_mult_206_U2742 ( .B1(DP_mult_206_n536), .B2(DP_mult_206_n487), 
        .A(DP_mult_206_n488), .ZN(DP_mult_206_n486) );
  OAI21_X1 DP_mult_206_U2741 ( .B1(DP_mult_206_n536), .B2(DP_mult_206_n2167), 
        .A(DP_mult_206_n535), .ZN(DP_mult_206_n533) );
  XNOR2_X1 DP_mult_206_U2740 ( .A(DP_coeffs_ff_int[21]), .B(DP_mult_206_n2271), 
        .ZN(DP_mult_206_n253) );
  XNOR2_X1 DP_mult_206_U2739 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1769) );
  XNOR2_X1 DP_mult_206_U2738 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1765) );
  XNOR2_X1 DP_mult_206_U2737 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1761) );
  XNOR2_X1 DP_mult_206_U2736 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1767) );
  XNOR2_X1 DP_mult_206_U2735 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1759) );
  XNOR2_X1 DP_mult_206_U2734 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1763) );
  OAI22_X1 DP_mult_206_U2733 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1742), 
        .B1(DP_mult_206_n2266), .B2(DP_mult_206_n1741), .ZN(DP_mult_206_n1443)
         );
  OAI22_X1 DP_mult_206_U2732 ( .A1(DP_mult_206_n2240), .A2(DP_mult_206_n1737), 
        .B1(DP_mult_206_n1736), .B2(DP_mult_206_n2267), .ZN(DP_mult_206_n1438)
         );
  OAI22_X1 DP_mult_206_U2731 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1743), 
        .B1(DP_mult_206_n1742), .B2(DP_mult_206_n2267), .ZN(DP_mult_206_n1444)
         );
  OAI22_X1 DP_mult_206_U2730 ( .A1(DP_mult_206_n2240), .A2(DP_mult_206_n1734), 
        .B1(DP_mult_206_n2267), .B2(DP_mult_206_n1733), .ZN(DP_mult_206_n1435)
         );
  OAI22_X1 DP_mult_206_U2729 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1739), 
        .B1(DP_mult_206_n1738), .B2(DP_mult_206_n2266), .ZN(DP_mult_206_n1440)
         );
  OAI22_X1 DP_mult_206_U2728 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1735), 
        .B1(DP_mult_206_n1734), .B2(DP_mult_206_n2267), .ZN(DP_mult_206_n1436)
         );
  OAI22_X1 DP_mult_206_U2727 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1736), 
        .B1(DP_mult_206_n2266), .B2(DP_mult_206_n1735), .ZN(DP_mult_206_n1437)
         );
  OAI22_X1 DP_mult_206_U2726 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1740), 
        .B1(DP_mult_206_n2265), .B2(DP_mult_206_n1739), .ZN(DP_mult_206_n1441)
         );
  OAI22_X1 DP_mult_206_U2725 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1741), 
        .B1(DP_mult_206_n1740), .B2(DP_mult_206_n2265), .ZN(DP_mult_206_n1442)
         );
  OAI22_X1 DP_mult_206_U2724 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1738), 
        .B1(DP_mult_206_n2265), .B2(DP_mult_206_n1737), .ZN(DP_mult_206_n1439)
         );
  OAI22_X1 DP_mult_206_U2723 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n2280), 
        .B1(DP_mult_206_n1756), .B2(DP_mult_206_n2266), .ZN(DP_mult_206_n1192)
         );
  INV_X1 DP_mult_206_U2722 ( .A(DP_mult_206_n490), .ZN(DP_mult_206_n492) );
  AOI21_X1 DP_mult_206_U2721 ( .B1(DP_mult_206_n508), .B2(DP_mult_206_n489), 
        .A(DP_mult_206_n1935), .ZN(DP_mult_206_n488) );
  XNOR2_X1 DP_mult_206_U2720 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2299), .ZN(
        DP_mult_206_n1642) );
  XNOR2_X1 DP_mult_206_U2719 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2297), .ZN(
        DP_mult_206_n1640) );
  XNOR2_X1 DP_mult_206_U2718 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2298), .ZN(
        DP_mult_206_n1644) );
  XNOR2_X1 DP_mult_206_U2717 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2297), .ZN(
        DP_mult_206_n1638) );
  OAI22_X1 DP_mult_206_U2716 ( .A1(DP_mult_206_n2230), .A2(DP_mult_206_n1608), 
        .B1(DP_mult_206_n1607), .B2(DP_mult_206_n2257), .ZN(DP_mult_206_n746)
         );
  XNOR2_X1 DP_mult_206_U2715 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2299), .ZN(
        DP_mult_206_n1634) );
  XNOR2_X1 DP_mult_206_U2714 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2299), .ZN(
        DP_mult_206_n1636) );
  OAI22_X1 DP_mult_206_U2713 ( .A1(DP_mult_206_n2229), .A2(DP_mult_206_n1614), 
        .B1(DP_mult_206_n1613), .B2(DP_mult_206_n2257), .ZN(DP_mult_206_n1320)
         );
  OAI22_X1 DP_mult_206_U2712 ( .A1(DP_mult_206_n2229), .A2(DP_mult_206_n1616), 
        .B1(DP_mult_206_n1615), .B2(DP_mult_206_n2258), .ZN(DP_mult_206_n1322)
         );
  OAI22_X1 DP_mult_206_U2711 ( .A1(DP_mult_206_n2229), .A2(DP_mult_206_n1618), 
        .B1(DP_mult_206_n1617), .B2(DP_mult_206_n2258), .ZN(DP_mult_206_n1324)
         );
  OAI22_X1 DP_mult_206_U2710 ( .A1(DP_mult_206_n2060), .A2(DP_mult_206_n2306), 
        .B1(DP_mult_206_n1631), .B2(DP_mult_206_n2258), .ZN(DP_mult_206_n1187)
         );
  OAI22_X1 DP_mult_206_U2709 ( .A1(DP_mult_206_n2061), .A2(DP_mult_206_n1609), 
        .B1(DP_mult_206_n2257), .B2(DP_mult_206_n1608), .ZN(DP_mult_206_n1315)
         );
  INV_X1 DP_mult_206_U2708 ( .A(DP_mult_206_n746), .ZN(DP_mult_206_n747) );
  OAI22_X1 DP_mult_206_U2707 ( .A1(DP_mult_206_n2230), .A2(DP_mult_206_n1611), 
        .B1(DP_mult_206_n2257), .B2(DP_mult_206_n1610), .ZN(DP_mult_206_n1317)
         );
  OAI22_X1 DP_mult_206_U2706 ( .A1(DP_mult_206_n2230), .A2(DP_mult_206_n1615), 
        .B1(DP_mult_206_n2257), .B2(DP_mult_206_n1614), .ZN(DP_mult_206_n1321)
         );
  OAI22_X1 DP_mult_206_U2705 ( .A1(DP_mult_206_n2060), .A2(DP_mult_206_n1617), 
        .B1(DP_mult_206_n2258), .B2(DP_mult_206_n1616), .ZN(DP_mult_206_n1323)
         );
  OAI22_X1 DP_mult_206_U2704 ( .A1(DP_mult_206_n2060), .A2(DP_mult_206_n1610), 
        .B1(DP_mult_206_n1609), .B2(DP_mult_206_n2258), .ZN(DP_mult_206_n1316)
         );
  OAI22_X1 DP_mult_206_U2703 ( .A1(DP_mult_206_n2060), .A2(DP_mult_206_n1612), 
        .B1(DP_mult_206_n1611), .B2(DP_mult_206_n2258), .ZN(DP_mult_206_n1318)
         );
  OAI22_X1 DP_mult_206_U2702 ( .A1(DP_mult_206_n2061), .A2(DP_mult_206_n1613), 
        .B1(DP_mult_206_n2258), .B2(DP_mult_206_n1612), .ZN(DP_mult_206_n1319)
         );
  NAND2_X1 DP_mult_206_U2701 ( .A1(DP_mult_206_n717), .A2(DP_mult_206_n726), 
        .ZN(DP_mult_206_n418) );
  NAND2_X1 DP_mult_206_U2700 ( .A1(DP_mult_206_n345), .A2(DP_mult_206_n2185), 
        .ZN(DP_mult_206_n336) );
  INV_X1 DP_mult_206_U2699 ( .A(DP_mult_206_n345), .ZN(DP_mult_206_n343) );
  INV_X1 DP_mult_206_U2698 ( .A(DP_mult_206_n325), .ZN(
        DP_pipe0_coeff_pipe00[23]) );
  OAI21_X1 DP_mult_206_U2697 ( .B1(DP_mult_206_n506), .B2(DP_mult_206_n452), 
        .A(DP_mult_206_n453), .ZN(DP_mult_206_n451) );
  OAI22_X1 DP_mult_206_U2696 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n2300), 
        .B1(DP_mult_206_n1656), .B2(DP_mult_206_n2259), .ZN(DP_mult_206_n1188)
         );
  XNOR2_X1 DP_mult_206_U2695 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2302), .ZN(
        DP_mult_206_n1615) );
  XNOR2_X1 DP_mult_206_U2694 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2302), .ZN(
        DP_mult_206_n1619) );
  XNOR2_X1 DP_mult_206_U2693 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2302), .ZN(
        DP_mult_206_n1617) );
  XNOR2_X1 DP_mult_206_U2692 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2302), .ZN(
        DP_mult_206_n1613) );
  XNOR2_X1 DP_mult_206_U2691 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2007), .ZN(
        DP_mult_206_n1609) );
  OAI22_X1 DP_mult_206_U2690 ( .A1(DP_mult_206_n1988), .A2(DP_mult_206_n1605), 
        .B1(DP_mult_206_n1604), .B2(DP_mult_206_n2255), .ZN(DP_mult_206_n1312)
         );
  XNOR2_X1 DP_mult_206_U2689 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2007), .ZN(
        DP_mult_206_n1611) );
  OAI22_X1 DP_mult_206_U2688 ( .A1(DP_mult_206_n2024), .A2(DP_mult_206_n1599), 
        .B1(DP_mult_206_n1598), .B2(DP_mult_206_n2256), .ZN(DP_mult_206_n1306)
         );
  OAI22_X1 DP_mult_206_U2687 ( .A1(DP_mult_206_n1987), .A2(DP_mult_206_n1604), 
        .B1(DP_mult_206_n2256), .B2(DP_mult_206_n1603), .ZN(DP_mult_206_n1311)
         );
  OAI22_X1 DP_mult_206_U2686 ( .A1(DP_mult_206_n2227), .A2(DP_mult_206_n1595), 
        .B1(DP_mult_206_n1594), .B2(DP_mult_206_n2256), .ZN(DP_mult_206_n1302)
         );
  OAI22_X1 DP_mult_206_U2685 ( .A1(DP_mult_206_n2024), .A2(DP_mult_206_n1603), 
        .B1(DP_mult_206_n1602), .B2(DP_mult_206_n2255), .ZN(DP_mult_206_n1310)
         );
  OAI22_X1 DP_mult_206_U2684 ( .A1(DP_mult_206_n2227), .A2(DP_mult_206_n1597), 
        .B1(DP_mult_206_n1596), .B2(DP_mult_206_n2256), .ZN(DP_mult_206_n1304)
         );
  OAI22_X1 DP_mult_206_U2683 ( .A1(DP_mult_206_n2024), .A2(DP_mult_206_n1598), 
        .B1(DP_mult_206_n2256), .B2(DP_mult_206_n1597), .ZN(DP_mult_206_n1305)
         );
  OAI22_X1 DP_mult_206_U2682 ( .A1(DP_mult_206_n1987), .A2(DP_mult_206_n1596), 
        .B1(DP_mult_206_n2255), .B2(DP_mult_206_n1595), .ZN(DP_mult_206_n1303)
         );
  OAI22_X1 DP_mult_206_U2681 ( .A1(DP_mult_206_n1987), .A2(DP_mult_206_n1594), 
        .B1(DP_mult_206_n2255), .B2(DP_mult_206_n1593), .ZN(DP_mult_206_n1301)
         );
  OAI22_X1 DP_mult_206_U2680 ( .A1(DP_mult_206_n1987), .A2(DP_mult_206_n1601), 
        .B1(DP_mult_206_n1600), .B2(DP_mult_206_n2255), .ZN(DP_mult_206_n1308)
         );
  OAI22_X1 DP_mult_206_U2679 ( .A1(DP_mult_206_n2227), .A2(DP_mult_206_n1600), 
        .B1(DP_mult_206_n2255), .B2(DP_mult_206_n1599), .ZN(DP_mult_206_n1307)
         );
  OAI22_X1 DP_mult_206_U2678 ( .A1(DP_mult_206_n2024), .A2(DP_mult_206_n1602), 
        .B1(DP_mult_206_n2256), .B2(DP_mult_206_n1601), .ZN(DP_mult_206_n1309)
         );
  OAI21_X1 DP_mult_206_U2677 ( .B1(DP_mult_206_n572), .B2(DP_mult_206_n569), 
        .A(DP_mult_206_n570), .ZN(DP_mult_206_n568) );
  XNOR2_X1 DP_mult_206_U2676 ( .A(DP_mult_206_n430), .B(DP_mult_206_n310), 
        .ZN(DP_pipe0_coeff_pipe00[14]) );
  AOI21_X1 DP_mult_206_U2675 ( .B1(DP_mult_206_n540), .B2(DP_mult_206_n553), 
        .A(DP_mult_206_n541), .ZN(DP_mult_206_n539) );
  NAND2_X1 DP_mult_206_U2674 ( .A1(DP_mult_206_n540), .A2(DP_mult_206_n552), 
        .ZN(DP_mult_206_n538) );
  OAI22_X1 DP_mult_206_U2673 ( .A1(DP_mult_206_n2126), .A2(DP_mult_206_n1527), 
        .B1(DP_mult_206_n2247), .B2(DP_mult_206_n1526), .ZN(DP_mult_206_n1237)
         );
  OAI22_X1 DP_mult_206_U2672 ( .A1(DP_mult_206_n2221), .A2(DP_mult_206_n1528), 
        .B1(DP_mult_206_n1527), .B2(DP_mult_206_n2246), .ZN(DP_mult_206_n1238)
         );
  OAI22_X1 DP_mult_206_U2671 ( .A1(DP_mult_206_n2127), .A2(DP_mult_206_n1530), 
        .B1(DP_mult_206_n1529), .B2(DP_mult_206_n2048), .ZN(DP_mult_206_n1240)
         );
  OAI22_X1 DP_mult_206_U2670 ( .A1(DP_mult_206_n2221), .A2(DP_mult_206_n1526), 
        .B1(DP_mult_206_n1525), .B2(DP_mult_206_n2247), .ZN(DP_mult_206_n1236)
         );
  OAI22_X1 DP_mult_206_U2669 ( .A1(DP_mult_206_n2126), .A2(DP_mult_206_n1524), 
        .B1(DP_mult_206_n1523), .B2(DP_mult_206_n2246), .ZN(DP_mult_206_n1234)
         );
  OAI22_X1 DP_mult_206_U2668 ( .A1(DP_mult_206_n2222), .A2(DP_mult_206_n1529), 
        .B1(DP_mult_206_n2048), .B2(DP_mult_206_n1528), .ZN(DP_mult_206_n1239)
         );
  OAI22_X1 DP_mult_206_U2667 ( .A1(DP_mult_206_n2126), .A2(DP_mult_206_n1525), 
        .B1(DP_mult_206_n2246), .B2(DP_mult_206_n1524), .ZN(DP_mult_206_n1235)
         );
  OAI22_X1 DP_mult_206_U2666 ( .A1(DP_mult_206_n2222), .A2(DP_mult_206_n1523), 
        .B1(DP_mult_206_n2247), .B2(DP_mult_206_n1522), .ZN(DP_mult_206_n1233)
         );
  OAI22_X1 DP_mult_206_U2665 ( .A1(DP_mult_206_n2222), .A2(DP_mult_206_n1519), 
        .B1(DP_mult_206_n2247), .B2(DP_mult_206_n1518), .ZN(DP_mult_206_n1229)
         );
  OAI22_X1 DP_mult_206_U2664 ( .A1(DP_mult_206_n2127), .A2(DP_mult_206_n1520), 
        .B1(DP_mult_206_n1519), .B2(DP_mult_206_n2048), .ZN(DP_mult_206_n1230)
         );
  OAI22_X1 DP_mult_206_U2663 ( .A1(DP_mult_206_n2127), .A2(DP_mult_206_n1521), 
        .B1(DP_mult_206_n2048), .B2(DP_mult_206_n1520), .ZN(DP_mult_206_n1231)
         );
  OAI22_X1 DP_mult_206_U2662 ( .A1(DP_mult_206_n2222), .A2(DP_mult_206_n1522), 
        .B1(DP_mult_206_n1521), .B2(DP_mult_206_n2247), .ZN(DP_mult_206_n1232)
         );
  XNOR2_X1 DP_mult_206_U2661 ( .A(DP_mult_206_n419), .B(DP_mult_206_n309), 
        .ZN(DP_pipe0_coeff_pipe00[15]) );
  OAI22_X1 DP_mult_206_U2660 ( .A1(DP_mult_206_n1948), .A2(DP_mult_206_n1498), 
        .B1(DP_mult_206_n1986), .B2(DP_mult_206_n1497), .ZN(DP_mult_206_n1209)
         );
  OAI22_X1 DP_mult_206_U2659 ( .A1(DP_mult_206_n1948), .A2(DP_mult_206_n1504), 
        .B1(DP_mult_206_n1986), .B2(DP_mult_206_n1503), .ZN(DP_mult_206_n1215)
         );
  OAI22_X1 DP_mult_206_U2658 ( .A1(DP_mult_206_n1948), .A2(DP_mult_206_n1505), 
        .B1(DP_mult_206_n1504), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n1216)
         );
  OAI22_X1 DP_mult_206_U2657 ( .A1(DP_mult_206_n1948), .A2(DP_mult_206_n1499), 
        .B1(DP_mult_206_n1498), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n1210)
         );
  OAI22_X1 DP_mult_206_U2656 ( .A1(DP_mult_206_n1948), .A2(DP_mult_206_n1503), 
        .B1(DP_mult_206_n1502), .B2(DP_mult_206_n1986), .ZN(DP_mult_206_n1214)
         );
  OAI22_X1 DP_mult_206_U2655 ( .A1(DP_mult_206_n2220), .A2(DP_mult_206_n1494), 
        .B1(DP_mult_206_n1986), .B2(DP_mult_206_n1493), .ZN(DP_mult_206_n1205)
         );
  OAI22_X1 DP_mult_206_U2654 ( .A1(DP_mult_206_n1948), .A2(DP_mult_206_n1501), 
        .B1(DP_mult_206_n1500), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n1212)
         );
  OAI22_X1 DP_mult_206_U2653 ( .A1(DP_mult_206_n1948), .A2(DP_mult_206_n1502), 
        .B1(DP_mult_206_n2244), .B2(DP_mult_206_n1501), .ZN(DP_mult_206_n1213)
         );
  OAI22_X1 DP_mult_206_U2652 ( .A1(DP_mult_206_n2220), .A2(DP_mult_206_n1500), 
        .B1(DP_mult_206_n1986), .B2(DP_mult_206_n1499), .ZN(DP_mult_206_n1211)
         );
  OAI22_X1 DP_mult_206_U2651 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1495), 
        .B1(DP_mult_206_n1494), .B2(DP_mult_206_n1986), .ZN(DP_mult_206_n1206)
         );
  OAI22_X1 DP_mult_206_U2650 ( .A1(DP_mult_206_n2220), .A2(DP_mult_206_n1496), 
        .B1(DP_mult_206_n2244), .B2(DP_mult_206_n1495), .ZN(DP_mult_206_n1207)
         );
  OAI22_X1 DP_mult_206_U2649 ( .A1(DP_mult_206_n2220), .A2(DP_mult_206_n1497), 
        .B1(DP_mult_206_n1496), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n1208)
         );
  XNOR2_X1 DP_mult_206_U2648 ( .A(DP_mult_206_n410), .B(DP_mult_206_n308), 
        .ZN(DP_pipe0_coeff_pipe00[16]) );
  XNOR2_X1 DP_mult_206_U2647 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1540) );
  XNOR2_X1 DP_mult_206_U2646 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1544) );
  XNOR2_X1 DP_mult_206_U2645 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1538) );
  XNOR2_X1 DP_mult_206_U2644 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1542) );
  OR2_X1 DP_mult_206_U2643 ( .A1(DP_mult_206_n1237), .A2(DP_mult_206_n1215), 
        .ZN(DP_mult_206_n938) );
  XNOR2_X1 DP_mult_206_U2642 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1534) );
  XNOR2_X1 DP_mult_206_U2641 ( .A(DP_mult_206_n1237), .B(DP_mult_206_n1215), 
        .ZN(DP_mult_206_n939) );
  XNOR2_X1 DP_mult_206_U2640 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1536) );
  XNOR2_X1 DP_mult_206_U2639 ( .A(DP_mult_206_n397), .B(DP_mult_206_n307), 
        .ZN(DP_pipe0_coeff_pipe00[17]) );
  XNOR2_X1 DP_mult_206_U2638 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2287), .ZN(
        DP_mult_206_n1692) );
  XNOR2_X1 DP_mult_206_U2637 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2288), .ZN(
        DP_mult_206_n1694) );
  XNOR2_X1 DP_mult_206_U2636 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2288), .ZN(
        DP_mult_206_n1684) );
  XNOR2_X1 DP_mult_206_U2635 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2287), .ZN(
        DP_mult_206_n1686) );
  XNOR2_X1 DP_mult_206_U2634 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2287), .ZN(
        DP_mult_206_n1690) );
  XNOR2_X1 DP_mult_206_U2633 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2287), .ZN(
        DP_mult_206_n1688) );
  OAI22_X1 DP_mult_206_U2632 ( .A1(DP_mult_206_n1941), .A2(DP_mult_206_n1668), 
        .B1(DP_mult_206_n1667), .B2(DP_mult_206_n2201), .ZN(DP_mult_206_n1372)
         );
  OAI22_X1 DP_mult_206_U2631 ( .A1(DP_mult_206_n1942), .A2(DP_mult_206_n1659), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1658), .ZN(DP_mult_206_n1363)
         );
  OAI22_X1 DP_mult_206_U2630 ( .A1(DP_mult_206_n2234), .A2(DP_mult_206_n1662), 
        .B1(DP_mult_206_n1661), .B2(DP_mult_206_n2201), .ZN(DP_mult_206_n1366)
         );
  OAI22_X1 DP_mult_206_U2629 ( .A1(DP_mult_206_n1941), .A2(DP_mult_206_n1658), 
        .B1(DP_mult_206_n1657), .B2(DP_mult_206_n2201), .ZN(DP_mult_206_n802)
         );
  OAI22_X1 DP_mult_206_U2628 ( .A1(DP_mult_206_n1942), .A2(DP_mult_206_n1665), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1664), .ZN(DP_mult_206_n1369)
         );
  OAI22_X1 DP_mult_206_U2627 ( .A1(DP_mult_206_n2234), .A2(DP_mult_206_n1664), 
        .B1(DP_mult_206_n1663), .B2(DP_mult_206_n2201), .ZN(DP_mult_206_n1368)
         );
  OAI22_X1 DP_mult_206_U2626 ( .A1(DP_mult_206_n1941), .A2(DP_mult_206_n1667), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1666), .ZN(DP_mult_206_n1371)
         );
  OAI22_X1 DP_mult_206_U2625 ( .A1(DP_mult_206_n2233), .A2(DP_mult_206_n2295), 
        .B1(DP_mult_206_n1681), .B2(DP_mult_206_n2201), .ZN(DP_mult_206_n1189)
         );
  OAI22_X1 DP_mult_206_U2624 ( .A1(DP_mult_206_n1941), .A2(DP_mult_206_n1663), 
        .B1(DP_mult_206_n2201), .B2(DP_mult_206_n1662), .ZN(DP_mult_206_n1367)
         );
  OAI22_X1 DP_mult_206_U2623 ( .A1(DP_mult_206_n2233), .A2(DP_mult_206_n1660), 
        .B1(DP_mult_206_n1659), .B2(DP_mult_206_n2201), .ZN(DP_mult_206_n1364)
         );
  OAI22_X1 DP_mult_206_U2622 ( .A1(DP_mult_206_n1941), .A2(DP_mult_206_n1661), 
        .B1(DP_mult_206_n2201), .B2(DP_mult_206_n1660), .ZN(DP_mult_206_n1365)
         );
  XNOR2_X1 DP_mult_206_U2621 ( .A(DP_mult_206_n388), .B(DP_mult_206_n306), 
        .ZN(DP_pipe0_coeff_pipe00[18]) );
  OAI22_X1 DP_mult_206_U2620 ( .A1(DP_mult_206_n1948), .A2(DP_mult_206_n2326), 
        .B1(DP_mult_206_n1506), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n1182)
         );
  OAI22_X1 DP_mult_206_U2619 ( .A1(DP_mult_206_n2220), .A2(DP_mult_206_n1493), 
        .B1(DP_mult_206_n1492), .B2(DP_mult_206_n1986), .ZN(DP_mult_206_n1204)
         );
  OAI22_X1 DP_mult_206_U2618 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1489), 
        .B1(DP_mult_206_n1488), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n1200)
         );
  OAI22_X1 DP_mult_206_U2617 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1492), 
        .B1(DP_mult_206_n2244), .B2(DP_mult_206_n1491), .ZN(DP_mult_206_n1203)
         );
  OAI22_X1 DP_mult_206_U2616 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1486), 
        .B1(DP_mult_206_n2244), .B2(DP_mult_206_n1485), .ZN(DP_mult_206_n1197)
         );
  OAI22_X1 DP_mult_206_U2615 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1490), 
        .B1(DP_mult_206_n1986), .B2(DP_mult_206_n1489), .ZN(DP_mult_206_n1201)
         );
  OAI22_X1 DP_mult_206_U2614 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1487), 
        .B1(DP_mult_206_n1486), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n1198)
         );
  OAI22_X1 DP_mult_206_U2613 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1488), 
        .B1(DP_mult_206_n1986), .B2(DP_mult_206_n1487), .ZN(DP_mult_206_n1199)
         );
  OAI22_X1 DP_mult_206_U2612 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1491), 
        .B1(DP_mult_206_n1490), .B2(DP_mult_206_n1986), .ZN(DP_mult_206_n1202)
         );
  OAI22_X1 DP_mult_206_U2611 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1485), 
        .B1(DP_mult_206_n1484), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n1196)
         );
  OAI22_X1 DP_mult_206_U2610 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1484), 
        .B1(DP_mult_206_n1986), .B2(DP_mult_206_n1483), .ZN(DP_mult_206_n1195)
         );
  OAI22_X1 DP_mult_206_U2609 ( .A1(DP_mult_206_n2104), .A2(DP_mult_206_n1483), 
        .B1(DP_mult_206_n1482), .B2(DP_mult_206_n2244), .ZN(DP_mult_206_n676)
         );
  OAI21_X1 DP_mult_206_U2608 ( .B1(DP_mult_206_n421), .B2(DP_mult_206_n402), 
        .A(DP_mult_206_n405), .ZN(DP_mult_206_n401) );
  OAI21_X1 DP_mult_206_U2607 ( .B1(DP_mult_206_n421), .B2(DP_mult_206_n347), 
        .A(DP_mult_206_n348), .ZN(DP_mult_206_n346) );
  INV_X1 DP_mult_206_U2606 ( .A(DP_mult_206_n421), .ZN(DP_mult_206_n423) );
  XNOR2_X1 DP_mult_206_U2605 ( .A(DP_mult_206_n370), .B(DP_mult_206_n304), 
        .ZN(DP_pipe0_coeff_pipe00[20]) );
  NAND2_X1 DP_mult_206_U2604 ( .A1(DP_mult_206_n1812), .A2(DP_mult_206_n2133), 
        .ZN(DP_mult_206_n285) );
  OAI22_X1 DP_mult_206_U2603 ( .A1(DP_mult_206_n2231), .A2(DP_mult_206_n1643), 
        .B1(DP_mult_206_n1642), .B2(DP_mult_206_n2259), .ZN(DP_mult_206_n1348)
         );
  OAI22_X1 DP_mult_206_U2602 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1655), 
        .B1(DP_mult_206_n1654), .B2(DP_mult_206_n2056), .ZN(DP_mult_206_n1360)
         );
  OAI22_X1 DP_mult_206_U2601 ( .A1(DP_mult_206_n2231), .A2(DP_mult_206_n1641), 
        .B1(DP_mult_206_n1640), .B2(DP_mult_206_n2259), .ZN(DP_mult_206_n1346)
         );
  OAI22_X1 DP_mult_206_U2600 ( .A1(DP_mult_206_n2231), .A2(DP_mult_206_n1642), 
        .B1(DP_mult_206_n2259), .B2(DP_mult_206_n1641), .ZN(DP_mult_206_n1347)
         );
  OAI22_X1 DP_mult_206_U2599 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1633), 
        .B1(DP_mult_206_n1632), .B2(DP_mult_206_n2259), .ZN(DP_mult_206_n772)
         );
  OAI22_X1 DP_mult_206_U2598 ( .A1(DP_mult_206_n2231), .A2(DP_mult_206_n1638), 
        .B1(DP_mult_206_n2259), .B2(DP_mult_206_n1637), .ZN(DP_mult_206_n1343)
         );
  OAI22_X1 DP_mult_206_U2597 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1640), 
        .B1(DP_mult_206_n2056), .B2(DP_mult_206_n1639), .ZN(DP_mult_206_n1345)
         );
  OAI22_X1 DP_mult_206_U2596 ( .A1(DP_mult_206_n2231), .A2(DP_mult_206_n1639), 
        .B1(DP_mult_206_n1638), .B2(DP_mult_206_n2259), .ZN(DP_mult_206_n1344)
         );
  OAI22_X1 DP_mult_206_U2595 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1653), 
        .B1(DP_mult_206_n1652), .B2(DP_mult_206_n2259), .ZN(DP_mult_206_n1358)
         );
  OAI22_X1 DP_mult_206_U2594 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1635), 
        .B1(DP_mult_206_n1634), .B2(DP_mult_206_n2259), .ZN(DP_mult_206_n1340)
         );
  OAI22_X1 DP_mult_206_U2593 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1634), 
        .B1(DP_mult_206_n2259), .B2(DP_mult_206_n1633), .ZN(DP_mult_206_n1339)
         );
  OAI22_X1 DP_mult_206_U2592 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1636), 
        .B1(DP_mult_206_n2259), .B2(DP_mult_206_n1635), .ZN(DP_mult_206_n1341)
         );
  OAI22_X1 DP_mult_206_U2591 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1637), 
        .B1(DP_mult_206_n1636), .B2(DP_mult_206_n2056), .ZN(DP_mult_206_n1342)
         );
  OAI22_X1 DP_mult_206_U2590 ( .A1(DP_mult_206_n2226), .A2(DP_mult_206_n1568), 
        .B1(DP_mult_206_n1567), .B2(DP_mult_206_n2252), .ZN(DP_mult_206_n1276)
         );
  OAI22_X1 DP_mult_206_U2589 ( .A1(DP_mult_206_n2202), .A2(DP_mult_206_n1558), 
        .B1(DP_mult_206_n1557), .B2(DP_mult_206_n2253), .ZN(DP_mult_206_n706)
         );
  OAI22_X1 DP_mult_206_U2588 ( .A1(DP_mult_206_n2169), .A2(DP_mult_206_n1565), 
        .B1(DP_mult_206_n2253), .B2(DP_mult_206_n1564), .ZN(DP_mult_206_n1273)
         );
  OAI22_X1 DP_mult_206_U2587 ( .A1(DP_mult_206_n2168), .A2(DP_mult_206_n1578), 
        .B1(DP_mult_206_n1577), .B2(DP_mult_206_n2253), .ZN(DP_mult_206_n1286)
         );
  OAI22_X1 DP_mult_206_U2586 ( .A1(DP_mult_206_n2226), .A2(DP_mult_206_n1580), 
        .B1(DP_mult_206_n1579), .B2(DP_mult_206_n2252), .ZN(DP_mult_206_n1288)
         );
  OAI22_X1 DP_mult_206_U2585 ( .A1(DP_mult_206_n2168), .A2(DP_mult_206_n2313), 
        .B1(DP_mult_206_n1581), .B2(DP_mult_206_n2252), .ZN(DP_mult_206_n1185)
         );
  OAI22_X1 DP_mult_206_U2584 ( .A1(DP_mult_206_n2168), .A2(DP_mult_206_n1562), 
        .B1(DP_mult_206_n1561), .B2(DP_mult_206_n2253), .ZN(DP_mult_206_n1270)
         );
  OAI22_X1 DP_mult_206_U2583 ( .A1(DP_mult_206_n2168), .A2(DP_mult_206_n1564), 
        .B1(DP_mult_206_n1563), .B2(DP_mult_206_n2253), .ZN(DP_mult_206_n1272)
         );
  OAI22_X1 DP_mult_206_U2582 ( .A1(DP_mult_206_n2168), .A2(DP_mult_206_n1566), 
        .B1(DP_mult_206_n1565), .B2(DP_mult_206_n2253), .ZN(DP_mult_206_n1274)
         );
  OAI22_X1 DP_mult_206_U2581 ( .A1(DP_mult_206_n2169), .A2(DP_mult_206_n1567), 
        .B1(DP_mult_206_n2252), .B2(DP_mult_206_n1566), .ZN(DP_mult_206_n1275)
         );
  OAI22_X1 DP_mult_206_U2580 ( .A1(DP_mult_206_n2202), .A2(DP_mult_206_n1559), 
        .B1(DP_mult_206_n2253), .B2(DP_mult_206_n1558), .ZN(DP_mult_206_n1267)
         );
  OAI22_X1 DP_mult_206_U2579 ( .A1(DP_mult_206_n2226), .A2(DP_mult_206_n1560), 
        .B1(DP_mult_206_n1559), .B2(DP_mult_206_n2252), .ZN(DP_mult_206_n1268)
         );
  OAI22_X1 DP_mult_206_U2578 ( .A1(DP_mult_206_n2169), .A2(DP_mult_206_n1561), 
        .B1(DP_mult_206_n2252), .B2(DP_mult_206_n1560), .ZN(DP_mult_206_n1269)
         );
  OAI22_X1 DP_mult_206_U2577 ( .A1(DP_mult_206_n2168), .A2(DP_mult_206_n1563), 
        .B1(DP_mult_206_n2253), .B2(DP_mult_206_n1562), .ZN(DP_mult_206_n1271)
         );
  OAI22_X1 DP_mult_206_U2576 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1755), 
        .B1(DP_mult_206_n1754), .B2(DP_mult_206_n2265), .ZN(DP_mult_206_n1456)
         );
  OAI22_X1 DP_mult_206_U2575 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1751), 
        .B1(DP_mult_206_n1750), .B2(DP_mult_206_n2266), .ZN(DP_mult_206_n1452)
         );
  OAI22_X1 DP_mult_206_U2574 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1752), 
        .B1(DP_mult_206_n2266), .B2(DP_mult_206_n1751), .ZN(DP_mult_206_n1453)
         );
  OAI22_X1 DP_mult_206_U2573 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1754), 
        .B1(DP_mult_206_n2265), .B2(DP_mult_206_n1753), .ZN(DP_mult_206_n1455)
         );
  OAI22_X1 DP_mult_206_U2572 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1746), 
        .B1(DP_mult_206_n2265), .B2(DP_mult_206_n1745), .ZN(DP_mult_206_n1447)
         );
  OAI22_X1 DP_mult_206_U2571 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1744), 
        .B1(DP_mult_206_n2266), .B2(DP_mult_206_n1743), .ZN(DP_mult_206_n1445)
         );
  OAI22_X1 DP_mult_206_U2570 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1748), 
        .B1(DP_mult_206_n2265), .B2(DP_mult_206_n1747), .ZN(DP_mult_206_n1449)
         );
  OAI22_X1 DP_mult_206_U2569 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1745), 
        .B1(DP_mult_206_n1744), .B2(DP_mult_206_n2266), .ZN(DP_mult_206_n1446)
         );
  OAI22_X1 DP_mult_206_U2568 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1749), 
        .B1(DP_mult_206_n1748), .B2(DP_mult_206_n2265), .ZN(DP_mult_206_n1450)
         );
  OAI22_X1 DP_mult_206_U2567 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1750), 
        .B1(DP_mult_206_n2266), .B2(DP_mult_206_n1749), .ZN(DP_mult_206_n1451)
         );
  OAI22_X1 DP_mult_206_U2566 ( .A1(DP_mult_206_n2031), .A2(DP_mult_206_n1747), 
        .B1(DP_mult_206_n1746), .B2(DP_mult_206_n2266), .ZN(DP_mult_206_n1448)
         );
  OAI22_X1 DP_mult_206_U2565 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1753), 
        .B1(DP_mult_206_n1752), .B2(DP_mult_206_n2266), .ZN(DP_mult_206_n1454)
         );
  OAI21_X1 DP_mult_206_U2564 ( .B1(DP_mult_206_n594), .B2(DP_mult_206_n582), 
        .A(DP_mult_206_n583), .ZN(DP_mult_206_n581) );
  XNOR2_X1 DP_mult_206_U2563 ( .A(DP_mult_206_n379), .B(DP_mult_206_n305), 
        .ZN(DP_pipe0_coeff_pipe00[19]) );
  INV_X1 DP_mult_206_U2562 ( .A(DP_mult_206_n2109), .ZN(DP_mult_206_n671) );
  XNOR2_X1 DP_mult_206_U2561 ( .A(DP_mult_206_n353), .B(DP_mult_206_n303), 
        .ZN(DP_pipe0_coeff_pipe00[21]) );
  OAI22_X1 DP_mult_206_U2560 ( .A1(DP_mult_206_n2033), .A2(DP_mult_206_n1553), 
        .B1(DP_mult_206_n1552), .B2(DP_mult_206_n2250), .ZN(DP_mult_206_n1262)
         );
  OAI22_X1 DP_mult_206_U2559 ( .A1(DP_mult_206_n2129), .A2(DP_mult_206_n1554), 
        .B1(DP_mult_206_n2249), .B2(DP_mult_206_n1553), .ZN(DP_mult_206_n1263)
         );
  OAI22_X1 DP_mult_206_U2558 ( .A1(DP_mult_206_n2130), .A2(DP_mult_206_n1545), 
        .B1(DP_mult_206_n1544), .B2(DP_mult_206_n2250), .ZN(DP_mult_206_n1254)
         );
  OAI22_X1 DP_mult_206_U2557 ( .A1(DP_mult_206_n2033), .A2(DP_mult_206_n1547), 
        .B1(DP_mult_206_n1546), .B2(DP_mult_206_n2249), .ZN(DP_mult_206_n1256)
         );
  OAI22_X1 DP_mult_206_U2556 ( .A1(DP_mult_206_n2223), .A2(DP_mult_206_n1548), 
        .B1(DP_mult_206_n2249), .B2(DP_mult_206_n1547), .ZN(DP_mult_206_n1257)
         );
  OAI22_X1 DP_mult_206_U2555 ( .A1(DP_mult_206_n1944), .A2(DP_mult_206_n1549), 
        .B1(DP_mult_206_n1548), .B2(DP_mult_206_n2249), .ZN(DP_mult_206_n1258)
         );
  OAI22_X1 DP_mult_206_U2554 ( .A1(DP_mult_206_n2224), .A2(DP_mult_206_n1546), 
        .B1(DP_mult_206_n2250), .B2(DP_mult_206_n1545), .ZN(DP_mult_206_n1255)
         );
  OAI22_X1 DP_mult_206_U2553 ( .A1(DP_mult_206_n1550), .A2(DP_mult_206_n2033), 
        .B1(DP_mult_206_n2249), .B2(DP_mult_206_n1549), .ZN(DP_mult_206_n1259)
         );
  OAI22_X1 DP_mult_206_U2552 ( .A1(DP_mult_206_n2130), .A2(DP_mult_206_n1555), 
        .B1(DP_mult_206_n1554), .B2(DP_mult_206_n2249), .ZN(DP_mult_206_n1264)
         );
  OAI22_X1 DP_mult_206_U2551 ( .A1(DP_mult_206_n2224), .A2(DP_mult_206_n1552), 
        .B1(DP_mult_206_n2249), .B2(DP_mult_206_n1551), .ZN(DP_mult_206_n1261)
         );
  OAI22_X1 DP_mult_206_U2550 ( .A1(DP_mult_206_n1944), .A2(DP_mult_206_n1544), 
        .B1(DP_mult_206_n2250), .B2(DP_mult_206_n1543), .ZN(DP_mult_206_n1253)
         );
  XNOR2_X1 DP_mult_206_U2549 ( .A(DP_mult_206_n342), .B(DP_mult_206_n302), 
        .ZN(DP_pipe0_coeff_pipe00[22]) );
  INV_X1 DP_mult_206_U2548 ( .A(DP_mult_206_n1952), .ZN(DP_mult_206_n917) );
  XNOR2_X1 DP_mult_206_U2547 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2321), .ZN(
        DP_mult_206_n1515) );
  XNOR2_X1 DP_mult_206_U2546 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2321), .ZN(
        DP_mult_206_n1511) );
  XNOR2_X1 DP_mult_206_U2545 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2321), .ZN(
        DP_mult_206_n1517) );
  XNOR2_X1 DP_mult_206_U2544 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2320), .ZN(
        DP_mult_206_n1509) );
  XNOR2_X1 DP_mult_206_U2543 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2321), .ZN(
        DP_mult_206_n1519) );
  XNOR2_X1 DP_mult_206_U2542 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2320), .ZN(
        DP_mult_206_n1513) );
  INV_X1 DP_mult_206_U2541 ( .A(DP_mult_206_n401), .ZN(DP_mult_206_n399) );
  OAI22_X1 DP_mult_206_U2540 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1703), 
        .B1(DP_mult_206_n1702), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1406)
         );
  OAI22_X1 DP_mult_206_U2539 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1705), 
        .B1(DP_mult_206_n1704), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1408)
         );
  NAND2_X1 DP_mult_206_U2538 ( .A1(DP_mult_206_n761), .A2(DP_mult_206_n774), 
        .ZN(DP_mult_206_n461) );
  NAND2_X1 DP_mult_206_U2537 ( .A1(DP_mult_206_n919), .A2(DP_mult_206_n940), 
        .ZN(DP_mult_206_n543) );
  AOI21_X1 DP_mult_206_U2536 ( .B1(DP_mult_206_n589), .B2(DP_mult_206_n2175), 
        .A(DP_mult_206_n1974), .ZN(DP_mult_206_n583) );
  NAND2_X1 DP_mult_206_U2535 ( .A1(DP_mult_206_n588), .A2(DP_mult_206_n2175), 
        .ZN(DP_mult_206_n582) );
  OAI22_X1 DP_mult_206_U2534 ( .A1(DP_mult_206_n2130), .A2(DP_mult_206_n1539), 
        .B1(DP_mult_206_n1538), .B2(DP_mult_206_n2250), .ZN(DP_mult_206_n1248)
         );
  OAI22_X1 DP_mult_206_U2533 ( .A1(DP_mult_206_n2223), .A2(DP_mult_206_n1540), 
        .B1(DP_mult_206_n2250), .B2(DP_mult_206_n1539), .ZN(DP_mult_206_n1249)
         );
  OAI22_X1 DP_mult_206_U2532 ( .A1(DP_mult_206_n2129), .A2(DP_mult_206_n1533), 
        .B1(DP_mult_206_n1532), .B2(DP_mult_206_n2250), .ZN(DP_mult_206_n692)
         );
  OAI22_X1 DP_mult_206_U2531 ( .A1(DP_mult_206_n2129), .A2(DP_mult_206_n1541), 
        .B1(DP_mult_206_n1540), .B2(DP_mult_206_n2250), .ZN(DP_mult_206_n1250)
         );
  OAI22_X1 DP_mult_206_U2530 ( .A1(DP_mult_206_n2224), .A2(DP_mult_206_n1538), 
        .B1(DP_mult_206_n2249), .B2(DP_mult_206_n1537), .ZN(DP_mult_206_n1247)
         );
  OAI22_X1 DP_mult_206_U2529 ( .A1(DP_mult_206_n2130), .A2(DP_mult_206_n1542), 
        .B1(DP_mult_206_n2249), .B2(DP_mult_206_n1541), .ZN(DP_mult_206_n1251)
         );
  OAI22_X1 DP_mult_206_U2528 ( .A1(DP_mult_206_n2224), .A2(DP_mult_206_n1543), 
        .B1(DP_mult_206_n1542), .B2(DP_mult_206_n2250), .ZN(DP_mult_206_n1252)
         );
  OAI22_X1 DP_mult_206_U2527 ( .A1(DP_mult_206_n2129), .A2(DP_mult_206_n2318), 
        .B1(DP_mult_206_n1556), .B2(DP_mult_206_n2249), .ZN(DP_mult_206_n1184)
         );
  OAI22_X1 DP_mult_206_U2526 ( .A1(DP_mult_206_n2130), .A2(DP_mult_206_n1534), 
        .B1(DP_mult_206_n2249), .B2(DP_mult_206_n1533), .ZN(DP_mult_206_n1243)
         );
  OAI22_X1 DP_mult_206_U2525 ( .A1(DP_mult_206_n1944), .A2(DP_mult_206_n1537), 
        .B1(DP_mult_206_n1536), .B2(DP_mult_206_n2250), .ZN(DP_mult_206_n1246)
         );
  OAI22_X1 DP_mult_206_U2524 ( .A1(DP_mult_206_n2224), .A2(DP_mult_206_n1535), 
        .B1(DP_mult_206_n1534), .B2(DP_mult_206_n2250), .ZN(DP_mult_206_n1244)
         );
  OAI22_X1 DP_mult_206_U2523 ( .A1(DP_mult_206_n2129), .A2(DP_mult_206_n1536), 
        .B1(DP_mult_206_n2250), .B2(DP_mult_206_n1535), .ZN(DP_mult_206_n1245)
         );
  OAI22_X1 DP_mult_206_U2522 ( .A1(DP_mult_206_n1988), .A2(DP_mult_206_n2310), 
        .B1(DP_mult_206_n1606), .B2(DP_mult_206_n2255), .ZN(DP_mult_206_n1186)
         );
  OAI22_X1 DP_mult_206_U2521 ( .A1(DP_mult_206_n1988), .A2(DP_mult_206_n1585), 
        .B1(DP_mult_206_n1584), .B2(DP_mult_206_n2256), .ZN(DP_mult_206_n1292)
         );
  OAI22_X1 DP_mult_206_U2520 ( .A1(DP_mult_206_n2228), .A2(DP_mult_206_n1586), 
        .B1(DP_mult_206_n2256), .B2(DP_mult_206_n1585), .ZN(DP_mult_206_n1293)
         );
  OAI22_X1 DP_mult_206_U2519 ( .A1(DP_mult_206_n2228), .A2(DP_mult_206_n1592), 
        .B1(DP_mult_206_n2256), .B2(DP_mult_206_n1591), .ZN(DP_mult_206_n1299)
         );
  OAI22_X1 DP_mult_206_U2518 ( .A1(DP_mult_206_n2227), .A2(DP_mult_206_n1591), 
        .B1(DP_mult_206_n1590), .B2(DP_mult_206_n2256), .ZN(DP_mult_206_n1298)
         );
  OAI22_X1 DP_mult_206_U2517 ( .A1(DP_mult_206_n1988), .A2(DP_mult_206_n1587), 
        .B1(DP_mult_206_n1586), .B2(DP_mult_206_n2256), .ZN(DP_mult_206_n1294)
         );
  OAI22_X1 DP_mult_206_U2516 ( .A1(DP_mult_206_n2024), .A2(DP_mult_206_n1583), 
        .B1(DP_mult_206_n1582), .B2(DP_mult_206_n2256), .ZN(DP_mult_206_n724)
         );
  OAI22_X1 DP_mult_206_U2515 ( .A1(DP_mult_206_n1988), .A2(DP_mult_206_n1588), 
        .B1(DP_mult_206_n2255), .B2(DP_mult_206_n1587), .ZN(DP_mult_206_n1295)
         );
  OAI22_X1 DP_mult_206_U2514 ( .A1(DP_mult_206_n2228), .A2(DP_mult_206_n1589), 
        .B1(DP_mult_206_n1588), .B2(DP_mult_206_n2255), .ZN(DP_mult_206_n1296)
         );
  OAI22_X1 DP_mult_206_U2513 ( .A1(DP_mult_206_n2228), .A2(DP_mult_206_n1590), 
        .B1(DP_mult_206_n2255), .B2(DP_mult_206_n1589), .ZN(DP_mult_206_n1297)
         );
  OAI22_X1 DP_mult_206_U2512 ( .A1(DP_mult_206_n2228), .A2(DP_mult_206_n1584), 
        .B1(DP_mult_206_n2256), .B2(DP_mult_206_n1583), .ZN(DP_mult_206_n1291)
         );
  OAI22_X1 DP_mult_206_U2511 ( .A1(DP_mult_206_n1987), .A2(DP_mult_206_n1593), 
        .B1(DP_mult_206_n1592), .B2(DP_mult_206_n2255), .ZN(DP_mult_206_n1300)
         );
  OAI21_X1 DP_mult_206_U2510 ( .B1(DP_mult_206_n2144), .B2(DP_mult_206_n521), 
        .A(DP_mult_206_n514), .ZN(DP_mult_206_n512) );
  OAI22_X1 DP_mult_206_U2509 ( .A1(DP_mult_206_n2234), .A2(DP_mult_206_n1674), 
        .B1(DP_mult_206_n1673), .B2(DP_mult_206_n2260), .ZN(DP_mult_206_n1378)
         );
  OAI22_X1 DP_mult_206_U2508 ( .A1(DP_mult_206_n2233), .A2(DP_mult_206_n1680), 
        .B1(DP_mult_206_n1679), .B2(DP_mult_206_n2201), .ZN(DP_mult_206_n1384)
         );
  OAI22_X1 DP_mult_206_U2507 ( .A1(DP_mult_206_n1941), .A2(DP_mult_206_n1678), 
        .B1(DP_mult_206_n1677), .B2(DP_mult_206_n2201), .ZN(DP_mult_206_n1382)
         );
  OAI22_X1 DP_mult_206_U2506 ( .A1(DP_mult_206_n2233), .A2(DP_mult_206_n1676), 
        .B1(DP_mult_206_n1675), .B2(DP_mult_206_n2260), .ZN(DP_mult_206_n1380)
         );
  OAI22_X1 DP_mult_206_U2505 ( .A1(DP_mult_206_n1942), .A2(DP_mult_206_n1679), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1678), .ZN(DP_mult_206_n1383)
         );
  OAI22_X1 DP_mult_206_U2504 ( .A1(DP_mult_206_n1942), .A2(DP_mult_206_n1673), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1672), .ZN(DP_mult_206_n1377)
         );
  OAI22_X1 DP_mult_206_U2503 ( .A1(DP_mult_206_n1942), .A2(DP_mult_206_n1677), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1676), .ZN(DP_mult_206_n1381)
         );
  OAI22_X1 DP_mult_206_U2502 ( .A1(DP_mult_206_n2233), .A2(DP_mult_206_n1671), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1670), .ZN(DP_mult_206_n1375)
         );
  OAI22_X1 DP_mult_206_U2501 ( .A1(DP_mult_206_n2233), .A2(DP_mult_206_n1672), 
        .B1(DP_mult_206_n1671), .B2(DP_mult_206_n2260), .ZN(DP_mult_206_n1376)
         );
  OAI22_X1 DP_mult_206_U2500 ( .A1(DP_mult_206_n1942), .A2(DP_mult_206_n1670), 
        .B1(DP_mult_206_n1669), .B2(DP_mult_206_n2260), .ZN(DP_mult_206_n1374)
         );
  OAI22_X1 DP_mult_206_U2499 ( .A1(DP_mult_206_n2233), .A2(DP_mult_206_n1669), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1668), .ZN(DP_mult_206_n1373)
         );
  OAI22_X1 DP_mult_206_U2498 ( .A1(DP_mult_206_n1941), .A2(DP_mult_206_n1675), 
        .B1(DP_mult_206_n2260), .B2(DP_mult_206_n1674), .ZN(DP_mult_206_n1379)
         );
  XNOR2_X1 DP_mult_206_U2497 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1594) );
  XNOR2_X1 DP_mult_206_U2496 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1586) );
  XNOR2_X1 DP_mult_206_U2495 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1584) );
  XNOR2_X1 DP_mult_206_U2494 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1590) );
  XNOR2_X1 DP_mult_206_U2493 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1592) );
  XNOR2_X1 DP_mult_206_U2492 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1588) );
  INV_X1 DP_mult_206_U2491 ( .A(DP_mult_206_n706), .ZN(DP_mult_206_n707) );
  AOI21_X1 DP_mult_206_U2490 ( .B1(DP_mult_206_n346), .B2(DP_mult_206_n2185), 
        .A(DP_mult_206_n339), .ZN(DP_mult_206_n337) );
  AOI21_X1 DP_mult_206_U2489 ( .B1(DP_mult_206_n383), .B2(DP_mult_206_n2182), 
        .A(DP_mult_206_n376), .ZN(DP_mult_206_n372) );
  AOI21_X1 DP_mult_206_U2488 ( .B1(DP_mult_206_n423), .B2(DP_mult_206_n356), 
        .A(DP_mult_206_n359), .ZN(DP_mult_206_n355) );
  NAND2_X1 DP_mult_206_U2487 ( .A1(DP_mult_206_n382), .A2(DP_mult_206_n2182), 
        .ZN(DP_mult_206_n371) );
  NAND2_X1 DP_mult_206_U2486 ( .A1(DP_mult_206_n422), .A2(DP_mult_206_n356), 
        .ZN(DP_mult_206_n354) );
  INV_X1 DP_mult_206_U2485 ( .A(DP_mult_206_n346), .ZN(DP_mult_206_n344) );
  NAND2_X1 DP_mult_206_U2484 ( .A1(DP_mult_206_n2182), .A2(DP_mult_206_n378), 
        .ZN(DP_mult_206_n305) );
  OAI22_X1 DP_mult_206_U2483 ( .A1(DP_mult_206_n2238), .A2(DP_mult_206_n1712), 
        .B1(DP_mult_206_n1711), .B2(DP_mult_206_n2263), .ZN(DP_mult_206_n1414)
         );
  OAI22_X1 DP_mult_206_U2482 ( .A1(DP_mult_206_n2238), .A2(DP_mult_206_n1710), 
        .B1(DP_mult_206_n1709), .B2(DP_mult_206_n2263), .ZN(DP_mult_206_n1412)
         );
  OAI22_X1 DP_mult_206_U2481 ( .A1(DP_mult_206_n2237), .A2(DP_mult_206_n1708), 
        .B1(DP_mult_206_n1707), .B2(DP_mult_206_n2264), .ZN(DP_mult_206_n874)
         );
  OAI22_X1 DP_mult_206_U2480 ( .A1(DP_mult_206_n2160), .A2(DP_mult_206_n1709), 
        .B1(DP_mult_206_n2263), .B2(DP_mult_206_n1708), .ZN(DP_mult_206_n1411)
         );
  OAI22_X1 DP_mult_206_U2479 ( .A1(DP_mult_206_n2160), .A2(DP_mult_206_n1717), 
        .B1(DP_mult_206_n2264), .B2(DP_mult_206_n1716), .ZN(DP_mult_206_n1419)
         );
  OAI22_X1 DP_mult_206_U2478 ( .A1(DP_mult_206_n2159), .A2(DP_mult_206_n1715), 
        .B1(DP_mult_206_n2264), .B2(DP_mult_206_n1714), .ZN(DP_mult_206_n1417)
         );
  OAI22_X1 DP_mult_206_U2477 ( .A1(DP_mult_206_n2237), .A2(DP_mult_206_n1716), 
        .B1(DP_mult_206_n1715), .B2(DP_mult_206_n2263), .ZN(DP_mult_206_n1418)
         );
  OAI22_X1 DP_mult_206_U2476 ( .A1(DP_mult_206_n2159), .A2(DP_mult_206_n1713), 
        .B1(DP_mult_206_n2263), .B2(DP_mult_206_n1712), .ZN(DP_mult_206_n1415)
         );
  OAI22_X1 DP_mult_206_U2475 ( .A1(DP_mult_206_n2160), .A2(DP_mult_206_n1711), 
        .B1(DP_mult_206_n2264), .B2(DP_mult_206_n1710), .ZN(DP_mult_206_n1413)
         );
  OAI22_X1 DP_mult_206_U2474 ( .A1(DP_mult_206_n2160), .A2(DP_mult_206_n1718), 
        .B1(DP_mult_206_n1717), .B2(DP_mult_206_n2263), .ZN(DP_mult_206_n1420)
         );
  OAI22_X1 DP_mult_206_U2473 ( .A1(DP_mult_206_n2237), .A2(DP_mult_206_n2285), 
        .B1(DP_mult_206_n1731), .B2(DP_mult_206_n2263), .ZN(DP_mult_206_n1191)
         );
  NAND2_X1 DP_mult_206_U2472 ( .A1(DP_mult_206_n839), .A2(DP_mult_206_n856), 
        .ZN(DP_mult_206_n514) );
  XNOR2_X1 DP_mult_206_U2471 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2294), .ZN(
        DP_mult_206_n1659) );
  XNOR2_X1 DP_mult_206_U2470 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2294), .ZN(
        DP_mult_206_n1667) );
  XNOR2_X1 DP_mult_206_U2469 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2293), .ZN(
        DP_mult_206_n1665) );
  XNOR2_X1 DP_mult_206_U2468 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2293), .ZN(
        DP_mult_206_n1661) );
  XNOR2_X1 DP_mult_206_U2467 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2294), .ZN(
        DP_mult_206_n1669) );
  OAI22_X1 DP_mult_206_U2466 ( .A1(DP_mult_206_n2231), .A2(DP_mult_206_n1651), 
        .B1(DP_mult_206_n1650), .B2(DP_mult_206_n2056), .ZN(DP_mult_206_n1356)
         );
  XNOR2_X1 DP_mult_206_U2465 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2293), .ZN(
        DP_mult_206_n1663) );
  OAI22_X1 DP_mult_206_U2464 ( .A1(DP_mult_206_n2231), .A2(DP_mult_206_n1646), 
        .B1(DP_mult_206_n2259), .B2(DP_mult_206_n1645), .ZN(DP_mult_206_n1351)
         );
  OAI22_X1 DP_mult_206_U2463 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1650), 
        .B1(DP_mult_206_n2056), .B2(DP_mult_206_n1649), .ZN(DP_mult_206_n1355)
         );
  OAI22_X1 DP_mult_206_U2462 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1654), 
        .B1(DP_mult_206_n2056), .B2(DP_mult_206_n1653), .ZN(DP_mult_206_n1359)
         );
  OAI22_X1 DP_mult_206_U2461 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1644), 
        .B1(DP_mult_206_n2259), .B2(DP_mult_206_n1643), .ZN(DP_mult_206_n1349)
         );
  OAI22_X1 DP_mult_206_U2460 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1648), 
        .B1(DP_mult_206_n2056), .B2(DP_mult_206_n1647), .ZN(DP_mult_206_n1353)
         );
  OAI22_X1 DP_mult_206_U2459 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1645), 
        .B1(DP_mult_206_n1644), .B2(DP_mult_206_n2056), .ZN(DP_mult_206_n1350)
         );
  OAI22_X1 DP_mult_206_U2458 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1649), 
        .B1(DP_mult_206_n1648), .B2(DP_mult_206_n2259), .ZN(DP_mult_206_n1354)
         );
  OAI22_X1 DP_mult_206_U2457 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1647), 
        .B1(DP_mult_206_n1646), .B2(DP_mult_206_n2056), .ZN(DP_mult_206_n1352)
         );
  OAI22_X1 DP_mult_206_U2456 ( .A1(DP_mult_206_n2035), .A2(DP_mult_206_n1652), 
        .B1(DP_mult_206_n2056), .B2(DP_mult_206_n1651), .ZN(DP_mult_206_n1357)
         );
  OAI21_X1 DP_mult_206_U2455 ( .B1(DP_mult_206_n2232), .B2(DP_mult_206_n2192), 
        .A(DP_mult_206_n2333), .ZN(DP_mult_206_n1338) );
  OAI22_X1 DP_mult_206_U2454 ( .A1(DP_mult_206_n2061), .A2(DP_mult_206_n1628), 
        .B1(DP_mult_206_n1627), .B2(DP_mult_206_n2258), .ZN(DP_mult_206_n1334)
         );
  OAI22_X1 DP_mult_206_U2453 ( .A1(DP_mult_206_n2229), .A2(DP_mult_206_n1624), 
        .B1(DP_mult_206_n1623), .B2(DP_mult_206_n2258), .ZN(DP_mult_206_n1330)
         );
  OAI22_X1 DP_mult_206_U2452 ( .A1(DP_mult_206_n2230), .A2(DP_mult_206_n1622), 
        .B1(DP_mult_206_n1621), .B2(DP_mult_206_n2257), .ZN(DP_mult_206_n1328)
         );
  OAI22_X1 DP_mult_206_U2451 ( .A1(DP_mult_206_n2060), .A2(DP_mult_206_n1627), 
        .B1(DP_mult_206_n2258), .B2(DP_mult_206_n1626), .ZN(DP_mult_206_n1333)
         );
  OAI22_X1 DP_mult_206_U2450 ( .A1(DP_mult_206_n2060), .A2(DP_mult_206_n1619), 
        .B1(DP_mult_206_n2257), .B2(DP_mult_206_n1618), .ZN(DP_mult_206_n1325)
         );
  OAI22_X1 DP_mult_206_U2449 ( .A1(DP_mult_206_n2061), .A2(DP_mult_206_n1621), 
        .B1(DP_mult_206_n2258), .B2(DP_mult_206_n1620), .ZN(DP_mult_206_n1327)
         );
  OAI22_X1 DP_mult_206_U2448 ( .A1(DP_mult_206_n2230), .A2(DP_mult_206_n1630), 
        .B1(DP_mult_206_n1629), .B2(DP_mult_206_n2257), .ZN(DP_mult_206_n1336)
         );
  OAI22_X1 DP_mult_206_U2447 ( .A1(DP_mult_206_n2060), .A2(DP_mult_206_n1623), 
        .B1(DP_mult_206_n2257), .B2(DP_mult_206_n1622), .ZN(DP_mult_206_n1329)
         );
  OAI22_X1 DP_mult_206_U2446 ( .A1(DP_mult_206_n2061), .A2(DP_mult_206_n1625), 
        .B1(DP_mult_206_n2258), .B2(DP_mult_206_n1624), .ZN(DP_mult_206_n1331)
         );
  OAI22_X1 DP_mult_206_U2445 ( .A1(DP_mult_206_n2230), .A2(DP_mult_206_n1626), 
        .B1(DP_mult_206_n1625), .B2(DP_mult_206_n2257), .ZN(DP_mult_206_n1332)
         );
  OAI22_X1 DP_mult_206_U2444 ( .A1(DP_mult_206_n2061), .A2(DP_mult_206_n1629), 
        .B1(DP_mult_206_n2258), .B2(DP_mult_206_n1628), .ZN(DP_mult_206_n1335)
         );
  OAI22_X1 DP_mult_206_U2443 ( .A1(DP_mult_206_n2230), .A2(DP_mult_206_n1620), 
        .B1(DP_mult_206_n1619), .B2(DP_mult_206_n2257), .ZN(DP_mult_206_n1326)
         );
  AOI21_X1 DP_mult_206_U2442 ( .B1(DP_mult_206_n490), .B2(DP_mult_206_n454), 
        .A(DP_mult_206_n455), .ZN(DP_mult_206_n453) );
  NAND2_X1 DP_mult_206_U2441 ( .A1(DP_mult_206_n489), .A2(DP_mult_206_n454), 
        .ZN(DP_mult_206_n452) );
  NAND2_X1 DP_mult_206_U2440 ( .A1(DP_mult_206_n805), .A2(DP_mult_206_n820), 
        .ZN(DP_mult_206_n496) );
  OAI21_X1 DP_mult_206_U2439 ( .B1(DP_mult_206_n492), .B2(DP_mult_206_n480), 
        .A(DP_mult_206_n481), .ZN(DP_mult_206_n479) );
  OAI21_X1 DP_mult_206_U2438 ( .B1(DP_mult_206_n492), .B2(DP_mult_206_n467), 
        .A(DP_mult_206_n468), .ZN(DP_mult_206_n466) );
  XNOR2_X1 DP_mult_206_U2437 ( .A(DP_mult_206_n475), .B(DP_mult_206_n314), 
        .ZN(DP_pipe0_coeff_pipe00[10]) );
  INV_X1 DP_mult_206_U2436 ( .A(DP_mult_206_n542), .ZN(DP_mult_206_n673) );
  NOR2_X1 DP_mult_206_U2435 ( .A1(DP_mult_206_n547), .A2(DP_mult_206_n542), 
        .ZN(DP_mult_206_n540) );
  OAI21_X1 DP_mult_206_U2434 ( .B1(DP_mult_206_n542), .B2(DP_mult_206_n550), 
        .A(DP_mult_206_n543), .ZN(DP_mult_206_n541) );
  INV_X1 DP_mult_206_U2433 ( .A(DP_mult_206_n474), .ZN(DP_mult_206_n472) );
  NAND2_X1 DP_mult_206_U2432 ( .A1(DP_mult_206_n1989), .A2(DP_mult_206_n474), 
        .ZN(DP_mult_206_n314) );
  NAND2_X1 DP_mult_206_U2431 ( .A1(DP_mult_206_n511), .A2(DP_mult_206_n525), 
        .ZN(DP_mult_206_n505) );
  NAND2_X1 DP_mult_206_U2430 ( .A1(DP_mult_206_n465), .A2(DP_mult_206_n507), 
        .ZN(DP_mult_206_n463) );
  NAND2_X1 DP_mult_206_U2429 ( .A1(DP_mult_206_n1963), .A2(DP_mult_206_n670), 
        .ZN(DP_mult_206_n516) );
  NAND2_X1 DP_mult_206_U2428 ( .A1(DP_mult_206_n507), .A2(DP_mult_206_n668), 
        .ZN(DP_mult_206_n498) );
  NAND2_X1 DP_mult_206_U2427 ( .A1(DP_mult_206_n507), .A2(DP_mult_206_n489), 
        .ZN(DP_mult_206_n487) );
  INV_X1 DP_mult_206_U2426 ( .A(DP_mult_206_n1963), .ZN(DP_mult_206_n523) );
  NAND2_X1 DP_mult_206_U2425 ( .A1(DP_mult_206_n478), .A2(DP_mult_206_n507), 
        .ZN(DP_mult_206_n476) );
  AOI21_X1 DP_mult_206_U2424 ( .B1(DP_mult_206_n2153), .B2(DP_mult_206_n2002), 
        .A(DP_mult_206_n451), .ZN(DP_mult_206_n301) );
  AOI21_X1 DP_mult_206_U2423 ( .B1(DP_mult_206_n537), .B2(DP_mult_206_n450), 
        .A(DP_mult_206_n451), .ZN(DP_mult_206_n2218) );
  AOI21_X1 DP_mult_206_U2422 ( .B1(DP_mult_206_n2153), .B2(DP_mult_206_n450), 
        .A(DP_mult_206_n451), .ZN(DP_mult_206_n2219) );
  NAND2_X1 DP_mult_206_U2421 ( .A1(DP_mult_206_n1171), .A2(DP_mult_206_n1174), 
        .ZN(DP_mult_206_n634) );
  NOR2_X1 DP_mult_206_U2420 ( .A1(DP_mult_206_n1171), .A2(DP_mult_206_n1174), 
        .ZN(DP_mult_206_n633) );
  INV_X1 DP_mult_206_U2419 ( .A(DP_mult_206_n382), .ZN(DP_mult_206_n380) );
  NOR2_X1 DP_mult_206_U2418 ( .A1(DP_mult_206_n897), .A2(DP_mult_206_n918), 
        .ZN(DP_mult_206_n534) );
  INV_X1 DP_mult_206_U2417 ( .A(DP_mult_206_n2203), .ZN(DP_mult_206_n508) );
  AOI21_X1 DP_mult_206_U2416 ( .B1(DP_mult_206_n2204), .B2(DP_mult_206_n670), 
        .A(DP_mult_206_n519), .ZN(DP_mult_206_n517) );
  INV_X1 DP_mult_206_U2415 ( .A(DP_mult_206_n2204), .ZN(DP_mult_206_n524) );
  NAND2_X1 DP_mult_206_U2414 ( .A1(DP_mult_206_n709), .A2(DP_mult_206_n716), 
        .ZN(DP_mult_206_n409) );
  AOI21_X1 DP_mult_206_U2413 ( .B1(DP_mult_206_n508), .B2(DP_mult_206_n465), 
        .A(DP_mult_206_n466), .ZN(DP_mult_206_n464) );
  AOI21_X1 DP_mult_206_U2412 ( .B1(DP_mult_206_n508), .B2(DP_mult_206_n668), 
        .A(DP_mult_206_n501), .ZN(DP_mult_206_n499) );
  AOI21_X1 DP_mult_206_U2411 ( .B1(DP_mult_206_n508), .B2(DP_mult_206_n478), 
        .A(DP_mult_206_n479), .ZN(DP_mult_206_n477) );
  XNOR2_X1 DP_mult_206_U2410 ( .A(DP_mult_206_n462), .B(DP_mult_206_n313), 
        .ZN(DP_pipe0_coeff_pipe00[11]) );
  NAND2_X1 DP_mult_206_U2409 ( .A1(DP_mult_206_n727), .A2(DP_mult_206_n736), 
        .ZN(DP_mult_206_n429) );
  NOR2_X1 DP_mult_206_U2408 ( .A1(DP_mult_206_n749), .A2(DP_mult_206_n760), 
        .ZN(DP_mult_206_n438) );
  NAND2_X1 DP_mult_206_U2407 ( .A1(DP_mult_206_n749), .A2(DP_mult_206_n760), 
        .ZN(DP_mult_206_n439) );
  OAI21_X1 DP_mult_206_U2406 ( .B1(DP_mult_206_n2137), .B2(DP_mult_206_n2019), 
        .A(DP_mult_206_n2339), .ZN(DP_mult_206_n1194) );
  XNOR2_X1 DP_mult_206_U2405 ( .A(DP_mult_206_n533), .B(DP_mult_206_n320), 
        .ZN(DP_pipe0_coeff_pipe00[4]) );
  NOR2_X1 DP_mult_206_U2404 ( .A1(DP_mult_206_n737), .A2(DP_mult_206_n748), 
        .ZN(DP_mult_206_n435) );
  OAI21_X1 DP_mult_206_U2403 ( .B1(DP_mult_206_n2158), .B2(DP_mult_206_n503), 
        .A(DP_mult_206_n496), .ZN(DP_mult_206_n490) );
  NOR2_X1 DP_mult_206_U2402 ( .A1(DP_mult_206_n805), .A2(DP_mult_206_n820), 
        .ZN(DP_mult_206_n495) );
  NAND2_X1 DP_mult_206_U2401 ( .A1(DP_mult_206_n1989), .A2(DP_mult_206_n2173), 
        .ZN(DP_mult_206_n456) );
  XNOR2_X1 DP_mult_206_U2400 ( .A(DP_mult_206_n504), .B(DP_mult_206_n317), 
        .ZN(DP_pipe0_coeff_pipe00[7]) );
  OAI21_X1 DP_mult_206_U2399 ( .B1(DP_mult_206_n2194), .B2(DP_mult_206_n1982), 
        .A(DP_mult_206_n2330), .ZN(DP_mult_206_n1410) );
  XNOR2_X1 DP_mult_206_U2398 ( .A(DP_mult_206_n522), .B(DP_mult_206_n319), 
        .ZN(DP_pipe0_coeff_pipe00[5]) );
  OAI22_X1 DP_mult_206_U2397 ( .A1(DP_mult_206_n1950), .A2(DP_mult_206_n1774), 
        .B1(DP_mult_206_n1773), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1475)
         );
  OAI22_X1 DP_mult_206_U2396 ( .A1(DP_mult_206_n2241), .A2(DP_mult_206_n1770), 
        .B1(DP_mult_206_n1769), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1471)
         );
  OAI22_X1 DP_mult_206_U2395 ( .A1(DP_mult_206_n2242), .A2(DP_mult_206_n1775), 
        .B1(DP_mult_206_n1774), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1476)
         );
  OAI22_X1 DP_mult_206_U2394 ( .A1(DP_mult_206_n2241), .A2(DP_mult_206_n1778), 
        .B1(DP_mult_206_n1777), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1479)
         );
  OAI22_X1 DP_mult_206_U2393 ( .A1(DP_mult_206_n2242), .A2(DP_mult_206_n1769), 
        .B1(DP_mult_206_n1768), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1470)
         );
  OAI22_X1 DP_mult_206_U2392 ( .A1(DP_mult_206_n2241), .A2(DP_mult_206_n1779), 
        .B1(DP_mult_206_n1778), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1480)
         );
  OAI22_X1 DP_mult_206_U2391 ( .A1(DP_mult_206_n2241), .A2(DP_mult_206_n1771), 
        .B1(DP_mult_206_n1770), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1472)
         );
  OAI22_X1 DP_mult_206_U2390 ( .A1(DP_mult_206_n1950), .A2(DP_mult_206_n1776), 
        .B1(DP_mult_206_n1775), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1477)
         );
  OAI22_X1 DP_mult_206_U2389 ( .A1(DP_mult_206_n1950), .A2(DP_mult_206_n1780), 
        .B1(DP_mult_206_n1779), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1481)
         );
  OAI22_X1 DP_mult_206_U2388 ( .A1(DP_mult_206_n1951), .A2(DP_mult_206_n1777), 
        .B1(DP_mult_206_n1776), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1478)
         );
  OAI22_X1 DP_mult_206_U2387 ( .A1(DP_mult_206_n1951), .A2(DP_mult_206_n1773), 
        .B1(DP_mult_206_n1772), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1474)
         );
  OAI22_X1 DP_mult_206_U2386 ( .A1(DP_mult_206_n2242), .A2(DP_mult_206_n1772), 
        .B1(DP_mult_206_n1771), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1473)
         );
  NAND2_X1 DP_mult_206_U2385 ( .A1(DP_mult_206_n1165), .A2(DP_mult_206_n1170), 
        .ZN(DP_mult_206_n632) );
  XNOR2_X1 DP_mult_206_U2384 ( .A(DP_mult_206_n515), .B(DP_mult_206_n318), 
        .ZN(DP_pipe0_coeff_pipe00[6]) );
  XNOR2_X1 DP_mult_206_U2383 ( .A(DP_mult_206_n497), .B(DP_mult_206_n316), 
        .ZN(DP_pipe0_coeff_pipe00[8]) );
  NOR2_X2 DP_mult_206_U2382 ( .A1(DP_mult_206_n789), .A2(DP_mult_206_n804), 
        .ZN(DP_mult_206_n480) );
  XNOR2_X1 DP_mult_206_U2381 ( .A(DP_mult_206_n486), .B(DP_mult_206_n315), 
        .ZN(DP_pipe0_coeff_pipe00[9]) );
  OAI21_X1 DP_mult_206_U2380 ( .B1(DP_mult_206_n2006), .B2(DP_mult_206_n2191), 
        .A(DP_mult_206_n2331), .ZN(DP_mult_206_n1386) );
  AOI21_X1 DP_mult_206_U2379 ( .B1(DP_mult_206_n1989), .B2(DP_mult_206_n483), 
        .A(DP_mult_206_n472), .ZN(DP_mult_206_n468) );
  INV_X1 DP_mult_206_U2378 ( .A(DP_mult_206_n418), .ZN(DP_mult_206_n416) );
  OAI21_X1 DP_mult_206_U2377 ( .B1(DP_mult_206_n337), .B2(DP_mult_206_n334), 
        .A(DP_mult_206_n335), .ZN(DP_mult_206_n333) );
  NAND2_X1 DP_mult_206_U2376 ( .A1(DP_mult_206_n2177), .A2(DP_mult_206_n418), 
        .ZN(DP_mult_206_n309) );
  NAND2_X1 DP_mult_206_U2375 ( .A1(DP_mult_206_n2172), .A2(DP_mult_206_n2174), 
        .ZN(DP_mult_206_n571) );
  AOI21_X1 DP_mult_206_U2374 ( .B1(DP_mult_206_n2172), .B2(DP_mult_206_n1966), 
        .A(DP_mult_206_n1972), .ZN(DP_mult_206_n572) );
  NOR2_X1 DP_mult_206_U2373 ( .A1(DP_mult_206_n520), .A2(DP_mult_206_n513), 
        .ZN(DP_mult_206_n511) );
  INV_X1 DP_mult_206_U2372 ( .A(DP_mult_206_n480), .ZN(DP_mult_206_n666) );
  NOR2_X1 DP_mult_206_U2371 ( .A1(DP_mult_206_n456), .A2(DP_mult_206_n480), 
        .ZN(DP_mult_206_n454) );
  NOR2_X1 DP_mult_206_U2370 ( .A1(DP_mult_206_n491), .A2(DP_mult_206_n480), 
        .ZN(DP_mult_206_n478) );
  OAI21_X1 DP_mult_206_U2369 ( .B1(DP_mult_206_n428), .B2(DP_mult_206_n436), 
        .A(DP_mult_206_n429), .ZN(DP_mult_206_n427) );
  INV_X1 DP_mult_206_U2368 ( .A(DP_mult_206_n428), .ZN(DP_mult_206_n661) );
  AOI21_X1 DP_mult_206_U2367 ( .B1(DP_mult_206_n423), .B2(DP_mult_206_n2177), 
        .A(DP_mult_206_n416), .ZN(DP_mult_206_n412) );
  NAND2_X1 DP_mult_206_U2366 ( .A1(DP_mult_206_n422), .A2(DP_mult_206_n2177), 
        .ZN(DP_mult_206_n411) );
  NAND2_X1 DP_mult_206_U2365 ( .A1(DP_mult_206_n332), .A2(DP_mult_206_n2186), 
        .ZN(DP_mult_206_n326) );
  NOR2_X1 DP_mult_206_U2364 ( .A1(DP_mult_206_n821), .A2(DP_mult_206_n838), 
        .ZN(DP_mult_206_n502) );
  OAI21_X1 DP_mult_206_U2363 ( .B1(DP_mult_206_n531), .B2(DP_mult_206_n535), 
        .A(DP_mult_206_n532), .ZN(DP_mult_206_n526) );
  NAND2_X1 DP_mult_206_U2362 ( .A1(DP_mult_206_n897), .A2(DP_mult_206_n918), 
        .ZN(DP_mult_206_n535) );
  OAI22_X1 DP_mult_206_U2361 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1699), 
        .B1(DP_mult_206_n1698), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1402)
         );
  OAI22_X1 DP_mult_206_U2360 ( .A1(DP_mult_206_n2135), .A2(DP_mult_206_n1700), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1699), .ZN(DP_mult_206_n1403)
         );
  OAI22_X1 DP_mult_206_U2359 ( .A1(DP_mult_206_n2134), .A2(DP_mult_206_n1697), 
        .B1(DP_mult_206_n1696), .B2(DP_mult_206_n2261), .ZN(DP_mult_206_n1400)
         );
  OAI22_X1 DP_mult_206_U2358 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1702), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1701), .ZN(DP_mult_206_n1405)
         );
  OAI22_X1 DP_mult_206_U2357 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1698), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1697), .ZN(DP_mult_206_n1401)
         );
  OAI22_X1 DP_mult_206_U2356 ( .A1(DP_mult_206_n2135), .A2(DP_mult_206_n1701), 
        .B1(DP_mult_206_n1700), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1404)
         );
  OAI22_X1 DP_mult_206_U2355 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1696), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1695), .ZN(DP_mult_206_n1399)
         );
  OAI22_X1 DP_mult_206_U2354 ( .A1(DP_mult_206_n2135), .A2(DP_mult_206_n1704), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1703), .ZN(DP_mult_206_n1407)
         );
  OAI22_X1 DP_mult_206_U2353 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1694), 
        .B1(DP_mult_206_n2039), .B2(DP_mult_206_n1693), .ZN(DP_mult_206_n1397)
         );
  OAI22_X1 DP_mult_206_U2352 ( .A1(DP_mult_206_n2235), .A2(DP_mult_206_n1695), 
        .B1(DP_mult_206_n1694), .B2(DP_mult_206_n2039), .ZN(DP_mult_206_n1398)
         );
  OAI21_X1 DP_mult_206_U2351 ( .B1(DP_mult_206_n456), .B2(DP_mult_206_n481), 
        .A(DP_mult_206_n457), .ZN(DP_mult_206_n455) );
  INV_X1 DP_mult_206_U2350 ( .A(DP_mult_206_n2158), .ZN(DP_mult_206_n667) );
  INV_X1 DP_mult_206_U2349 ( .A(DP_mult_206_n253), .ZN(DP_mult_206_n2268) );
  INV_X1 DP_mult_206_U2348 ( .A(DP_mult_206_n489), .ZN(DP_mult_206_n491) );
  INV_X1 DP_mult_206_U2347 ( .A(DP_mult_206_n502), .ZN(DP_mult_206_n668) );
  NAND2_X1 DP_mult_206_U2346 ( .A1(DP_mult_206_n1071), .A2(DP_mult_206_n1084), 
        .ZN(DP_mult_206_n591) );
  NOR2_X1 DP_mult_206_U2345 ( .A1(DP_mult_206_n633), .A2(DP_mult_206_n631), 
        .ZN(DP_mult_206_n629) );
  OAI21_X1 DP_mult_206_U2344 ( .B1(DP_mult_206_n631), .B2(DP_mult_206_n634), 
        .A(DP_mult_206_n632), .ZN(DP_mult_206_n630) );
  NOR2_X1 DP_mult_206_U2343 ( .A1(DP_mult_206_n1165), .A2(DP_mult_206_n1170), 
        .ZN(DP_mult_206_n631) );
  NAND2_X1 DP_mult_206_U2342 ( .A1(DP_mult_206_n941), .A2(DP_mult_206_n962), 
        .ZN(DP_mult_206_n550) );
  NAND3_X1 DP_mult_206_U2341 ( .A1(DP_mult_206_n2215), .A2(DP_mult_206_n2216), 
        .A3(DP_mult_206_n2217), .ZN(DP_mult_206_n822) );
  NAND2_X1 DP_mult_206_U2340 ( .A1(DP_mult_206_n827), .A2(DP_mult_206_n844), 
        .ZN(DP_mult_206_n2217) );
  NAND2_X1 DP_mult_206_U2339 ( .A1(DP_mult_206_n842), .A2(DP_mult_206_n844), 
        .ZN(DP_mult_206_n2216) );
  NAND2_X1 DP_mult_206_U2338 ( .A1(DP_mult_206_n2052), .A2(DP_mult_206_n827), 
        .ZN(DP_mult_206_n2215) );
  OAI21_X1 DP_mult_206_U2337 ( .B1(DP_mult_206_n1931), .B2(DP_mult_206_n2268), 
        .A(DP_mult_206_n2329), .ZN(DP_mult_206_n1434) );
  OAI21_X1 DP_mult_206_U2336 ( .B1(DP_mult_206_n566), .B2(DP_mult_206_n538), 
        .A(DP_mult_206_n539), .ZN(DP_mult_206_n537) );
  XNOR2_X1 DP_mult_206_U2335 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1775) );
  XNOR2_X1 DP_mult_206_U2334 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1773) );
  XNOR2_X1 DP_mult_206_U2333 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1779) );
  XNOR2_X1 DP_mult_206_U2332 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1777) );
  AOI21_X1 DP_mult_206_U2331 ( .B1(DP_mult_206_n595), .B2(DP_mult_206_n609), 
        .A(DP_mult_206_n596), .ZN(DP_mult_206_n594) );
  OAI22_X1 DP_mult_206_U2330 ( .A1(DP_mult_206_n2225), .A2(DP_mult_206_n1576), 
        .B1(DP_mult_206_n1575), .B2(DP_mult_206_n2253), .ZN(DP_mult_206_n1284)
         );
  OAI22_X1 DP_mult_206_U2329 ( .A1(DP_mult_206_n2225), .A2(DP_mult_206_n1574), 
        .B1(DP_mult_206_n1573), .B2(DP_mult_206_n2252), .ZN(DP_mult_206_n1282)
         );
  OAI22_X1 DP_mult_206_U2328 ( .A1(DP_mult_206_n2226), .A2(DP_mult_206_n1579), 
        .B1(DP_mult_206_n2252), .B2(DP_mult_206_n1578), .ZN(DP_mult_206_n1287)
         );
  OAI22_X1 DP_mult_206_U2327 ( .A1(DP_mult_206_n2225), .A2(DP_mult_206_n1572), 
        .B1(DP_mult_206_n1571), .B2(DP_mult_206_n2253), .ZN(DP_mult_206_n1280)
         );
  OAI22_X1 DP_mult_206_U2326 ( .A1(DP_mult_206_n2169), .A2(DP_mult_206_n1577), 
        .B1(DP_mult_206_n2252), .B2(DP_mult_206_n1576), .ZN(DP_mult_206_n1285)
         );
  OAI22_X1 DP_mult_206_U2325 ( .A1(DP_mult_206_n2226), .A2(DP_mult_206_n1573), 
        .B1(DP_mult_206_n2252), .B2(DP_mult_206_n1572), .ZN(DP_mult_206_n1281)
         );
  OAI22_X1 DP_mult_206_U2324 ( .A1(DP_mult_206_n2225), .A2(DP_mult_206_n1569), 
        .B1(DP_mult_206_n2252), .B2(DP_mult_206_n1568), .ZN(DP_mult_206_n1277)
         );
  OAI22_X1 DP_mult_206_U2323 ( .A1(DP_mult_206_n2226), .A2(DP_mult_206_n1575), 
        .B1(DP_mult_206_n2252), .B2(DP_mult_206_n1574), .ZN(DP_mult_206_n1283)
         );
  OAI22_X1 DP_mult_206_U2322 ( .A1(DP_mult_206_n2169), .A2(DP_mult_206_n1571), 
        .B1(DP_mult_206_n2252), .B2(DP_mult_206_n1570), .ZN(DP_mult_206_n1279)
         );
  OAI22_X1 DP_mult_206_U2321 ( .A1(DP_mult_206_n2169), .A2(DP_mult_206_n1570), 
        .B1(DP_mult_206_n1569), .B2(DP_mult_206_n2252), .ZN(DP_mult_206_n1278)
         );
  NOR2_X1 DP_mult_206_U2320 ( .A1(DP_mult_206_n571), .A2(DP_mult_206_n569), 
        .ZN(DP_mult_206_n567) );
  NAND2_X1 DP_mult_206_U2319 ( .A1(DP_mult_206_n1099), .A2(DP_mult_206_n1110), 
        .ZN(DP_mult_206_n598) );
  XNOR2_X1 DP_mult_206_U2318 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1550) );
  XNOR2_X1 DP_mult_206_U2317 ( .A(DP_mult_206_n2315), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1551) );
  AOI21_X1 DP_mult_206_U2316 ( .B1(DP_mult_206_n526), .B2(DP_mult_206_n511), 
        .A(DP_mult_206_n512), .ZN(DP_mult_206_n506) );
  NAND2_X1 DP_mult_206_U2315 ( .A1(DP_mult_206_n2213), .A2(DP_mult_206_n2214), 
        .ZN(DP_mult_206_n1260) );
  OR2_X1 DP_mult_206_U2314 ( .A1(DP_mult_206_n1550), .A2(DP_mult_206_n2250), 
        .ZN(DP_mult_206_n2214) );
  OR2_X1 DP_mult_206_U2313 ( .A1(DP_mult_206_n2223), .A2(DP_mult_206_n1551), 
        .ZN(DP_mult_206_n2213) );
  INV_X1 DP_mult_206_U2312 ( .A(DP_mult_206_n508), .ZN(DP_mult_206_n2212) );
  NAND2_X1 DP_mult_206_U2311 ( .A1(DP_mult_206_n1348), .A2(DP_mult_206_n1182), 
        .ZN(DP_mult_206_n2211) );
  NAND2_X1 DP_mult_206_U2310 ( .A1(DP_mult_206_n1260), .A2(DP_mult_206_n1182), 
        .ZN(DP_mult_206_n2210) );
  NAND2_X1 DP_mult_206_U2309 ( .A1(DP_mult_206_n1260), .A2(DP_mult_206_n1348), 
        .ZN(DP_mult_206_n2209) );
  XOR2_X1 DP_mult_206_U2308 ( .A(DP_mult_206_n2128), .B(DP_mult_206_n2208), 
        .Z(DP_mult_206_n959) );
  XOR2_X1 DP_mult_206_U2307 ( .A(DP_mult_206_n1348), .B(DP_mult_206_n1182), 
        .Z(DP_mult_206_n2208) );
  XNOR2_X1 DP_mult_206_U2306 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1567) );
  XNOR2_X1 DP_mult_206_U2305 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1561) );
  XNOR2_X1 DP_mult_206_U2304 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1569) );
  XNOR2_X1 DP_mult_206_U2303 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1563) );
  XNOR2_X1 DP_mult_206_U2302 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1565) );
  XNOR2_X1 DP_mult_206_U2301 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1559) );
  OAI22_X1 DP_mult_206_U2300 ( .A1(DP_mult_206_n2122), .A2(DP_mult_206_n2322), 
        .B1(DP_mult_206_n1531), .B2(DP_mult_206_n2247), .ZN(DP_mult_206_n1183)
         );
  OAI22_X1 DP_mult_206_U2299 ( .A1(DP_mult_206_n2122), .A2(DP_mult_206_n1516), 
        .B1(DP_mult_206_n1515), .B2(DP_mult_206_n2247), .ZN(DP_mult_206_n1226)
         );
  OAI22_X1 DP_mult_206_U2298 ( .A1(DP_mult_206_n2222), .A2(DP_mult_206_n1512), 
        .B1(DP_mult_206_n1511), .B2(DP_mult_206_n2247), .ZN(DP_mult_206_n1222)
         );
  OAI22_X1 DP_mult_206_U2297 ( .A1(DP_mult_206_n2222), .A2(DP_mult_206_n1510), 
        .B1(DP_mult_206_n1509), .B2(DP_mult_206_n2048), .ZN(DP_mult_206_n1220)
         );
  OAI22_X1 DP_mult_206_U2296 ( .A1(DP_mult_206_n2122), .A2(DP_mult_206_n1514), 
        .B1(DP_mult_206_n1513), .B2(DP_mult_206_n2048), .ZN(DP_mult_206_n1224)
         );
  OAI22_X1 DP_mult_206_U2295 ( .A1(DP_mult_206_n2127), .A2(DP_mult_206_n1518), 
        .B1(DP_mult_206_n1517), .B2(DP_mult_206_n2048), .ZN(DP_mult_206_n1228)
         );
  OAI22_X1 DP_mult_206_U2294 ( .A1(DP_mult_206_n2127), .A2(DP_mult_206_n1508), 
        .B1(DP_mult_206_n1507), .B2(DP_mult_206_n2048), .ZN(DP_mult_206_n682)
         );
  INV_X1 DP_mult_206_U2293 ( .A(DP_mult_206_n439), .ZN(DP_mult_206_n445) );
  AOI21_X1 DP_mult_206_U2292 ( .B1(DP_mult_206_n401), .B2(DP_mult_206_n2176), 
        .A(DP_mult_206_n394), .ZN(DP_mult_206_n390) );
  OAI21_X1 DP_mult_206_U2291 ( .B1(DP_mult_206_n390), .B2(DP_mult_206_n384), 
        .A(DP_mult_206_n387), .ZN(DP_mult_206_n383) );
  NAND2_X1 DP_mult_206_U2290 ( .A1(DP_mult_206_n663), .A2(DP_mult_206_n439), 
        .ZN(DP_mult_206_n312) );
  NAND2_X1 DP_mult_206_U2289 ( .A1(DP_mult_206_n2181), .A2(DP_mult_206_n2179), 
        .ZN(DP_mult_206_n599) );
  OAI21_X1 DP_mult_206_U2288 ( .B1(DP_mult_206_n1984), .B2(DP_mult_206_n564), 
        .A(DP_mult_206_n559), .ZN(DP_mult_206_n553) );
  INV_X1 DP_mult_206_U2287 ( .A(DP_mult_206_n2058), .ZN(DP_mult_206_n555) );
  AOI21_X1 DP_mult_206_U2286 ( .B1(DP_mult_206_n1981), .B2(DP_mult_206_n552), 
        .A(DP_mult_206_n2118), .ZN(DP_mult_206_n551) );
  INV_X1 DP_mult_206_U2285 ( .A(DP_mult_206_n772), .ZN(DP_mult_206_n773) );
  NAND3_X1 DP_mult_206_U2284 ( .A1(DP_mult_206_n2205), .A2(DP_mult_206_n2206), 
        .A3(DP_mult_206_n2207), .ZN(DP_mult_206_n974) );
  NAND2_X1 DP_mult_206_U2283 ( .A1(DP_mult_206_n1415), .A2(DP_mult_206_n1393), 
        .ZN(DP_mult_206_n2207) );
  NAND2_X1 DP_mult_206_U2282 ( .A1(DP_mult_206_n1000), .A2(DP_mult_206_n1393), 
        .ZN(DP_mult_206_n2206) );
  NAND2_X1 DP_mult_206_U2281 ( .A1(DP_mult_206_n1000), .A2(DP_mult_206_n1415), 
        .ZN(DP_mult_206_n2205) );
  INV_X1 DP_mult_206_U2280 ( .A(DP_mult_206_n1945), .ZN(DP_mult_206_n565) );
  OAI21_X1 DP_mult_206_U2279 ( .B1(DP_mult_206_n535), .B2(DP_mult_206_n2109), 
        .A(DP_mult_206_n532), .ZN(DP_mult_206_n2204) );
  AOI21_X1 DP_mult_206_U2278 ( .B1(DP_mult_206_n2204), .B2(DP_mult_206_n2124), 
        .A(DP_mult_206_n2131), .ZN(DP_mult_206_n2203) );
  NAND2_X1 DP_mult_206_U2277 ( .A1(DP_mult_206_n666), .A2(DP_mult_206_n1989), 
        .ZN(DP_mult_206_n467) );
  OAI21_X1 DP_mult_206_U2276 ( .B1(DP_mult_206_n555), .B2(DP_mult_206_n2055), 
        .A(DP_mult_206_n550), .ZN(DP_mult_206_n546) );
  INV_X1 DP_mult_206_U2275 ( .A(DP_mult_206_n1933), .ZN(DP_mult_206_n674) );
  NAND2_X1 DP_mult_206_U2274 ( .A1(DP_mult_206_n685), .A2(DP_mult_206_n688), 
        .ZN(DP_mult_206_n369) );
  OAI21_X1 DP_mult_206_U2273 ( .B1(DP_mult_206_n2119), .B2(DP_mult_206_n2121), 
        .A(DP_mult_206_n2338), .ZN(DP_mult_206_n1218) );
  OAI21_X1 DP_mult_206_U2272 ( .B1(DP_mult_206_n2193), .B2(DP_mult_206_n2132), 
        .A(DP_mult_206_n2332), .ZN(DP_mult_206_n1362) );
  OAI21_X1 DP_mult_206_U2271 ( .B1(DP_mult_206_n1990), .B2(DP_mult_206_n2199), 
        .A(DP_mult_206_n2334), .ZN(DP_mult_206_n1314) );
  OAI22_X1 DP_mult_206_U2270 ( .A1(DP_mult_206_n1951), .A2(DP_mult_206_n1949), 
        .B1(DP_mult_206_n1781), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1193)
         );
  OAI21_X1 DP_mult_206_U2269 ( .B1(DP_mult_206_n2196), .B2(DP_mult_206_n2154), 
        .A(DP_mult_206_n2335), .ZN(DP_mult_206_n1290) );
  XNOR2_X1 DP_mult_206_U2268 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2325), .ZN(
        DP_mult_206_n1482) );
  XNOR2_X1 DP_mult_206_U2267 ( .A(DP_mult_206_n448), .B(DP_mult_206_n312), 
        .ZN(DP_pipe0_coeff_pipe00[12]) );
  INV_X1 DP_mult_206_U2266 ( .A(DP_coeffs_ff_int[23]), .ZN(DP_mult_206_n251)
         );
  XNOR2_X1 DP_mult_206_U2265 ( .A(DP_mult_206_n2274), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1780) );
  INV_X1 DP_mult_206_U2264 ( .A(DP_mult_206_n285), .ZN(DP_mult_206_n2232) );
  INV_X1 DP_mult_206_U2263 ( .A(DP_mult_206_n1757), .ZN(DP_mult_206_n2328) );
  OAI21_X1 DP_mult_206_U2262 ( .B1(DP_coeffs_ff_int[23]), .B2(
        DP_mult_206_n2189), .A(DP_mult_206_n2328), .ZN(DP_mult_206_n1458) );
  NAND2_X1 DP_mult_206_U2261 ( .A1(DP_mult_206_n2173), .A2(DP_mult_206_n461), 
        .ZN(DP_mult_206_n313) );
  NAND2_X1 DP_mult_206_U2260 ( .A1(DP_mult_206_n666), .A2(DP_mult_206_n481), 
        .ZN(DP_mult_206_n315) );
  NAND2_X1 DP_mult_206_U2259 ( .A1(DP_mult_206_n667), .A2(DP_mult_206_n496), 
        .ZN(DP_mult_206_n316) );
  NAND2_X1 DP_mult_206_U2258 ( .A1(DP_mult_206_n2049), .A2(DP_mult_206_n514), 
        .ZN(DP_mult_206_n318) );
  NAND2_X1 DP_mult_206_U2257 ( .A1(DP_mult_206_n670), .A2(DP_mult_206_n2063), 
        .ZN(DP_mult_206_n319) );
  NAND2_X1 DP_mult_206_U2256 ( .A1(DP_mult_206_n668), .A2(DP_mult_206_n503), 
        .ZN(DP_mult_206_n317) );
  NAND2_X1 DP_mult_206_U2255 ( .A1(DP_mult_206_n532), .A2(DP_mult_206_n671), 
        .ZN(DP_mult_206_n320) );
  AOI21_X1 DP_mult_206_U2254 ( .B1(DP_mult_206_n565), .B2(DP_mult_206_n545), 
        .A(DP_mult_206_n546), .ZN(DP_mult_206_n544) );
  AOI21_X1 DP_mult_206_U2253 ( .B1(DP_mult_206_n565), .B2(DP_mult_206_n561), 
        .A(DP_mult_206_n562), .ZN(DP_mult_206_n560) );
  XNOR2_X1 DP_mult_206_U2252 ( .A(DP_pipe00[11]), .B(DP_mult_206_n2325), .ZN(
        DP_mult_206_n1494) );
  XNOR2_X1 DP_mult_206_U2251 ( .A(DP_pipe00[21]), .B(DP_mult_206_n2325), .ZN(
        DP_mult_206_n1484) );
  XNOR2_X1 DP_mult_206_U2250 ( .A(DP_pipe00[19]), .B(DP_mult_206_n2325), .ZN(
        DP_mult_206_n1486) );
  XNOR2_X1 DP_mult_206_U2249 ( .A(DP_pipe00[15]), .B(DP_mult_206_n2325), .ZN(
        DP_mult_206_n1490) );
  XNOR2_X1 DP_mult_206_U2248 ( .A(DP_pipe00[17]), .B(DP_mult_206_n2325), .ZN(
        DP_mult_206_n1488) );
  XNOR2_X1 DP_mult_206_U2247 ( .A(DP_pipe00[13]), .B(DP_mult_206_n2324), .ZN(
        DP_mult_206_n1492) );
  XNOR2_X1 DP_mult_206_U2246 ( .A(DP_mult_206_n2299), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1655) );
  XNOR2_X1 DP_mult_206_U2245 ( .A(DP_mult_206_n2284), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1730) );
  XNOR2_X1 DP_mult_206_U2244 ( .A(DP_mult_206_n2312), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1580) );
  XNOR2_X1 DP_mult_206_U2243 ( .A(DP_mult_206_n2324), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1505) );
  XNOR2_X1 DP_mult_206_U2242 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2282), .ZN(
        DP_mult_206_n1725) );
  XNOR2_X1 DP_mult_206_U2241 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2287), .ZN(
        DP_mult_206_n1700) );
  XNOR2_X1 DP_mult_206_U2240 ( .A(DP_pipe00[5]), .B(DP_mult_206_n1985), .ZN(
        DP_mult_206_n1750) );
  XNOR2_X1 DP_mult_206_U2239 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2292), .ZN(
        DP_mult_206_n1675) );
  XNOR2_X1 DP_mult_206_U2238 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2319), .ZN(
        DP_mult_206_n1525) );
  XNOR2_X1 DP_mult_206_U2237 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2297), .ZN(
        DP_mult_206_n1650) );
  XNOR2_X1 DP_mult_206_U2236 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2007), .ZN(
        DP_mult_206_n1625) );
  XNOR2_X1 DP_mult_206_U2235 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1600) );
  XNOR2_X1 DP_mult_206_U2234 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2324), .ZN(
        DP_mult_206_n1500) );
  XNOR2_X1 DP_mult_206_U2233 ( .A(DP_pipe00[5]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1575) );
  XNOR2_X1 DP_mult_206_U2232 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2289), .ZN(
        DP_mult_206_n1704) );
  XNOR2_X1 DP_mult_206_U2231 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2282), .ZN(
        DP_mult_206_n1727) );
  XNOR2_X1 DP_mult_206_U2230 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2299), .ZN(
        DP_mult_206_n1652) );
  XNOR2_X1 DP_mult_206_U2229 ( .A(DP_pipe00[7]), .B(DP_mult_206_n1985), .ZN(
        DP_mult_206_n1748) );
  XNOR2_X1 DP_mult_206_U2228 ( .A(DP_pipe00[3]), .B(DP_mult_206_n1985), .ZN(
        DP_mult_206_n1752) );
  XNOR2_X1 DP_mult_206_U2227 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2292), .ZN(
        DP_mult_206_n1677) );
  XNOR2_X1 DP_mult_206_U2226 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2282), .ZN(
        DP_mult_206_n1729) );
  XNOR2_X1 DP_mult_206_U2225 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2289), .ZN(
        DP_mult_206_n1698) );
  XNOR2_X1 DP_mult_206_U2224 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2319), .ZN(
        DP_mult_206_n1523) );
  XNOR2_X1 DP_mult_206_U2223 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2007), .ZN(
        DP_mult_206_n1629) );
  XNOR2_X1 DP_mult_206_U2222 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2293), .ZN(
        DP_mult_206_n1679) );
  XNOR2_X1 DP_mult_206_U2221 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1552) );
  XNOR2_X1 DP_mult_206_U2220 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2299), .ZN(
        DP_mult_206_n1654) );
  XNOR2_X1 DP_mult_206_U2219 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2289), .ZN(
        DP_mult_206_n1702) );
  XNOR2_X1 DP_mult_206_U2218 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2292), .ZN(
        DP_mult_206_n1673) );
  XNOR2_X1 DP_mult_206_U2217 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2319), .ZN(
        DP_mult_206_n1529) );
  XNOR2_X1 DP_mult_206_U2216 ( .A(DP_pipe00[1]), .B(DP_mult_206_n1985), .ZN(
        DP_mult_206_n1754) );
  XNOR2_X1 DP_mult_206_U2215 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1604) );
  XNOR2_X1 DP_mult_206_U2214 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2282), .ZN(
        DP_mult_206_n1723) );
  XNOR2_X1 DP_mult_206_U2213 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2302), .ZN(
        DP_mult_206_n1627) );
  XNOR2_X1 DP_mult_206_U2212 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2298), .ZN(
        DP_mult_206_n1648) );
  XNOR2_X1 DP_mult_206_U2211 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1602) );
  XNOR2_X1 DP_mult_206_U2210 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1579) );
  XNOR2_X1 DP_mult_206_U2209 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1577) );
  XNOR2_X1 DP_mult_206_U2208 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1554) );
  XNOR2_X1 DP_mult_206_U2207 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2302), .ZN(
        DP_mult_206_n1623) );
  XNOR2_X1 DP_mult_206_U2206 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1598) );
  XNOR2_X1 DP_mult_206_U2205 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1548) );
  XNOR2_X1 DP_mult_206_U2204 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2324), .ZN(
        DP_mult_206_n1502) );
  XNOR2_X1 DP_mult_206_U2203 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2324), .ZN(
        DP_mult_206_n1498) );
  XNOR2_X1 DP_mult_206_U2202 ( .A(DP_pipe00[7]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1573) );
  XNOR2_X1 DP_mult_206_U2201 ( .A(DP_pipe00[3]), .B(DP_mult_206_n2319), .ZN(
        DP_mult_206_n1527) );
  XNOR2_X1 DP_mult_206_U2200 ( .A(DP_pipe00[1]), .B(DP_mult_206_n2324), .ZN(
        DP_mult_206_n1504) );
  XNOR2_X1 DP_mult_206_U2199 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2319), .ZN(
        DP_mult_206_n1521) );
  XNOR2_X1 DP_mult_206_U2198 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1771) );
  XNOR2_X1 DP_mult_206_U2197 ( .A(DP_pipe00[9]), .B(DP_mult_206_n1985), .ZN(
        DP_mult_206_n1746) );
  XNOR2_X1 DP_mult_206_U2196 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2282), .ZN(
        DP_mult_206_n1721) );
  XNOR2_X1 DP_mult_206_U2195 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2288), .ZN(
        DP_mult_206_n1696) );
  XNOR2_X1 DP_mult_206_U2194 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2292), .ZN(
        DP_mult_206_n1671) );
  XNOR2_X1 DP_mult_206_U2193 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2298), .ZN(
        DP_mult_206_n1646) );
  XNOR2_X1 DP_mult_206_U2192 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2324), .ZN(
        DP_mult_206_n1496) );
  XNOR2_X1 DP_mult_206_U2191 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2007), .ZN(
        DP_mult_206_n1621) );
  XNOR2_X1 DP_mult_206_U2190 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1546) );
  XNOR2_X1 DP_mult_206_U2189 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1596) );
  XNOR2_X1 DP_mult_206_U2188 ( .A(DP_pipe00[9]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1571) );
  XNOR2_X1 DP_mult_206_U2187 ( .A(DP_mult_206_n2287), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1705) );
  XNOR2_X1 DP_mult_206_U2186 ( .A(DP_mult_206_n2316), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1555) );
  XNOR2_X1 DP_mult_206_U2185 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2319), .ZN(
        DP_mult_206_n1507) );
  XNOR2_X1 DP_mult_206_U2184 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2314), .ZN(
        DP_mult_206_n1532) );
  XNOR2_X1 DP_mult_206_U2183 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2307), .ZN(
        DP_mult_206_n1582) );
  XNOR2_X1 DP_mult_206_U2182 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2038), .ZN(
        DP_mult_206_n1557) );
  XNOR2_X1 DP_mult_206_U2181 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2007), .ZN(
        DP_mult_206_n1607) );
  XNOR2_X1 DP_mult_206_U2180 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2298), .ZN(
        DP_mult_206_n1632) );
  XNOR2_X1 DP_mult_206_U2179 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2292), .ZN(
        DP_mult_206_n1657) );
  XNOR2_X1 DP_mult_206_U2178 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2277), .ZN(
        DP_mult_206_n1732) );
  XNOR2_X1 DP_mult_206_U2177 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2282), .ZN(
        DP_mult_206_n1707) );
  XNOR2_X1 DP_mult_206_U2176 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2287), .ZN(
        DP_mult_206_n1682) );
  XNOR2_X1 DP_mult_206_U2175 ( .A(DP_mult_206_n2287), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1701) );
  XNOR2_X1 DP_mult_206_U2174 ( .A(DP_mult_206_n2303), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1626) );
  XNOR2_X1 DP_mult_206_U2173 ( .A(DP_mult_206_n2278), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1751) );
  XNOR2_X1 DP_mult_206_U2172 ( .A(DP_mult_206_n2299), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1651) );
  XNOR2_X1 DP_mult_206_U2171 ( .A(DP_mult_206_n2283), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1726) );
  XNOR2_X1 DP_mult_206_U2170 ( .A(DP_mult_206_n2293), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1676) );
  XNOR2_X1 DP_mult_206_U2169 ( .A(DP_mult_206_n2320), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1526) );
  XNOR2_X1 DP_mult_206_U2168 ( .A(DP_mult_206_n2308), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1601) );
  XNOR2_X1 DP_mult_206_U2167 ( .A(DP_mult_206_n2311), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1576) );
  XNOR2_X1 DP_mult_206_U2166 ( .A(DP_mult_206_n2324), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1501) );
  XNOR2_X1 DP_mult_206_U2165 ( .A(DP_mult_206_n2273), .B(DP_pipe00[4]), .ZN(
        DP_mult_206_n1776) );
  XNOR2_X1 DP_mult_206_U2164 ( .A(DP_mult_206_n2278), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1747) );
  XNOR2_X1 DP_mult_206_U2163 ( .A(DP_mult_206_n2278), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1753) );
  XNOR2_X1 DP_mult_206_U2162 ( .A(DP_mult_206_n2278), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1749) );
  XNOR2_X1 DP_mult_206_U2161 ( .A(DP_mult_206_n2320), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1522) );
  XNOR2_X1 DP_mult_206_U2160 ( .A(DP_mult_206_n2288), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1699) );
  XNOR2_X1 DP_mult_206_U2159 ( .A(DP_mult_206_n2283), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1728) );
  XNOR2_X1 DP_mult_206_U2158 ( .A(DP_mult_206_n2288), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1703) );
  XNOR2_X1 DP_mult_206_U2157 ( .A(DP_mult_206_n2298), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1653) );
  XNOR2_X1 DP_mult_206_U2156 ( .A(DP_mult_206_n2298), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1649) );
  XNOR2_X1 DP_mult_206_U2155 ( .A(DP_mult_206_n2308), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1603) );
  XNOR2_X1 DP_mult_206_U2154 ( .A(DP_mult_206_n2320), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1524) );
  XNOR2_X1 DP_mult_206_U2153 ( .A(DP_mult_206_n2287), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1697) );
  XNOR2_X1 DP_mult_206_U2152 ( .A(DP_mult_206_n2283), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1722) );
  XNOR2_X1 DP_mult_206_U2151 ( .A(DP_mult_206_n2293), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1672) );
  XNOR2_X1 DP_mult_206_U2150 ( .A(DP_mult_206_n2293), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1678) );
  XNOR2_X1 DP_mult_206_U2149 ( .A(DP_mult_206_n2293), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1674) );
  XNOR2_X1 DP_mult_206_U2148 ( .A(DP_mult_206_n2303), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1628) );
  XNOR2_X1 DP_mult_206_U2147 ( .A(DP_mult_206_n2283), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1724) );
  XNOR2_X1 DP_mult_206_U2146 ( .A(DP_mult_206_n2303), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1624) );
  XNOR2_X1 DP_mult_206_U2145 ( .A(DP_mult_206_n2298), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1647) );
  XNOR2_X1 DP_mult_206_U2144 ( .A(DP_mult_206_n2315), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1553) );
  XNOR2_X1 DP_mult_206_U2143 ( .A(DP_mult_206_n2311), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1578) );
  XNOR2_X1 DP_mult_206_U2142 ( .A(DP_mult_206_n2303), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1622) );
  XNOR2_X1 DP_mult_206_U2141 ( .A(DP_mult_206_n2308), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1599) );
  XNOR2_X1 DP_mult_206_U2140 ( .A(DP_mult_206_n2324), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1497) );
  XNOR2_X1 DP_mult_206_U2139 ( .A(DP_mult_206_n2315), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1547) );
  XNOR2_X1 DP_mult_206_U2138 ( .A(DP_mult_206_n2311), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1574) );
  XNOR2_X1 DP_mult_206_U2137 ( .A(DP_mult_206_n2308), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1597) );
  XNOR2_X1 DP_mult_206_U2136 ( .A(DP_mult_206_n2324), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1499) );
  XNOR2_X1 DP_mult_206_U2135 ( .A(DP_mult_206_n2315), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1549) );
  XNOR2_X1 DP_mult_206_U2134 ( .A(DP_mult_206_n2324), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1503) );
  XNOR2_X1 DP_mult_206_U2133 ( .A(DP_mult_206_n2311), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1572) );
  XNOR2_X1 DP_mult_206_U2132 ( .A(DP_mult_206_n2320), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1528) );
  XNOR2_X1 DP_mult_206_U2131 ( .A(DP_mult_206_n2273), .B(DP_pipe00[8]), .ZN(
        DP_mult_206_n1772) );
  XNOR2_X1 DP_mult_206_U2130 ( .A(DP_mult_206_n2273), .B(DP_pipe00[6]), .ZN(
        DP_mult_206_n1774) );
  XNOR2_X1 DP_mult_206_U2129 ( .A(DP_mult_206_n2273), .B(DP_pipe00[2]), .ZN(
        DP_mult_206_n1778) );
  XNOR2_X1 DP_mult_206_U2128 ( .A(DP_pipe00[23]), .B(DP_mult_206_n2272), .ZN(
        DP_mult_206_n1757) );
  XNOR2_X1 DP_mult_206_U2127 ( .A(DP_mult_206_n2325), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1483) );
  XNOR2_X1 DP_mult_206_U2126 ( .A(DP_mult_206_n2316), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1535) );
  XNOR2_X1 DP_mult_206_U2125 ( .A(DP_mult_206_n2325), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1485) );
  XNOR2_X1 DP_mult_206_U2124 ( .A(DP_mult_206_n2325), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1487) );
  XNOR2_X1 DP_mult_206_U2123 ( .A(DP_mult_206_n2312), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1560) );
  XNOR2_X1 DP_mult_206_U2122 ( .A(DP_mult_206_n2320), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1520) );
  XNOR2_X1 DP_mult_206_U2121 ( .A(DP_mult_206_n2320), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1518) );
  XNOR2_X1 DP_mult_206_U2120 ( .A(DP_mult_206_n2316), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1533) );
  XNOR2_X1 DP_mult_206_U2119 ( .A(DP_mult_206_n2311), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1562) );
  XNOR2_X1 DP_mult_206_U2118 ( .A(DP_mult_206_n2309), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1583) );
  XNOR2_X1 DP_mult_206_U2117 ( .A(DP_mult_206_n2325), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1489) );
  XNOR2_X1 DP_mult_206_U2116 ( .A(DP_mult_206_n2325), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1493) );
  XNOR2_X1 DP_mult_206_U2115 ( .A(DP_mult_206_n2278), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1745) );
  XNOR2_X1 DP_mult_206_U2114 ( .A(DP_mult_206_n2315), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1537) );
  XNOR2_X1 DP_mult_206_U2113 ( .A(DP_mult_206_n2283), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1720) );
  XNOR2_X1 DP_mult_206_U2112 ( .A(DP_mult_206_n2309), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1585) );
  XNOR2_X1 DP_mult_206_U2111 ( .A(DP_mult_206_n2316), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1539) );
  XNOR2_X1 DP_mult_206_U2110 ( .A(DP_mult_206_n2312), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1558) );
  XNOR2_X1 DP_mult_206_U2109 ( .A(DP_mult_206_n2325), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1491) );
  XNOR2_X1 DP_mult_206_U2108 ( .A(DP_mult_206_n2278), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1741) );
  XNOR2_X1 DP_mult_206_U2107 ( .A(DP_mult_206_n2278), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1743) );
  XNOR2_X1 DP_mult_206_U2106 ( .A(DP_mult_206_n2304), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1608) );
  XNOR2_X1 DP_mult_206_U2105 ( .A(DP_mult_206_n2289), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1695) );
  XNOR2_X1 DP_mult_206_U2104 ( .A(DP_mult_206_n2283), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1718) );
  XNOR2_X1 DP_mult_206_U2103 ( .A(DP_mult_206_n2293), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1670) );
  XNOR2_X1 DP_mult_206_U2102 ( .A(DP_mult_206_n2298), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1633) );
  XNOR2_X1 DP_mult_206_U2101 ( .A(DP_mult_206_n2288), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1693) );
  XNOR2_X1 DP_mult_206_U2100 ( .A(DP_mult_206_n2279), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1739) );
  XNOR2_X1 DP_mult_206_U2099 ( .A(DP_mult_206_n2283), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1716) );
  XNOR2_X1 DP_mult_206_U2098 ( .A(DP_mult_206_n2298), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1645) );
  XNOR2_X1 DP_mult_206_U2097 ( .A(DP_mult_206_n2284), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1714) );
  XNOR2_X1 DP_mult_206_U2096 ( .A(DP_mult_206_n2293), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1668) );
  XNOR2_X1 DP_mult_206_U2095 ( .A(DP_mult_206_n2312), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1564) );
  XNOR2_X1 DP_mult_206_U2094 ( .A(DP_mult_206_n2308), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1587) );
  XNOR2_X1 DP_mult_206_U2093 ( .A(DP_mult_206_n2287), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1683) );
  XNOR2_X1 DP_mult_206_U2092 ( .A(DP_mult_206_n2284), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1708) );
  XNOR2_X1 DP_mult_206_U2091 ( .A(DP_mult_206_n2278), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1737) );
  XNOR2_X1 DP_mult_206_U2090 ( .A(DP_mult_206_n2304), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1610) );
  XNOR2_X1 DP_mult_206_U2089 ( .A(DP_mult_206_n2297), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1637) );
  XNOR2_X1 DP_mult_206_U2088 ( .A(DP_mult_206_n2289), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1691) );
  XNOR2_X1 DP_mult_206_U2087 ( .A(DP_mult_206_n2303), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1620) );
  XNOR2_X1 DP_mult_206_U2086 ( .A(DP_mult_206_n2325), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1495) );
  XNOR2_X1 DP_mult_206_U2085 ( .A(DP_mult_206_n2315), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1541) );
  XNOR2_X1 DP_mult_206_U2084 ( .A(DP_mult_206_n2303), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1612) );
  XNOR2_X1 DP_mult_206_U2083 ( .A(DP_mult_206_n2303), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1616) );
  XNOR2_X1 DP_mult_206_U2082 ( .A(DP_mult_206_n2279), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1735) );
  XNOR2_X1 DP_mult_206_U2081 ( .A(DP_mult_206_n2293), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1666) );
  XNOR2_X1 DP_mult_206_U2080 ( .A(DP_mult_206_n2289), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1689) );
  XNOR2_X1 DP_mult_206_U2079 ( .A(DP_mult_206_n2294), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1658) );
  XNOR2_X1 DP_mult_206_U2078 ( .A(DP_mult_206_n2308), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1591) );
  XNOR2_X1 DP_mult_206_U2077 ( .A(DP_mult_206_n2283), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1712) );
  XNOR2_X1 DP_mult_206_U2076 ( .A(DP_mult_206_n2284), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1710) );
  XNOR2_X1 DP_mult_206_U2075 ( .A(DP_mult_206_n2311), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1566) );
  XNOR2_X1 DP_mult_206_U2074 ( .A(DP_mult_206_n2309), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1589) );
  XNOR2_X1 DP_mult_206_U2073 ( .A(DP_mult_206_n2298), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1643) );
  XNOR2_X1 DP_mult_206_U2072 ( .A(DP_mult_206_n2297), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1639) );
  XNOR2_X1 DP_mult_206_U2071 ( .A(DP_mult_206_n2294), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1660) );
  XNOR2_X1 DP_mult_206_U2070 ( .A(DP_mult_206_n2311), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1568) );
  XNOR2_X1 DP_mult_206_U2069 ( .A(DP_mult_206_n2293), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1662) );
  XNOR2_X1 DP_mult_206_U2068 ( .A(DP_mult_206_n2311), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1570) );
  XNOR2_X1 DP_mult_206_U2067 ( .A(DP_mult_206_n2288), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1685) );
  XNOR2_X1 DP_mult_206_U2066 ( .A(DP_mult_206_n2315), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1545) );
  XNOR2_X1 DP_mult_206_U2065 ( .A(DP_mult_206_n2304), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1614) );
  XNOR2_X1 DP_mult_206_U2064 ( .A(DP_mult_206_n2279), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1733) );
  XNOR2_X1 DP_mult_206_U2063 ( .A(DP_mult_206_n2298), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1635) );
  XNOR2_X1 DP_mult_206_U2062 ( .A(DP_mult_206_n2315), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1543) );
  XNOR2_X1 DP_mult_206_U2061 ( .A(DP_mult_206_n2297), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1641) );
  XNOR2_X1 DP_mult_206_U2060 ( .A(DP_mult_206_n2303), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1618) );
  XNOR2_X1 DP_mult_206_U2059 ( .A(DP_mult_206_n2308), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1595) );
  XNOR2_X1 DP_mult_206_U2058 ( .A(DP_mult_206_n2308), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1593) );
  XNOR2_X1 DP_mult_206_U2057 ( .A(DP_mult_206_n2289), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1687) );
  XNOR2_X1 DP_mult_206_U2056 ( .A(DP_mult_206_n2294), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1664) );
  XNOR2_X1 DP_mult_206_U2055 ( .A(DP_mult_206_n2273), .B(DP_pipe00[10]), .ZN(
        DP_mult_206_n1770) );
  XNOR2_X1 DP_mult_206_U2054 ( .A(DP_mult_206_n2321), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1508) );
  XNOR2_X1 DP_mult_206_U2053 ( .A(DP_mult_206_n2321), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1510) );
  XNOR2_X1 DP_mult_206_U2052 ( .A(DP_mult_206_n2321), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1514) );
  XNOR2_X1 DP_mult_206_U2051 ( .A(DP_mult_206_n2320), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1512) );
  XNOR2_X1 DP_mult_206_U2050 ( .A(DP_mult_206_n2320), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1516) );
  XNOR2_X1 DP_mult_206_U2049 ( .A(DP_mult_206_n2273), .B(DP_pipe00[12]), .ZN(
        DP_mult_206_n1768) );
  XNOR2_X1 DP_mult_206_U2048 ( .A(DP_mult_206_n2274), .B(DP_pipe00[16]), .ZN(
        DP_mult_206_n1764) );
  XNOR2_X1 DP_mult_206_U2047 ( .A(DP_mult_206_n2273), .B(DP_pipe00[14]), .ZN(
        DP_mult_206_n1766) );
  XNOR2_X1 DP_mult_206_U2046 ( .A(DP_mult_206_n2273), .B(DP_pipe00[18]), .ZN(
        DP_mult_206_n1762) );
  XNOR2_X1 DP_mult_206_U2045 ( .A(DP_mult_206_n2274), .B(DP_pipe00[20]), .ZN(
        DP_mult_206_n1760) );
  XNOR2_X1 DP_mult_206_U2044 ( .A(DP_mult_206_n2274), .B(DP_pipe00[22]), .ZN(
        DP_mult_206_n1758) );
  XNOR2_X1 DP_mult_206_U2043 ( .A(DP_mult_206_n2294), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1680) );
  XNOR2_X1 DP_mult_206_U2042 ( .A(DP_mult_206_n2304), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1630) );
  XNOR2_X1 DP_mult_206_U2041 ( .A(DP_mult_206_n2279), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1755) );
  XNOR2_X1 DP_mult_206_U2040 ( .A(DP_mult_206_n2309), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1605) );
  XNOR2_X1 DP_mult_206_U2039 ( .A(DP_mult_206_n2321), .B(DP_pipe00[0]), .ZN(
        DP_mult_206_n1530) );
  INV_X1 DP_mult_206_U2038 ( .A(DP_mult_206_n1482), .ZN(DP_mult_206_n2339) );
  INV_X1 DP_mult_206_U2037 ( .A(DP_mult_206_n1582), .ZN(DP_mult_206_n2335) );
  INV_X1 DP_mult_206_U2036 ( .A(DP_mult_206_n1657), .ZN(DP_mult_206_n2332) );
  INV_X1 DP_mult_206_U2035 ( .A(DP_mult_206_n1732), .ZN(DP_mult_206_n2329) );
  INV_X1 DP_mult_206_U2034 ( .A(DP_mult_206_n802), .ZN(DP_mult_206_n803) );
  OAI22_X1 DP_mult_206_U2033 ( .A1(DP_mult_206_n1951), .A2(DP_mult_206_n1767), 
        .B1(DP_mult_206_n1766), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1468)
         );
  INV_X1 DP_mult_206_U2032 ( .A(DP_mult_206_n1607), .ZN(DP_mult_206_n2334) );
  INV_X1 DP_mult_206_U2031 ( .A(DP_mult_206_n1557), .ZN(DP_mult_206_n2336) );
  OAI21_X1 DP_mult_206_U2030 ( .B1(DP_mult_206_n2195), .B2(DP_mult_206_n2108), 
        .A(DP_mult_206_n2336), .ZN(DP_mult_206_n1266) );
  OAI22_X1 DP_mult_206_U2029 ( .A1(DP_mult_206_n1951), .A2(DP_mult_206_n1764), 
        .B1(DP_mult_206_n1763), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1465)
         );
  XNOR2_X1 DP_mult_206_U2028 ( .A(DP_mult_206_n1415), .B(DP_mult_206_n1393), 
        .ZN(DP_mult_206_n2188) );
  XNOR2_X1 DP_mult_206_U2027 ( .A(DP_mult_206_n1000), .B(DP_mult_206_n2188), 
        .ZN(DP_mult_206_n975) );
  INV_X1 DP_mult_206_U2026 ( .A(DP_mult_206_n874), .ZN(DP_mult_206_n875) );
  NOR2_X1 DP_mult_206_U2025 ( .A1(DP_mult_206_n2257), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1337) );
  NOR2_X1 DP_mult_206_U2024 ( .A1(DP_mult_206_n2253), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1289) );
  INV_X1 DP_mult_206_U2023 ( .A(DP_mult_206_n724), .ZN(DP_mult_206_n725) );
  OAI22_X1 DP_mult_206_U2022 ( .A1(DP_mult_206_n2122), .A2(DP_mult_206_n1513), 
        .B1(DP_mult_206_n2247), .B2(DP_mult_206_n1512), .ZN(DP_mult_206_n1223)
         );
  OAI22_X1 DP_mult_206_U2021 ( .A1(DP_mult_206_n1950), .A2(DP_mult_206_n1765), 
        .B1(DP_mult_206_n1764), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1466)
         );
  INV_X1 DP_mult_206_U2020 ( .A(DP_mult_206_n1707), .ZN(DP_mult_206_n2330) );
  OAI22_X1 DP_mult_206_U2019 ( .A1(DP_mult_206_n2242), .A2(DP_mult_206_n1768), 
        .B1(DP_mult_206_n1767), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1469)
         );
  NOR2_X1 DP_mult_206_U2018 ( .A1(DP_mult_206_n2247), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1241) );
  NOR2_X1 DP_mult_206_U2017 ( .A1(DP_mult_206_n2056), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1361) );
  NOR2_X1 DP_mult_206_U2016 ( .A1(DP_mult_206_n2249), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1265) );
  OAI22_X1 DP_mult_206_U2015 ( .A1(DP_mult_206_n2122), .A2(DP_mult_206_n1517), 
        .B1(DP_mult_206_n2048), .B2(DP_mult_206_n1516), .ZN(DP_mult_206_n1227)
         );
  INV_X1 DP_mult_206_U2014 ( .A(DP_mult_206_n1682), .ZN(DP_mult_206_n2331) );
  OAI22_X1 DP_mult_206_U2013 ( .A1(DP_mult_206_n2122), .A2(DP_mult_206_n1509), 
        .B1(DP_mult_206_n2247), .B2(DP_mult_206_n1508), .ZN(DP_mult_206_n1219)
         );
  OAI22_X1 DP_mult_206_U2012 ( .A1(DP_mult_206_n2241), .A2(DP_mult_206_n1759), 
        .B1(DP_mult_206_n1758), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1460)
         );
  NOR2_X1 DP_mult_206_U2011 ( .A1(DP_mult_206_n2255), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1313) );
  OAI22_X1 DP_mult_206_U2010 ( .A1(DP_mult_206_n2242), .A2(DP_mult_206_n1763), 
        .B1(DP_mult_206_n1762), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1464)
         );
  NOR2_X1 DP_mult_206_U2009 ( .A1(DP_mult_206_n1986), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1217) );
  OAI22_X1 DP_mult_206_U2008 ( .A1(DP_mult_206_n2127), .A2(DP_mult_206_n1511), 
        .B1(DP_mult_206_n2048), .B2(DP_mult_206_n1510), .ZN(DP_mult_206_n1221)
         );
  NOR2_X1 DP_mult_206_U2007 ( .A1(DP_mult_206_n2039), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1409) );
  INV_X1 DP_mult_206_U2006 ( .A(DP_mult_206_n1532), .ZN(DP_mult_206_n2337) );
  OAI21_X1 DP_mult_206_U2005 ( .B1(DP_mult_206_n1943), .B2(DP_mult_206_n1991), 
        .A(DP_mult_206_n2337), .ZN(DP_mult_206_n1242) );
  INV_X1 DP_mult_206_U2004 ( .A(DP_mult_206_n1632), .ZN(DP_mult_206_n2333) );
  INV_X1 DP_mult_206_U2003 ( .A(DP_mult_206_n692), .ZN(DP_mult_206_n693) );
  NOR2_X1 DP_mult_206_U2002 ( .A1(DP_mult_206_n1181), .A2(DP_mult_206_n1192), 
        .ZN(DP_mult_206_n644) );
  NAND2_X1 DP_mult_206_U2001 ( .A1(DP_mult_206_n1181), .A2(DP_mult_206_n1192), 
        .ZN(DP_mult_206_n645) );
  NAND2_X1 DP_mult_206_U2000 ( .A1(DP_mult_206_n2315), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1556) );
  NAND2_X1 DP_mult_206_U1999 ( .A1(DP_mult_206_n2311), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1581) );
  NAND2_X1 DP_mult_206_U1998 ( .A1(DP_mult_206_n2288), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1706) );
  NAND2_X1 DP_mult_206_U1997 ( .A1(DP_mult_206_n2273), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1781) );
  NAND2_X1 DP_mult_206_U1996 ( .A1(DP_mult_206_n2303), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1631) );
  NAND2_X1 DP_mult_206_U1995 ( .A1(DP_mult_206_n2308), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1606) );
  NAND2_X1 DP_mult_206_U1994 ( .A1(DP_mult_206_n2298), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1656) );
  NAND2_X1 DP_mult_206_U1993 ( .A1(DP_mult_206_n2325), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1506) );
  AOI21_X1 DP_mult_206_U1992 ( .B1(DP_mult_206_n1965), .B2(DP_mult_206_n1964), 
        .A(DP_mult_206_n1971), .ZN(DP_mult_206_n646) );
  NAND2_X1 DP_mult_206_U1991 ( .A1(DP_mult_206_n2320), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1531) );
  NAND2_X1 DP_mult_206_U1990 ( .A1(DP_mult_206_n2293), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1681) );
  NOR2_X1 DP_mult_206_U1989 ( .A1(DP_mult_206_n2264), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1433) );
  INV_X1 DP_mult_206_U1988 ( .A(DP_mult_206_n1990), .ZN(DP_mult_206_n2257) );
  INV_X1 DP_mult_206_U1987 ( .A(DP_mult_206_n2190), .ZN(DP_mult_206_n2244) );
  INV_X1 DP_mult_206_U1986 ( .A(DP_mult_206_n1943), .ZN(DP_mult_206_n2224) );
  NOR2_X1 DP_mult_206_U1985 ( .A1(DP_mult_206_n2260), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1385) );
  NAND2_X1 DP_mult_206_U1984 ( .A1(DP_mult_206_n2283), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1731) );
  INV_X1 DP_mult_206_U1983 ( .A(DP_mult_206_n682), .ZN(DP_mult_206_n683) );
  INV_X1 DP_mult_206_U1982 ( .A(DP_mult_206_n1507), .ZN(DP_mult_206_n2338) );
  OAI22_X1 DP_mult_206_U1981 ( .A1(DP_mult_206_n2241), .A2(DP_mult_206_n1766), 
        .B1(DP_mult_206_n1765), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1467)
         );
  OAI22_X1 DP_mult_206_U1980 ( .A1(DP_mult_206_n1950), .A2(DP_mult_206_n1760), 
        .B1(DP_mult_206_n1759), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1461)
         );
  OAI22_X1 DP_mult_206_U1979 ( .A1(DP_mult_206_n2122), .A2(DP_mult_206_n1515), 
        .B1(DP_mult_206_n2247), .B2(DP_mult_206_n1514), .ZN(DP_mult_206_n1225)
         );
  OAI22_X1 DP_mult_206_U1978 ( .A1(DP_mult_206_n1951), .A2(DP_mult_206_n1761), 
        .B1(DP_mult_206_n1760), .B2(DP_mult_206_n2269), .ZN(DP_mult_206_n1462)
         );
  OAI22_X1 DP_mult_206_U1977 ( .A1(DP_mult_206_n1950), .A2(DP_mult_206_n1758), 
        .B1(DP_mult_206_n1757), .B2(DP_mult_206_n2269), .ZN(DP_mult_206_n1459)
         );
  OAI22_X1 DP_mult_206_U1976 ( .A1(DP_mult_206_n2242), .A2(DP_mult_206_n1762), 
        .B1(DP_mult_206_n1761), .B2(DP_mult_206_n2270), .ZN(DP_mult_206_n1463)
         );
  NOR2_X1 DP_mult_206_U1975 ( .A1(DP_mult_206_n2265), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1457) );
  INV_X1 DP_mult_206_U1974 ( .A(DP_mult_206_n2276), .ZN(DP_mult_206_n2273) );
  INV_X1 DP_mult_206_U1973 ( .A(DP_mult_206_n2281), .ZN(DP_mult_206_n2278) );
  NAND2_X1 DP_mult_206_U1972 ( .A1(DP_mult_206_n2278), .A2(DP_mult_206_n2327), 
        .ZN(DP_mult_206_n1756) );
  AND2_X1 DP_mult_206_U1971 ( .A1(DP_mult_206_n1194), .A2(DP_mult_206_n676), 
        .ZN(DP_mult_206_n2187) );
  OR2_X1 DP_mult_206_U1970 ( .A1(DP_mult_206_n1194), .A2(DP_mult_206_n676), 
        .ZN(DP_mult_206_n2186) );
  NAND2_X1 DP_mult_206_U1969 ( .A1(DP_mult_206_n1159), .A2(DP_mult_206_n1161), 
        .ZN(DP_mult_206_n627) );
  NAND2_X1 DP_mult_206_U1968 ( .A1(DP_mult_206_n1175), .A2(DP_mult_206_n1178), 
        .ZN(DP_mult_206_n637) );
  NAND2_X1 DP_mult_206_U1967 ( .A1(DP_mult_206_n679), .A2(DP_mult_206_n680), 
        .ZN(DP_mult_206_n341) );
  NAND2_X1 DP_mult_206_U1966 ( .A1(DP_mult_206_n681), .A2(DP_mult_206_n684), 
        .ZN(DP_mult_206_n352) );
  OR2_X1 DP_mult_206_U1965 ( .A1(DP_mult_206_n679), .A2(DP_mult_206_n680), 
        .ZN(DP_mult_206_n2185) );
  NOR2_X1 DP_mult_206_U1964 ( .A1(DP_mult_206_n678), .A2(DP_mult_206_n677), 
        .ZN(DP_mult_206_n334) );
  NOR2_X1 DP_mult_206_U1963 ( .A1(DP_mult_206_n1175), .A2(DP_mult_206_n1178), 
        .ZN(DP_mult_206_n636) );
  NOR2_X1 DP_mult_206_U1962 ( .A1(DP_mult_206_n1159), .A2(DP_mult_206_n1161), 
        .ZN(DP_mult_206_n626) );
  INV_X1 DP_mult_206_U1961 ( .A(DP_mult_206_n341), .ZN(DP_mult_206_n339) );
  NAND2_X1 DP_mult_206_U1960 ( .A1(DP_mult_206_n678), .A2(DP_mult_206_n677), 
        .ZN(DP_mult_206_n335) );
  OR2_X1 DP_mult_206_U1959 ( .A1(DP_mult_206_n681), .A2(DP_mult_206_n684), 
        .ZN(DP_mult_206_n2184) );
  OAI21_X1 DP_mult_206_U1958 ( .B1(DP_mult_206_n646), .B2(DP_mult_206_n644), 
        .A(DP_mult_206_n645), .ZN(DP_mult_206_n643) );
  AOI21_X1 DP_mult_206_U1957 ( .B1(DP_mult_206_n643), .B2(DP_mult_206_n1967), 
        .A(DP_mult_206_n1973), .ZN(DP_mult_206_n638) );
  OR2_X1 DP_mult_206_U1956 ( .A1(DP_mult_206_n685), .A2(DP_mult_206_n688), 
        .ZN(DP_mult_206_n2183) );
  INV_X1 DP_mult_206_U1955 ( .A(DP_mult_206_n676), .ZN(DP_mult_206_n677) );
  AOI21_X1 DP_mult_206_U1954 ( .B1(DP_mult_206_n2181), .B2(DP_mult_206_n1969), 
        .A(DP_mult_206_n1976), .ZN(DP_mult_206_n600) );
  NAND2_X1 DP_mult_206_U1953 ( .A1(DP_mult_206_n2184), .A2(DP_mult_206_n352), 
        .ZN(DP_mult_206_n303) );
  NAND2_X1 DP_mult_206_U1952 ( .A1(DP_mult_206_n2185), .A2(DP_mult_206_n341), 
        .ZN(DP_mult_206_n302) );
  NAND2_X1 DP_mult_206_U1951 ( .A1(DP_mult_206_n2183), .A2(DP_mult_206_n369), 
        .ZN(DP_mult_206_n304) );
  NOR2_X1 DP_mult_206_U1950 ( .A1(DP_mult_206_n336), .A2(DP_mult_206_n334), 
        .ZN(DP_mult_206_n332) );
  NAND2_X1 DP_mult_206_U1949 ( .A1(DP_mult_206_n2170), .A2(DP_mult_206_n2180), 
        .ZN(DP_mult_206_n610) );
  NAND2_X1 DP_mult_206_U1948 ( .A1(DP_mult_206_n694), .A2(DP_mult_206_n689), 
        .ZN(DP_mult_206_n378) );
  INV_X1 DP_mult_206_U1947 ( .A(DP_mult_206_n369), .ZN(DP_mult_206_n367) );
  NAND2_X1 DP_mult_206_U1946 ( .A1(DP_mult_206_n1085), .A2(DP_mult_206_n1098), 
        .ZN(DP_mult_206_n593) );
  OR2_X1 DP_mult_206_U1945 ( .A1(DP_mult_206_n694), .A2(DP_mult_206_n689), 
        .ZN(DP_mult_206_n2182) );
  NAND2_X1 DP_mult_206_U1944 ( .A1(DP_mult_206_n701), .A2(DP_mult_206_n708), 
        .ZN(DP_mult_206_n396) );
  NAND2_X1 DP_mult_206_U1943 ( .A1(DP_mult_206_n695), .A2(DP_mult_206_n700), 
        .ZN(DP_mult_206_n387) );
  OR2_X1 DP_mult_206_U1942 ( .A1(DP_mult_206_n1111), .A2(DP_mult_206_n1122), 
        .ZN(DP_mult_206_n2181) );
  OR2_X1 DP_mult_206_U1941 ( .A1(DP_mult_206_n1133), .A2(DP_mult_206_n1142), 
        .ZN(DP_mult_206_n2180) );
  NOR2_X1 DP_mult_206_U1940 ( .A1(DP_mult_206_n1085), .A2(DP_mult_206_n1098), 
        .ZN(DP_mult_206_n592) );
  NOR2_X1 DP_mult_206_U1939 ( .A1(DP_mult_206_n590), .A2(DP_mult_206_n592), 
        .ZN(DP_mult_206_n588) );
  AOI21_X1 DP_mult_206_U1938 ( .B1(DP_mult_206_n376), .B2(DP_mult_206_n2183), 
        .A(DP_mult_206_n367), .ZN(DP_mult_206_n365) );
  OAI21_X1 DP_mult_206_U1937 ( .B1(DP_mult_206_n364), .B2(DP_mult_206_n387), 
        .A(DP_mult_206_n365), .ZN(DP_mult_206_n363) );
  AOI21_X1 DP_mult_206_U1936 ( .B1(DP_mult_206_n362), .B2(DP_mult_206_n394), 
        .A(DP_mult_206_n363), .ZN(DP_mult_206_n361) );
  OAI21_X1 DP_mult_206_U1935 ( .B1(DP_mult_206_n405), .B2(DP_mult_206_n360), 
        .A(DP_mult_206_n361), .ZN(DP_mult_206_n359) );
  NAND2_X1 DP_mult_206_U1934 ( .A1(DP_mult_206_n2182), .A2(DP_mult_206_n2183), 
        .ZN(DP_mult_206_n364) );
  AOI21_X1 DP_mult_206_U1933 ( .B1(DP_mult_206_n2180), .B2(DP_mult_206_n1968), 
        .A(DP_mult_206_n1975), .ZN(DP_mult_206_n611) );
  OR2_X1 DP_mult_206_U1932 ( .A1(DP_mult_206_n1123), .A2(DP_mult_206_n1132), 
        .ZN(DP_mult_206_n2179) );
  OAI21_X1 DP_mult_206_U1931 ( .B1(DP_mult_206_n628), .B2(DP_mult_206_n626), 
        .A(DP_mult_206_n627), .ZN(DP_mult_206_n625) );
  AOI21_X1 DP_mult_206_U1930 ( .B1(DP_mult_206_n625), .B2(DP_mult_206_n1977), 
        .A(DP_mult_206_n1970), .ZN(DP_mult_206_n620) );
  OAI21_X1 DP_mult_206_U1929 ( .B1(DP_mult_206_n638), .B2(DP_mult_206_n636), 
        .A(DP_mult_206_n637), .ZN(DP_mult_206_n635) );
  AOI21_X1 DP_mult_206_U1928 ( .B1(DP_mult_206_n629), .B2(DP_mult_206_n635), 
        .A(DP_mult_206_n630), .ZN(DP_mult_206_n628) );
  OR2_X1 DP_mult_206_U1927 ( .A1(DP_mult_206_n709), .A2(DP_mult_206_n716), 
        .ZN(DP_mult_206_n2178) );
  OR2_X1 DP_mult_206_U1926 ( .A1(DP_mult_206_n717), .A2(DP_mult_206_n726), 
        .ZN(DP_mult_206_n2177) );
  NOR2_X1 DP_mult_206_U1925 ( .A1(DP_mult_206_n727), .A2(DP_mult_206_n736), 
        .ZN(DP_mult_206_n428) );
  OR2_X1 DP_mult_206_U1924 ( .A1(DP_mult_206_n701), .A2(DP_mult_206_n708), 
        .ZN(DP_mult_206_n2176) );
  INV_X1 DP_mult_206_U1923 ( .A(DP_mult_206_n352), .ZN(DP_mult_206_n350) );
  AOI21_X1 DP_mult_206_U1922 ( .B1(DP_mult_206_n359), .B2(DP_mult_206_n2184), 
        .A(DP_mult_206_n350), .ZN(DP_mult_206_n348) );
  NOR2_X1 DP_mult_206_U1921 ( .A1(DP_mult_206_n695), .A2(DP_mult_206_n700), 
        .ZN(DP_mult_206_n384) );
  NOR2_X1 DP_mult_206_U1920 ( .A1(DP_mult_206_n1099), .A2(DP_mult_206_n1110), 
        .ZN(DP_mult_206_n597) );
  NAND2_X1 DP_mult_206_U1919 ( .A1(DP_mult_206_n2176), .A2(DP_mult_206_n396), 
        .ZN(DP_mult_206_n307) );
  NAND2_X1 DP_mult_206_U1918 ( .A1(DP_mult_206_n661), .A2(DP_mult_206_n429), 
        .ZN(DP_mult_206_n310) );
  NAND2_X1 DP_mult_206_U1917 ( .A1(DP_mult_206_n2178), .A2(DP_mult_206_n409), 
        .ZN(DP_mult_206_n308) );
  OR2_X1 DP_mult_206_U1916 ( .A1(DP_mult_206_n1039), .A2(DP_mult_206_n1054), 
        .ZN(DP_mult_206_n2174) );
  NAND2_X1 DP_mult_206_U1915 ( .A1(DP_mult_206_n1003), .A2(DP_mult_206_n1020), 
        .ZN(DP_mult_206_n570) );
  INV_X1 DP_mult_206_U1914 ( .A(DP_mult_206_n384), .ZN(DP_mult_206_n657) );
  NAND2_X1 DP_mult_206_U1913 ( .A1(DP_mult_206_n657), .A2(DP_mult_206_n387), 
        .ZN(DP_mult_206_n306) );
  NAND2_X1 DP_mult_206_U1912 ( .A1(DP_mult_206_n400), .A2(DP_mult_206_n2176), 
        .ZN(DP_mult_206_n389) );
  NAND2_X1 DP_mult_206_U1911 ( .A1(DP_mult_206_n983), .A2(DP_mult_206_n1002), 
        .ZN(DP_mult_206_n564) );
  NOR2_X1 DP_mult_206_U1910 ( .A1(DP_mult_206_n389), .A2(DP_mult_206_n384), 
        .ZN(DP_mult_206_n382) );
  NAND2_X1 DP_mult_206_U1909 ( .A1(DP_mult_206_n963), .A2(DP_mult_206_n982), 
        .ZN(DP_mult_206_n559) );
  INV_X1 DP_mult_206_U1908 ( .A(DP_mult_206_n378), .ZN(DP_mult_206_n376) );
  INV_X1 DP_mult_206_U1907 ( .A(DP_mult_206_n396), .ZN(DP_mult_206_n394) );
  NAND2_X1 DP_mult_206_U1906 ( .A1(DP_mult_206_n362), .A2(DP_mult_206_n2176), 
        .ZN(DP_mult_206_n360) );
  NOR2_X1 DP_mult_206_U1905 ( .A1(DP_mult_206_n1003), .A2(DP_mult_206_n1020), 
        .ZN(DP_mult_206_n569) );
  OR2_X1 DP_mult_206_U1904 ( .A1(DP_mult_206_n761), .A2(DP_mult_206_n774), 
        .ZN(DP_mult_206_n2173) );
  OR2_X1 DP_mult_206_U1903 ( .A1(DP_mult_206_n1021), .A2(DP_mult_206_n1038), 
        .ZN(DP_mult_206_n2172) );
  NOR2_X1 DP_mult_206_U1902 ( .A1(DP_mult_206_n420), .A2(DP_mult_206_n347), 
        .ZN(DP_mult_206_n345) );
  NAND2_X1 DP_mult_206_U1901 ( .A1(DP_mult_206_n877), .A2(DP_mult_206_n896), 
        .ZN(DP_mult_206_n532) );
  NOR2_X1 DP_mult_206_U1900 ( .A1(DP_mult_206_n983), .A2(DP_mult_206_n1002), 
        .ZN(DP_mult_206_n563) );
  NAND2_X1 DP_mult_206_U1899 ( .A1(DP_mult_206_n737), .A2(DP_mult_206_n748), 
        .ZN(DP_mult_206_n436) );
  NAND2_X1 DP_mult_206_U1898 ( .A1(DP_mult_206_n821), .A2(DP_mult_206_n838), 
        .ZN(DP_mult_206_n503) );
  NAND2_X1 DP_mult_206_U1897 ( .A1(DP_mult_206_n857), .A2(DP_mult_206_n876), 
        .ZN(DP_mult_206_n521) );
  NOR2_X1 DP_mult_206_U1896 ( .A1(DP_mult_206_n857), .A2(DP_mult_206_n876), 
        .ZN(DP_mult_206_n520) );
  NAND2_X1 DP_mult_206_U1895 ( .A1(DP_mult_206_n789), .A2(DP_mult_206_n804), 
        .ZN(DP_mult_206_n481) );
  NOR2_X1 DP_mult_206_U1894 ( .A1(DP_mult_206_n384), .A2(DP_mult_206_n364), 
        .ZN(DP_mult_206_n362) );
  OAI21_X1 DP_mult_206_U1893 ( .B1(DP_mult_206_n620), .B2(DP_mult_206_n610), 
        .A(DP_mult_206_n611), .ZN(DP_mult_206_n609) );
  OAI21_X1 DP_mult_206_U1892 ( .B1(DP_mult_206_n600), .B2(DP_mult_206_n597), 
        .A(DP_mult_206_n598), .ZN(DP_mult_206_n596) );
  NOR2_X1 DP_mult_206_U1891 ( .A1(DP_mult_206_n597), .A2(DP_mult_206_n599), 
        .ZN(DP_mult_206_n595) );
  OAI21_X1 DP_mult_206_U1890 ( .B1(DP_mult_206_n590), .B2(DP_mult_206_n593), 
        .A(DP_mult_206_n591), .ZN(DP_mult_206_n589) );
  NOR2_X1 DP_mult_206_U1889 ( .A1(DP_mult_206_n435), .A2(DP_mult_206_n428), 
        .ZN(DP_mult_206_n426) );
  NAND2_X1 DP_mult_206_U1888 ( .A1(DP_mult_206_n2177), .A2(DP_mult_206_n2178), 
        .ZN(DP_mult_206_n402) );
  INV_X1 DP_mult_206_U1887 ( .A(DP_mult_206_n409), .ZN(DP_mult_206_n407) );
  AOI21_X1 DP_mult_206_U1886 ( .B1(DP_mult_206_n2178), .B2(DP_mult_206_n416), 
        .A(DP_mult_206_n407), .ZN(DP_mult_206_n405) );
  AOI21_X1 DP_mult_206_U1885 ( .B1(DP_mult_206_n426), .B2(DP_mult_206_n445), 
        .A(DP_mult_206_n427), .ZN(DP_mult_206_n421) );
  NOR2_X1 DP_mult_206_U1884 ( .A1(DP_mult_206_n1071), .A2(DP_mult_206_n1084), 
        .ZN(DP_mult_206_n590) );
  NAND2_X1 DP_mult_206_U1883 ( .A1(DP_mult_206_n662), .A2(DP_mult_206_n436), 
        .ZN(DP_mult_206_n311) );
  INV_X1 DP_mult_206_U1882 ( .A(DP_mult_206_n564), .ZN(DP_mult_206_n562) );
  INV_X1 DP_mult_206_U1881 ( .A(DP_mult_206_n563), .ZN(DP_mult_206_n561) );
  INV_X1 DP_mult_206_U1880 ( .A(DP_mult_206_n2123), .ZN(DP_mult_206_n670) );
  NOR2_X1 DP_mult_206_U1879 ( .A1(DP_mult_206_n402), .A2(DP_mult_206_n360), 
        .ZN(DP_mult_206_n356) );
  INV_X1 DP_mult_206_U1878 ( .A(DP_mult_206_n438), .ZN(DP_mult_206_n663) );
  INV_X1 DP_mult_206_U1877 ( .A(DP_mult_206_n461), .ZN(DP_mult_206_n459) );
  AOI21_X1 DP_mult_206_U1876 ( .B1(DP_mult_206_n2173), .B2(DP_mult_206_n472), 
        .A(DP_mult_206_n459), .ZN(DP_mult_206_n457) );
  NOR2_X1 DP_mult_206_U1875 ( .A1(DP_mult_206_n420), .A2(DP_mult_206_n402), 
        .ZN(DP_mult_206_n400) );
  INV_X1 DP_mult_206_U1874 ( .A(DP_mult_206_n521), .ZN(DP_mult_206_n519) );
  INV_X1 DP_mult_206_U1873 ( .A(DP_mult_206_n503), .ZN(DP_mult_206_n501) );
  INV_X1 DP_mult_206_U1872 ( .A(DP_mult_206_n481), .ZN(DP_mult_206_n483) );
  INV_X1 DP_mult_206_U1871 ( .A(DP_mult_206_n383), .ZN(DP_mult_206_n381) );
  INV_X1 DP_mult_206_U1870 ( .A(DP_mult_206_n436), .ZN(DP_mult_206_n434) );
  AOI21_X1 DP_mult_206_U1869 ( .B1(DP_mult_206_n662), .B2(DP_mult_206_n445), 
        .A(DP_mult_206_n434), .ZN(DP_mult_206_n432) );
  NAND2_X1 DP_mult_206_U1868 ( .A1(DP_mult_206_n663), .A2(DP_mult_206_n662), 
        .ZN(DP_mult_206_n431) );
  NAND2_X1 DP_mult_206_U1867 ( .A1(DP_mult_206_n426), .A2(DP_mult_206_n663), 
        .ZN(DP_mult_206_n420) );
  INV_X1 DP_mult_206_U1866 ( .A(DP_mult_206_n435), .ZN(DP_mult_206_n662) );
  NOR2_X1 DP_mult_206_U1865 ( .A1(DP_mult_206_n558), .A2(DP_mult_206_n563), 
        .ZN(DP_mult_206_n552) );
  INV_X1 DP_mult_206_U1864 ( .A(DP_mult_206_n420), .ZN(DP_mult_206_n422) );
  NOR2_X1 DP_mult_206_U1863 ( .A1(DP_mult_206_n491), .A2(DP_mult_206_n467), 
        .ZN(DP_mult_206_n465) );
  INV_X1 DP_mult_206_U1862 ( .A(DP_mult_206_n400), .ZN(DP_mult_206_n398) );
  INV_X1 DP_mult_206_U1861 ( .A(DP_mult_206_n505), .ZN(DP_mult_206_n507) );
  INV_X2 DP_mult_206_U1860 ( .A(DP_mult_206_n2290), .ZN(DP_mult_206_n2288) );
  INV_X2 DP_mult_206_U1859 ( .A(DP_mult_206_n2300), .ZN(DP_mult_206_n2298) );
  INV_X2 DP_mult_206_U1858 ( .A(DP_mult_206_n2305), .ZN(DP_mult_206_n2303) );
  INV_X2 DP_mult_206_U1857 ( .A(DP_mult_206_n2313), .ZN(DP_mult_206_n2311) );
  INV_X2 DP_mult_206_U1856 ( .A(DP_mult_206_n2310), .ZN(DP_mult_206_n2308) );
  INV_X2 DP_mult_206_U1855 ( .A(DP_mult_206_n2189), .ZN(DP_mult_206_n2242) );
  OR2_X1 DP_mult_206_U1854 ( .A1(DP_mult_206_n1143), .A2(DP_mult_206_n1150), 
        .ZN(DP_mult_206_n2170) );
  AND2_X2 DP_mult_206_U1853 ( .A1(DP_mult_206_n1809), .A2(DP_mult_206_n2251), 
        .ZN(DP_mult_206_n2195) );
  INV_X1 DP_mult_206_U1852 ( .A(DP_mult_206_n2195), .ZN(DP_mult_206_n2225) );
  AND2_X2 DP_mult_206_U1851 ( .A1(DP_mult_206_n1816), .A2(DP_mult_206_n253), 
        .ZN(DP_mult_206_n2197) );
  INV_X1 DP_mult_206_U1850 ( .A(DP_mult_206_n2125), .ZN(DP_mult_206_n2167) );
  INV_X2 DP_mult_206_U1849 ( .A(DP_mult_206_n537), .ZN(DP_mult_206_n536) );
  NAND3_X1 DP_mult_206_U1848 ( .A1(DP_mult_206_n2164), .A2(DP_mult_206_n2165), 
        .A3(DP_mult_206_n2166), .ZN(DP_mult_206_n842) );
  NAND2_X1 DP_mult_206_U1847 ( .A1(DP_mult_206_n849), .A2(DP_mult_206_n864), 
        .ZN(DP_mult_206_n2166) );
  NAND2_X1 DP_mult_206_U1846 ( .A1(DP_mult_206_n2053), .A2(DP_mult_206_n864), 
        .ZN(DP_mult_206_n2165) );
  NAND2_X1 DP_mult_206_U1845 ( .A1(DP_mult_206_n2053), .A2(DP_mult_206_n849), 
        .ZN(DP_mult_206_n2164) );
  XOR2_X1 DP_mult_206_U1844 ( .A(DP_mult_206_n2054), .B(DP_mult_206_n2163), 
        .Z(DP_mult_206_n843) );
  XOR2_X1 DP_mult_206_U1843 ( .A(DP_mult_206_n849), .B(DP_mult_206_n864), .Z(
        DP_mult_206_n2163) );
  INV_X1 DP_mult_206_U1842 ( .A(DP_mult_206_n2018), .ZN(DP_mult_206_n2255) );
  AND2_X2 DP_mult_206_U1841 ( .A1(DP_mult_206_n1810), .A2(DP_mult_206_n2254), 
        .ZN(DP_mult_206_n2196) );
  AND2_X2 DP_mult_206_U1840 ( .A1(DP_mult_206_n1815), .A2(DP_mult_206_n2262), 
        .ZN(DP_mult_206_n2194) );
  AND2_X2 DP_mult_206_U1839 ( .A1(DP_mult_206_n1811), .A2(DP_mult_206_n1932), 
        .ZN(DP_mult_206_n2199) );
  INV_X1 DP_mult_206_U1838 ( .A(DP_mult_206_n2194), .ZN(DP_mult_206_n2238) );
  NAND2_X1 DP_mult_206_U1837 ( .A1(DP_mult_206_n2161), .A2(DP_mult_206_n2162), 
        .ZN(DP_mult_206_n1416) );
  OR2_X1 DP_mult_206_U1836 ( .A1(DP_mult_206_n1713), .A2(DP_mult_206_n2263), 
        .ZN(DP_mult_206_n2162) );
  OR2_X1 DP_mult_206_U1835 ( .A1(DP_mult_206_n2238), .A2(DP_mult_206_n1714), 
        .ZN(DP_mult_206_n2161) );
  INV_X1 DP_mult_206_U1834 ( .A(DP_mult_206_n2194), .ZN(DP_mult_206_n2159) );
  NOR2_X1 DP_mult_206_U1833 ( .A1(DP_mult_206_n805), .A2(DP_mult_206_n820), 
        .ZN(DP_mult_206_n2158) );
  NAND2_X1 DP_mult_206_U1832 ( .A1(DP_mult_206_n873), .A2(DP_mult_206_n888), 
        .ZN(DP_mult_206_n2157) );
  NAND2_X1 DP_mult_206_U1831 ( .A1(DP_mult_206_n886), .A2(DP_mult_206_n888), 
        .ZN(DP_mult_206_n2156) );
  NAND2_X1 DP_mult_206_U1830 ( .A1(DP_mult_206_n886), .A2(DP_mult_206_n873), 
        .ZN(DP_mult_206_n2155) );
  OAI21_X1 DP_mult_206_U1829 ( .B1(DP_mult_206_n1945), .B2(DP_mult_206_n538), 
        .A(DP_mult_206_n2117), .ZN(DP_mult_206_n2153) );
  NAND3_X1 DP_mult_206_U1828 ( .A1(DP_mult_206_n2150), .A2(DP_mult_206_n2151), 
        .A3(DP_mult_206_n2152), .ZN(DP_mult_206_n918) );
  NAND2_X1 DP_mult_206_U1827 ( .A1(DP_mult_206_n942), .A2(DP_mult_206_n923), 
        .ZN(DP_mult_206_n2152) );
  NAND2_X1 DP_mult_206_U1826 ( .A1(DP_mult_206_n921), .A2(DP_mult_206_n923), 
        .ZN(DP_mult_206_n2151) );
  NAND2_X1 DP_mult_206_U1825 ( .A1(DP_mult_206_n921), .A2(DP_mult_206_n942), 
        .ZN(DP_mult_206_n2150) );
  INV_X1 DP_mult_206_U1824 ( .A(DP_mult_206_n2119), .ZN(DP_mult_206_n2221) );
  NAND3_X1 DP_mult_206_U1823 ( .A1(DP_mult_206_n2147), .A2(DP_mult_206_n2148), 
        .A3(DP_mult_206_n2149), .ZN(DP_mult_206_n884) );
  NAND2_X1 DP_mult_206_U1822 ( .A1(DP_mult_206_n891), .A2(DP_mult_206_n895), 
        .ZN(DP_mult_206_n2149) );
  NAND2_X1 DP_mult_206_U1821 ( .A1(DP_mult_206_n908), .A2(DP_mult_206_n895), 
        .ZN(DP_mult_206_n2148) );
  NAND2_X1 DP_mult_206_U1820 ( .A1(DP_mult_206_n908), .A2(DP_mult_206_n891), 
        .ZN(DP_mult_206_n2147) );
  XOR2_X1 DP_mult_206_U1819 ( .A(DP_mult_206_n908), .B(DP_mult_206_n2146), .Z(
        DP_mult_206_n885) );
  XOR2_X1 DP_mult_206_U1818 ( .A(DP_mult_206_n891), .B(DP_mult_206_n895), .Z(
        DP_mult_206_n2146) );
  INV_X1 DP_mult_206_U1817 ( .A(DP_mult_206_n2080), .ZN(DP_mult_206_n2262) );
  INV_X2 DP_mult_206_U1816 ( .A(DP_mult_206_n2280), .ZN(DP_mult_206_n2277) );
  INV_X1 DP_mult_206_U1815 ( .A(DP_mult_206_n1929), .ZN(DP_mult_206_n2248) );
  INV_X1 DP_mult_206_U1814 ( .A(DP_mult_206_n2089), .ZN(DP_mult_206_n2251) );
  INV_X1 DP_mult_206_U1813 ( .A(DP_mult_206_n2120), .ZN(DP_mult_206_n2245) );
  INV_X2 DP_mult_206_U1812 ( .A(DP_mult_206_n2290), .ZN(DP_mult_206_n2287) );
  INV_X1 DP_mult_206_U1811 ( .A(DP_coeffs_ff_int[0]), .ZN(DP_mult_206_n2326)
         );
  INV_X2 DP_mult_206_U1810 ( .A(DP_mult_206_n2310), .ZN(DP_mult_206_n2307) );
  XNOR2_X1 DP_mult_206_U1809 ( .A(DP_mult_206_n942), .B(DP_mult_206_n923), 
        .ZN(DP_mult_206_n2145) );
  XNOR2_X1 DP_mult_206_U1808 ( .A(DP_mult_206_n2145), .B(DP_mult_206_n921), 
        .ZN(DP_mult_206_n919) );
  INV_X1 DP_mult_206_U1807 ( .A(DP_mult_206_n2006), .ZN(DP_mult_206_n2236) );
  NOR2_X1 DP_mult_206_U1806 ( .A1(DP_mult_206_n856), .A2(DP_mult_206_n839), 
        .ZN(DP_mult_206_n513) );
  NOR2_X1 DP_mult_206_U1805 ( .A1(DP_mult_206_n839), .A2(DP_mult_206_n856), 
        .ZN(DP_mult_206_n2144) );
  INV_X1 DP_mult_206_U1804 ( .A(DP_mult_206_n2154), .ZN(DP_mult_206_n2254) );
  NAND3_X1 DP_mult_206_U1803 ( .A1(DP_mult_206_n2141), .A2(DP_mult_206_n2142), 
        .A3(DP_mult_206_n2143), .ZN(DP_mult_206_n972) );
  NAND2_X1 DP_mult_206_U1802 ( .A1(DP_mult_206_n1217), .A2(DP_mult_206_n994), 
        .ZN(DP_mult_206_n2143) );
  NAND2_X1 DP_mult_206_U1801 ( .A1(DP_mult_206_n996), .A2(DP_mult_206_n994), 
        .ZN(DP_mult_206_n2142) );
  NAND2_X1 DP_mult_206_U1800 ( .A1(DP_mult_206_n996), .A2(DP_mult_206_n1217), 
        .ZN(DP_mult_206_n2141) );
  NAND2_X1 DP_mult_206_U1799 ( .A1(DP_mult_206_n1416), .A2(DP_mult_206_n1328), 
        .ZN(DP_mult_206_n2140) );
  NAND2_X1 DP_mult_206_U1798 ( .A1(DP_mult_206_n1306), .A2(DP_mult_206_n1328), 
        .ZN(DP_mult_206_n2139) );
  NAND2_X1 DP_mult_206_U1797 ( .A1(DP_mult_206_n2091), .A2(DP_mult_206_n1306), 
        .ZN(DP_mult_206_n2138) );
  AND2_X1 DP_mult_206_U1796 ( .A1(DP_mult_206_n1806), .A2(DP_mult_206_n2243), 
        .ZN(DP_mult_206_n2136) );
  INV_X1 DP_mult_206_U1795 ( .A(DP_mult_206_n2005), .ZN(DP_mult_206_n2134) );
  INV_X1 DP_mult_206_U1794 ( .A(DP_mult_206_n2006), .ZN(DP_mult_206_n2135) );
  INV_X2 DP_mult_206_U1793 ( .A(DP_mult_206_n2192), .ZN(DP_mult_206_n2259) );
  INV_X2 DP_mult_206_U1792 ( .A(DP_mult_206_n2322), .ZN(DP_mult_206_n2319) );
  AND2_X2 DP_mult_206_U1791 ( .A1(DP_mult_206_n2171), .A2(DP_mult_206_n2036), 
        .ZN(DP_mult_206_n2193) );
  INV_X2 DP_mult_206_U1790 ( .A(DP_mult_206_n2193), .ZN(DP_mult_206_n2233) );
  INV_X1 DP_mult_206_U1789 ( .A(DP_mult_206_n2198), .ZN(DP_mult_206_n2223) );
  CLKBUF_X1 DP_mult_206_U1788 ( .A(DP_mult_206_n512), .Z(DP_mult_206_n2131) );
  INV_X1 DP_mult_206_U1787 ( .A(DP_mult_206_n2198), .ZN(DP_mult_206_n2130) );
  CLKBUF_X1 DP_mult_206_U1786 ( .A(DP_mult_206_n1260), .Z(DP_mult_206_n2128)
         );
  OR2_X1 DP_mult_206_U1785 ( .A1(DP_mult_206_n897), .A2(DP_mult_206_n918), 
        .ZN(DP_mult_206_n2125) );
  INV_X2 DP_mult_206_U1784 ( .A(DP_mult_206_n2285), .ZN(DP_mult_206_n2282) );
  CLKBUF_X1 DP_mult_206_U1783 ( .A(DP_mult_206_n511), .Z(DP_mult_206_n2124) );
  CLKBUF_X1 DP_mult_206_U1782 ( .A(DP_mult_206_n520), .Z(DP_mult_206_n2123) );
  INV_X1 DP_mult_206_U1781 ( .A(DP_mult_206_n2200), .ZN(DP_mult_206_n2122) );
  INV_X1 DP_mult_206_U1780 ( .A(DP_mult_206_n2197), .ZN(DP_mult_206_n2240) );
  CLKBUF_X1 DP_mult_206_U1779 ( .A(DP_mult_206_n2058), .Z(DP_mult_206_n2118)
         );
  AOI21_X1 DP_mult_206_U1778 ( .B1(DP_mult_206_n553), .B2(DP_mult_206_n540), 
        .A(DP_mult_206_n541), .ZN(DP_mult_206_n2117) );
  NOR2_X2 DP_mult_206_U1777 ( .A1(DP_mult_206_n502), .A2(DP_mult_206_n495), 
        .ZN(DP_mult_206_n489) );
  INV_X2 DP_mult_206_U1776 ( .A(DP_mult_206_n2276), .ZN(DP_mult_206_n2272) );
  INV_X1 DP_mult_206_U1775 ( .A(DP_mult_206_n2275), .ZN(DP_mult_206_n2271) );
  NAND3_X1 DP_mult_206_U1774 ( .A1(DP_mult_206_n2114), .A2(DP_mult_206_n2115), 
        .A3(DP_mult_206_n2116), .ZN(DP_mult_206_n992) );
  NAND2_X1 DP_mult_206_U1773 ( .A1(DP_mult_206_n1394), .A2(DP_mult_206_n1018), 
        .ZN(DP_mult_206_n2116) );
  NAND2_X1 DP_mult_206_U1772 ( .A1(DP_mult_206_n1001), .A2(DP_mult_206_n1018), 
        .ZN(DP_mult_206_n2115) );
  NAND2_X1 DP_mult_206_U1771 ( .A1(DP_mult_206_n1001), .A2(DP_mult_206_n1394), 
        .ZN(DP_mult_206_n2114) );
  NAND3_X1 DP_mult_206_U1770 ( .A1(DP_mult_206_n2111), .A2(DP_mult_206_n2112), 
        .A3(DP_mult_206_n2113), .ZN(DP_mult_206_n1018) );
  NAND2_X1 DP_mult_206_U1769 ( .A1(DP_mult_206_n1351), .A2(DP_mult_206_n1285), 
        .ZN(DP_mult_206_n2113) );
  NAND2_X1 DP_mult_206_U1768 ( .A1(DP_mult_206_n1263), .A2(DP_mult_206_n1285), 
        .ZN(DP_mult_206_n2112) );
  NAND2_X1 DP_mult_206_U1767 ( .A1(DP_mult_206_n1263), .A2(DP_mult_206_n1351), 
        .ZN(DP_mult_206_n2111) );
  XOR2_X1 DP_mult_206_U1766 ( .A(DP_mult_206_n2110), .B(DP_mult_206_n1285), 
        .Z(DP_mult_206_n1019) );
  XOR2_X1 DP_mult_206_U1765 ( .A(DP_mult_206_n1263), .B(DP_mult_206_n1351), 
        .Z(DP_mult_206_n2110) );
  NOR2_X1 DP_mult_206_U1764 ( .A1(DP_mult_206_n896), .A2(DP_mult_206_n877), 
        .ZN(DP_mult_206_n531) );
  NOR2_X1 DP_mult_206_U1763 ( .A1(DP_mult_206_n877), .A2(DP_mult_206_n896), 
        .ZN(DP_mult_206_n2109) );
  INV_X1 DP_mult_206_U1762 ( .A(DP_mult_206_n2253), .ZN(DP_mult_206_n2108) );
  NAND3_X1 DP_mult_206_U1761 ( .A1(DP_mult_206_n2105), .A2(DP_mult_206_n2106), 
        .A3(DP_mult_206_n2107), .ZN(DP_mult_206_n796) );
  NAND2_X1 DP_mult_206_U1760 ( .A1(DP_mult_206_n1274), .A2(DP_mult_206_n1296), 
        .ZN(DP_mult_206_n2107) );
  NAND2_X1 DP_mult_206_U1759 ( .A1(DP_mult_206_n818), .A2(DP_mult_206_n1296), 
        .ZN(DP_mult_206_n2106) );
  NAND2_X1 DP_mult_206_U1758 ( .A1(DP_mult_206_n818), .A2(DP_mult_206_n1274), 
        .ZN(DP_mult_206_n2105) );
  NAND3_X1 DP_mult_206_U1757 ( .A1(DP_mult_206_n2101), .A2(DP_mult_206_n2102), 
        .A3(DP_mult_206_n2103), .ZN(DP_mult_206_n928) );
  NAND2_X1 DP_mult_206_U1756 ( .A1(DP_mult_206_n956), .A2(DP_mult_206_n954), 
        .ZN(DP_mult_206_n2103) );
  NAND2_X1 DP_mult_206_U1755 ( .A1(DP_mult_206_n2032), .A2(DP_mult_206_n954), 
        .ZN(DP_mult_206_n2102) );
  NAND2_X1 DP_mult_206_U1754 ( .A1(DP_mult_206_n2032), .A2(DP_mult_206_n956), 
        .ZN(DP_mult_206_n2101) );
  XOR2_X1 DP_mult_206_U1753 ( .A(DP_mult_206_n2100), .B(DP_mult_206_n954), .Z(
        DP_mult_206_n929) );
  XOR2_X1 DP_mult_206_U1752 ( .A(DP_mult_206_n2032), .B(DP_mult_206_n1940), 
        .Z(DP_mult_206_n2100) );
  NAND2_X1 DP_mult_206_U1751 ( .A1(DP_mult_206_n1414), .A2(DP_mult_206_n1282), 
        .ZN(DP_mult_206_n2099) );
  NAND2_X1 DP_mult_206_U1750 ( .A1(DP_mult_206_n1304), .A2(DP_mult_206_n1282), 
        .ZN(DP_mult_206_n2098) );
  NAND2_X1 DP_mult_206_U1749 ( .A1(DP_mult_206_n1304), .A2(DP_mult_206_n1414), 
        .ZN(DP_mult_206_n2097) );
  XOR2_X1 DP_mult_206_U1748 ( .A(DP_mult_206_n2096), .B(DP_mult_206_n1282), 
        .Z(DP_mult_206_n955) );
  XOR2_X1 DP_mult_206_U1747 ( .A(DP_mult_206_n1304), .B(DP_mult_206_n1414), 
        .Z(DP_mult_206_n2096) );
  INV_X2 DP_mult_206_U1746 ( .A(DP_mult_206_n2306), .ZN(DP_mult_206_n2302) );
  NAND3_X1 DP_mult_206_U1745 ( .A1(DP_mult_206_n2093), .A2(DP_mult_206_n2094), 
        .A3(DP_mult_206_n2095), .ZN(DP_mult_206_n848) );
  NAND2_X1 DP_mult_206_U1744 ( .A1(DP_mult_206_n1365), .A2(DP_mult_206_n1410), 
        .ZN(DP_mult_206_n2095) );
  NAND2_X1 DP_mult_206_U1743 ( .A1(DP_mult_206_n872), .A2(DP_mult_206_n1410), 
        .ZN(DP_mult_206_n2094) );
  NAND2_X1 DP_mult_206_U1742 ( .A1(DP_mult_206_n872), .A2(DP_mult_206_n1365), 
        .ZN(DP_mult_206_n2093) );
  XOR2_X1 DP_mult_206_U1741 ( .A(DP_mult_206_n872), .B(DP_mult_206_n2092), .Z(
        DP_mult_206_n849) );
  XOR2_X1 DP_mult_206_U1740 ( .A(DP_mult_206_n1365), .B(DP_mult_206_n1410), 
        .Z(DP_mult_206_n2092) );
  NAND2_X1 DP_mult_206_U1739 ( .A1(DP_mult_206_n2161), .A2(DP_mult_206_n2162), 
        .ZN(DP_mult_206_n2091) );
  CLKBUF_X1 DP_mult_206_U1738 ( .A(DP_mult_206_n505), .Z(DP_mult_206_n2090) );
  INV_X1 DP_mult_206_U1737 ( .A(DP_mult_206_n1929), .ZN(DP_mult_206_n2250) );
  XOR2_X1 DP_mult_206_U1736 ( .A(DP_coeffs_ff_int[9]), .B(DP_coeffs_ff_int[10]), .Z(DP_mult_206_n2154) );
  INV_X1 DP_mult_206_U1735 ( .A(DP_mult_206_n2018), .ZN(DP_mult_206_n2256) );
  AND2_X1 DP_mult_206_U1734 ( .A1(DP_mult_206_n1807), .A2(DP_mult_206_n2245), 
        .ZN(DP_mult_206_n2119) );
  NAND3_X1 DP_mult_206_U1733 ( .A1(DP_mult_206_n2086), .A2(DP_mult_206_n2087), 
        .A3(DP_mult_206_n2088), .ZN(DP_mult_206_n824) );
  NAND2_X1 DP_mult_206_U1732 ( .A1(DP_mult_206_n829), .A2(DP_mult_206_n846), 
        .ZN(DP_mult_206_n2088) );
  NAND2_X1 DP_mult_206_U1731 ( .A1(DP_mult_206_n848), .A2(DP_mult_206_n846), 
        .ZN(DP_mult_206_n2087) );
  NAND2_X1 DP_mult_206_U1730 ( .A1(DP_mult_206_n848), .A2(DP_mult_206_n829), 
        .ZN(DP_mult_206_n2086) );
  XOR2_X1 DP_mult_206_U1729 ( .A(DP_mult_206_n2085), .B(DP_mult_206_n846), .Z(
        DP_mult_206_n825) );
  XOR2_X1 DP_mult_206_U1728 ( .A(DP_mult_206_n848), .B(DP_mult_206_n829), .Z(
        DP_mult_206_n2085) );
  NAND3_X1 DP_mult_206_U1727 ( .A1(DP_mult_206_n2082), .A2(DP_mult_206_n2083), 
        .A3(DP_mult_206_n2084), .ZN(DP_mult_206_n846) );
  NAND2_X1 DP_mult_206_U1726 ( .A1(DP_mult_206_n870), .A2(DP_mult_206_n851), 
        .ZN(DP_mult_206_n2084) );
  NAND2_X1 DP_mult_206_U1725 ( .A1(DP_mult_206_n868), .A2(DP_mult_206_n851), 
        .ZN(DP_mult_206_n2083) );
  NAND2_X1 DP_mult_206_U1724 ( .A1(DP_mult_206_n868), .A2(DP_mult_206_n870), 
        .ZN(DP_mult_206_n2082) );
  XOR2_X1 DP_mult_206_U1723 ( .A(DP_mult_206_n2081), .B(DP_mult_206_n851), .Z(
        DP_mult_206_n847) );
  XOR2_X1 DP_mult_206_U1722 ( .A(DP_mult_206_n868), .B(DP_mult_206_n870), .Z(
        DP_mult_206_n2081) );
  NAND3_X1 DP_mult_206_U1721 ( .A1(DP_mult_206_n2077), .A2(DP_mult_206_n2078), 
        .A3(DP_mult_206_n2079), .ZN(DP_mult_206_n1020) );
  NAND2_X1 DP_mult_206_U1720 ( .A1(DP_mult_206_n1025), .A2(DP_mult_206_n1023), 
        .ZN(DP_mult_206_n2079) );
  NAND2_X1 DP_mult_206_U1719 ( .A1(DP_mult_206_n1040), .A2(DP_mult_206_n1023), 
        .ZN(DP_mult_206_n2078) );
  NAND2_X1 DP_mult_206_U1718 ( .A1(DP_mult_206_n1040), .A2(DP_mult_206_n1025), 
        .ZN(DP_mult_206_n2077) );
  NAND3_X1 DP_mult_206_U1717 ( .A1(DP_mult_206_n2074), .A2(DP_mult_206_n2075), 
        .A3(DP_mult_206_n2076), .ZN(DP_mult_206_n1022) );
  NAND2_X1 DP_mult_206_U1716 ( .A1(DP_mult_206_n1044), .A2(DP_mult_206_n1042), 
        .ZN(DP_mult_206_n2076) );
  NAND2_X1 DP_mult_206_U1715 ( .A1(DP_mult_206_n1027), .A2(DP_mult_206_n1042), 
        .ZN(DP_mult_206_n2075) );
  NAND2_X1 DP_mult_206_U1714 ( .A1(DP_mult_206_n1027), .A2(DP_mult_206_n1044), 
        .ZN(DP_mult_206_n2074) );
  XOR2_X1 DP_mult_206_U1713 ( .A(DP_mult_206_n2073), .B(DP_mult_206_n1042), 
        .Z(DP_mult_206_n1023) );
  XOR2_X1 DP_mult_206_U1712 ( .A(DP_mult_206_n1027), .B(DP_mult_206_n1044), 
        .Z(DP_mult_206_n2073) );
  XNOR2_X1 DP_mult_206_U1711 ( .A(DP_coeffs_ff_int[3]), .B(DP_mult_206_n2322), 
        .ZN(DP_mult_206_n1807) );
  XNOR2_X1 DP_mult_206_U1710 ( .A(DP_mult_206_n1040), .B(DP_mult_206_n1025), 
        .ZN(DP_mult_206_n2072) );
  XNOR2_X1 DP_mult_206_U1709 ( .A(DP_mult_206_n2072), .B(DP_mult_206_n1023), 
        .ZN(DP_mult_206_n1021) );
  XNOR2_X1 DP_mult_206_U1708 ( .A(DP_mult_206_n2091), .B(DP_mult_206_n1306), 
        .ZN(DP_mult_206_n2071) );
  XNOR2_X1 DP_mult_206_U1707 ( .A(DP_mult_206_n2071), .B(DP_mult_206_n2003), 
        .ZN(DP_mult_206_n995) );
  NAND3_X1 DP_mult_206_U1706 ( .A1(DP_mult_206_n2068), .A2(DP_mult_206_n2069), 
        .A3(DP_mult_206_n2070), .ZN(DP_mult_206_n896) );
  NAND2_X1 DP_mult_206_U1705 ( .A1(DP_mult_206_n901), .A2(DP_mult_206_n899), 
        .ZN(DP_mult_206_n2070) );
  NAND2_X1 DP_mult_206_U1704 ( .A1(DP_mult_206_n920), .A2(DP_mult_206_n899), 
        .ZN(DP_mult_206_n2069) );
  NAND2_X1 DP_mult_206_U1703 ( .A1(DP_mult_206_n920), .A2(DP_mult_206_n901), 
        .ZN(DP_mult_206_n2068) );
  NAND3_X1 DP_mult_206_U1702 ( .A1(DP_mult_206_n2065), .A2(DP_mult_206_n2066), 
        .A3(DP_mult_206_n2067), .ZN(DP_mult_206_n898) );
  NAND2_X1 DP_mult_206_U1701 ( .A1(DP_mult_206_n922), .A2(DP_mult_206_n924), 
        .ZN(DP_mult_206_n2067) );
  NAND2_X1 DP_mult_206_U1700 ( .A1(DP_mult_206_n922), .A2(DP_mult_206_n903), 
        .ZN(DP_mult_206_n2066) );
  NAND2_X1 DP_mult_206_U1699 ( .A1(DP_mult_206_n903), .A2(DP_mult_206_n924), 
        .ZN(DP_mult_206_n2065) );
  XOR2_X1 DP_mult_206_U1698 ( .A(DP_mult_206_n922), .B(DP_mult_206_n2064), .Z(
        DP_mult_206_n899) );
  XOR2_X1 DP_mult_206_U1697 ( .A(DP_mult_206_n903), .B(DP_mult_206_n924), .Z(
        DP_mult_206_n2064) );
  INV_X2 DP_mult_206_U1696 ( .A(DP_mult_206_n2296), .ZN(DP_mult_206_n2293) );
  INV_X1 DP_mult_206_U1695 ( .A(DP_mult_206_n519), .ZN(DP_mult_206_n2063) );
  XNOR2_X1 DP_mult_206_U1694 ( .A(DP_coeffs_ff_int[17]), .B(
        DP_coeffs_ff_int[18]), .ZN(DP_mult_206_n2062) );
  XNOR2_X1 DP_mult_206_U1693 ( .A(DP_coeffs_ff_int[17]), .B(DP_mult_206_n2291), 
        .ZN(DP_mult_206_n1814) );
  AND2_X2 DP_mult_206_U1692 ( .A1(DP_mult_206_n1817), .A2(DP_mult_206_n2269), 
        .ZN(DP_mult_206_n2189) );
  INV_X2 DP_mult_206_U1691 ( .A(DP_mult_206_n2189), .ZN(DP_mult_206_n2241) );
  INV_X1 DP_mult_206_U1690 ( .A(DP_coeffs_ff_int[2]), .ZN(DP_mult_206_n2322)
         );
  INV_X1 DP_mult_206_U1689 ( .A(DP_mult_206_n2133), .ZN(DP_mult_206_n2192) );
  INV_X1 DP_mult_206_U1688 ( .A(DP_mult_206_n2199), .ZN(DP_mult_206_n2229) );
  INV_X1 DP_mult_206_U1687 ( .A(DP_mult_206_n2199), .ZN(DP_mult_206_n2061) );
  XNOR2_X1 DP_mult_206_U1686 ( .A(DP_mult_206_n996), .B(DP_mult_206_n1217), 
        .ZN(DP_mult_206_n2059) );
  XNOR2_X1 DP_mult_206_U1685 ( .A(DP_mult_206_n2059), .B(DP_mult_206_n994), 
        .ZN(DP_mult_206_n973) );
  INV_X1 DP_mult_206_U1684 ( .A(DP_mult_206_n2190), .ZN(DP_mult_206_n2243) );
  OAI21_X1 DP_mult_206_U1683 ( .B1(DP_mult_206_n1984), .B2(DP_mult_206_n564), 
        .A(DP_mult_206_n559), .ZN(DP_mult_206_n2058) );
  XNOR2_X1 DP_mult_206_U1682 ( .A(DP_mult_206_n920), .B(DP_mult_206_n901), 
        .ZN(DP_mult_206_n2057) );
  XNOR2_X1 DP_mult_206_U1681 ( .A(DP_mult_206_n2057), .B(DP_mult_206_n899), 
        .ZN(DP_mult_206_n897) );
  XNOR2_X1 DP_mult_206_U1680 ( .A(DP_coeffs_ff_int[13]), .B(
        DP_coeffs_ff_int[14]), .ZN(DP_mult_206_n2133) );
  NOR2_X1 DP_mult_206_U1679 ( .A1(DP_mult_206_n2109), .A2(DP_mult_206_n534), 
        .ZN(DP_mult_206_n525) );
  INV_X2 DP_mult_206_U1678 ( .A(DP_mult_206_n2192), .ZN(DP_mult_206_n2056) );
  NOR2_X1 DP_mult_206_U1677 ( .A1(DP_mult_206_n941), .A2(DP_mult_206_n962), 
        .ZN(DP_mult_206_n547) );
  INV_X1 DP_mult_206_U1676 ( .A(DP_mult_206_n674), .ZN(DP_mult_206_n2055) );
  NAND3_X1 DP_mult_206_U1675 ( .A1(DP_mult_206_n2155), .A2(DP_mult_206_n2156), 
        .A3(DP_mult_206_n2157), .ZN(DP_mult_206_n2053) );
  NAND3_X1 DP_mult_206_U1674 ( .A1(DP_mult_206_n2155), .A2(DP_mult_206_n2156), 
        .A3(DP_mult_206_n2157), .ZN(DP_mult_206_n2054) );
  NAND3_X1 DP_mult_206_U1673 ( .A1(DP_mult_206_n2164), .A2(DP_mult_206_n2165), 
        .A3(DP_mult_206_n2166), .ZN(DP_mult_206_n2052) );
  XNOR2_X1 DP_mult_206_U1672 ( .A(DP_mult_206_n873), .B(DP_mult_206_n888), 
        .ZN(DP_mult_206_n2051) );
  XNOR2_X1 DP_mult_206_U1671 ( .A(DP_mult_206_n1934), .B(DP_mult_206_n2051), 
        .ZN(DP_mult_206_n863) );
  XNOR2_X1 DP_mult_206_U1670 ( .A(DP_coeffs_ff_int[19]), .B(DP_mult_206_n2285), 
        .ZN(DP_mult_206_n1815) );
  OAI22_X1 DP_mult_206_U1669 ( .A1(DP_mult_206_n2239), .A2(DP_mult_206_n1733), 
        .B1(DP_mult_206_n1732), .B2(DP_mult_206_n2265), .ZN(DP_mult_206_n2050)
         );
  OR2_X1 DP_mult_206_U1668 ( .A1(DP_mult_206_n1992), .A2(DP_mult_206_n856), 
        .ZN(DP_mult_206_n2049) );
  INV_X1 DP_mult_206_U1667 ( .A(DP_mult_206_n2121), .ZN(DP_mult_206_n2246) );
  INV_X1 DP_mult_206_U1666 ( .A(DP_mult_206_n2121), .ZN(DP_mult_206_n2048) );
  NAND3_X1 DP_mult_206_U1665 ( .A1(DP_mult_206_n2045), .A2(DP_mult_206_n2046), 
        .A3(DP_mult_206_n2047), .ZN(DP_mult_206_n830) );
  NAND2_X1 DP_mult_206_U1664 ( .A1(DP_mult_206_n1298), .A2(DP_mult_206_n1320), 
        .ZN(DP_mult_206_n2047) );
  NAND2_X1 DP_mult_206_U1663 ( .A1(DP_mult_206_n1254), .A2(DP_mult_206_n1320), 
        .ZN(DP_mult_206_n2046) );
  NAND2_X1 DP_mult_206_U1662 ( .A1(DP_mult_206_n1254), .A2(DP_mult_206_n1298), 
        .ZN(DP_mult_206_n2045) );
  XOR2_X1 DP_mult_206_U1661 ( .A(DP_mult_206_n2044), .B(DP_mult_206_n2034), 
        .Z(DP_mult_206_n831) );
  XOR2_X1 DP_mult_206_U1660 ( .A(DP_mult_206_n1298), .B(DP_mult_206_n1320), 
        .Z(DP_mult_206_n2044) );
  INV_X2 DP_mult_206_U1659 ( .A(DP_mult_206_n2194), .ZN(DP_mult_206_n2160) );
  XNOR2_X1 DP_mult_206_U1658 ( .A(DP_coeffs_ff_int[1]), .B(DP_mult_206_n2326), 
        .ZN(DP_mult_206_n1806) );
  INV_X1 DP_mult_206_U1657 ( .A(DP_mult_206_n2062), .ZN(DP_mult_206_n2191) );
  NAND3_X1 DP_mult_206_U1656 ( .A1(DP_mult_206_n2041), .A2(DP_mult_206_n2042), 
        .A3(DP_mult_206_n2043), .ZN(DP_mult_206_n1038) );
  NAND2_X1 DP_mult_206_U1655 ( .A1(DP_mult_206_n1056), .A2(DP_mult_206_n1043), 
        .ZN(DP_mult_206_n2043) );
  NAND2_X1 DP_mult_206_U1654 ( .A1(DP_mult_206_n1041), .A2(DP_mult_206_n1043), 
        .ZN(DP_mult_206_n2042) );
  NAND2_X1 DP_mult_206_U1653 ( .A1(DP_mult_206_n1041), .A2(DP_mult_206_n1056), 
        .ZN(DP_mult_206_n2041) );
  XNOR2_X1 DP_mult_206_U1652 ( .A(DP_mult_206_n1274), .B(DP_mult_206_n1296), 
        .ZN(DP_mult_206_n2040) );
  XNOR2_X1 DP_mult_206_U1651 ( .A(DP_mult_206_n818), .B(DP_mult_206_n2040), 
        .ZN(DP_mult_206_n797) );
  XNOR2_X1 DP_mult_206_U1650 ( .A(DP_coeffs_ff_int[23]), .B(DP_mult_206_n2276), 
        .ZN(DP_mult_206_n1817) );
  INV_X2 DP_mult_206_U1649 ( .A(DP_mult_206_n2191), .ZN(DP_mult_206_n2039) );
  INV_X1 DP_mult_206_U1648 ( .A(DP_mult_206_n2198), .ZN(DP_mult_206_n2129) );
  INV_X2 DP_mult_206_U1647 ( .A(DP_mult_206_n2037), .ZN(DP_mult_206_n2038) );
  INV_X1 DP_mult_206_U1646 ( .A(DP_coeffs_ff_int[6]), .ZN(DP_mult_206_n2037)
         );
  INV_X2 DP_mult_206_U1645 ( .A(DP_mult_206_n2132), .ZN(DP_mult_206_n2260) );
  XNOR2_X1 DP_mult_206_U1644 ( .A(DP_coeffs_ff_int[16]), .B(
        DP_coeffs_ff_int[15]), .ZN(DP_mult_206_n2036) );
  XNOR2_X1 DP_mult_206_U1643 ( .A(DP_coeffs_ff_int[7]), .B(DP_mult_206_n2037), 
        .ZN(DP_mult_206_n1809) );
  BUF_X2 DP_mult_206_U1642 ( .A(DP_mult_206_n285), .Z(DP_mult_206_n2035) );
  INV_X2 DP_mult_206_U1641 ( .A(DP_mult_206_n2194), .ZN(DP_mult_206_n2237) );
  INV_X1 DP_mult_206_U1640 ( .A(DP_mult_206_n2080), .ZN(DP_mult_206_n2263) );
  XOR2_X1 DP_mult_206_U1639 ( .A(DP_coeffs_ff_int[7]), .B(DP_coeffs_ff_int[8]), 
        .Z(DP_mult_206_n2089) );
  INV_X1 DP_mult_206_U1638 ( .A(DP_mult_206_n1943), .ZN(DP_mult_206_n2033) );
  NAND3_X1 DP_mult_206_U1637 ( .A1(DP_mult_206_n2209), .A2(DP_mult_206_n2210), 
        .A3(DP_mult_206_n2211), .ZN(DP_mult_206_n2032) );
  INV_X2 DP_mult_206_U1636 ( .A(DP_mult_206_n2197), .ZN(DP_mult_206_n2031) );
  NAND2_X1 DP_mult_206_U1635 ( .A1(DP_mult_206_n2029), .A2(DP_mult_206_n2030), 
        .ZN(DP_mult_206_n836) );
  OR2_X1 DP_mult_206_U1634 ( .A1(DP_mult_206_n1682), .A2(DP_mult_206_n2261), 
        .ZN(DP_mult_206_n2030) );
  NAND3_X1 DP_mult_206_U1633 ( .A1(DP_mult_206_n2026), .A2(DP_mult_206_n2027), 
        .A3(DP_mult_206_n2028), .ZN(DP_mult_206_n834) );
  NAND2_X1 DP_mult_206_U1632 ( .A1(DP_mult_206_n1276), .A2(DP_mult_206_n1210), 
        .ZN(DP_mult_206_n2028) );
  NAND2_X1 DP_mult_206_U1631 ( .A1(DP_mult_206_n2004), .A2(DP_mult_206_n1210), 
        .ZN(DP_mult_206_n2027) );
  NAND2_X1 DP_mult_206_U1630 ( .A1(DP_mult_206_n2004), .A2(DP_mult_206_n1276), 
        .ZN(DP_mult_206_n2026) );
  XOR2_X1 DP_mult_206_U1629 ( .A(DP_mult_206_n2004), .B(DP_mult_206_n2025), 
        .Z(DP_mult_206_n835) );
  XOR2_X1 DP_mult_206_U1628 ( .A(DP_mult_206_n1276), .B(DP_mult_206_n1210), 
        .Z(DP_mult_206_n2025) );
  INV_X1 DP_mult_206_U1627 ( .A(DP_mult_206_n2196), .ZN(DP_mult_206_n2227) );
  NAND3_X1 DP_mult_206_U1626 ( .A1(DP_mult_206_n2021), .A2(DP_mult_206_n2022), 
        .A3(DP_mult_206_n2023), .ZN(DP_mult_206_n790) );
  NAND2_X1 DP_mult_206_U1625 ( .A1(DP_mult_206_n795), .A2(DP_mult_206_n810), 
        .ZN(DP_mult_206_n2023) );
  NAND2_X1 DP_mult_206_U1624 ( .A1(DP_mult_206_n808), .A2(DP_mult_206_n810), 
        .ZN(DP_mult_206_n2022) );
  NAND2_X1 DP_mult_206_U1623 ( .A1(DP_mult_206_n808), .A2(DP_mult_206_n795), 
        .ZN(DP_mult_206_n2021) );
  XOR2_X1 DP_mult_206_U1622 ( .A(DP_mult_206_n808), .B(DP_mult_206_n2020), .Z(
        DP_mult_206_n791) );
  XOR2_X1 DP_mult_206_U1621 ( .A(DP_mult_206_n795), .B(DP_mult_206_n810), .Z(
        DP_mult_206_n2020) );
  INV_X2 DP_mult_206_U1620 ( .A(DP_mult_206_n2291), .ZN(DP_mult_206_n2289) );
  XNOR2_X1 DP_mult_206_U1619 ( .A(DP_coeffs_ff_int[15]), .B(DP_mult_206_n2295), 
        .ZN(DP_mult_206_n2171) );
  XNOR2_X1 DP_mult_206_U1618 ( .A(DP_coeffs_ff_int[11]), .B(DP_mult_206_n2305), 
        .ZN(DP_mult_206_n1811) );
  INV_X1 DP_mult_206_U1617 ( .A(DP_mult_206_n2199), .ZN(DP_mult_206_n2060) );
  AND2_X2 DP_mult_206_U1616 ( .A1(DP_mult_206_n1807), .A2(DP_mult_206_n2245), 
        .ZN(DP_mult_206_n2200) );
  XOR2_X1 DP_mult_206_U1615 ( .A(DP_coeffs_ff_int[1]), .B(DP_coeffs_ff_int[2]), 
        .Z(DP_mult_206_n2190) );
  INV_X1 DP_mult_206_U1614 ( .A(DP_mult_206_n2243), .ZN(DP_mult_206_n2019) );
  XOR2_X1 DP_mult_206_U1613 ( .A(DP_coeffs_ff_int[9]), .B(DP_coeffs_ff_int[10]), .Z(DP_mult_206_n2018) );
  XNOR2_X1 DP_mult_206_U1612 ( .A(DP_mult_206_n827), .B(DP_mult_206_n844), 
        .ZN(DP_mult_206_n2017) );
  XNOR2_X1 DP_mult_206_U1611 ( .A(DP_mult_206_n2052), .B(DP_mult_206_n2017), 
        .ZN(DP_mult_206_n823) );
  XNOR2_X1 DP_mult_206_U1610 ( .A(DP_mult_206_n1001), .B(DP_mult_206_n1394), 
        .ZN(DP_mult_206_n2016) );
  XNOR2_X1 DP_mult_206_U1609 ( .A(DP_mult_206_n2016), .B(DP_mult_206_n1018), 
        .ZN(DP_mult_206_n993) );
  INV_X2 DP_mult_206_U1608 ( .A(DP_mult_206_n2232), .ZN(DP_mult_206_n2231) );
  NAND3_X1 DP_mult_206_U1607 ( .A1(DP_mult_206_n2013), .A2(DP_mult_206_n2014), 
        .A3(DP_mult_206_n2015), .ZN(DP_mult_206_n882) );
  NAND2_X1 DP_mult_206_U1606 ( .A1(DP_mult_206_n893), .A2(DP_mult_206_n889), 
        .ZN(DP_mult_206_n2015) );
  NAND2_X1 DP_mult_206_U1605 ( .A1(DP_mult_206_n906), .A2(DP_mult_206_n889), 
        .ZN(DP_mult_206_n2014) );
  NAND2_X1 DP_mult_206_U1604 ( .A1(DP_mult_206_n906), .A2(DP_mult_206_n893), 
        .ZN(DP_mult_206_n2013) );
  XOR2_X1 DP_mult_206_U1603 ( .A(DP_mult_206_n906), .B(DP_mult_206_n2012), .Z(
        DP_mult_206_n883) );
  XOR2_X1 DP_mult_206_U1602 ( .A(DP_mult_206_n893), .B(DP_mult_206_n889), .Z(
        DP_mult_206_n2012) );
  NAND3_X1 DP_mult_206_U1601 ( .A1(DP_mult_206_n2009), .A2(DP_mult_206_n2010), 
        .A3(DP_mult_206_n2011), .ZN(DP_mult_206_n908) );
  NAND2_X1 DP_mult_206_U1600 ( .A1(DP_mult_206_n1390), .A2(DP_mult_206_n1368), 
        .ZN(DP_mult_206_n2011) );
  NAND2_X1 DP_mult_206_U1599 ( .A1(DP_mult_206_n938), .A2(DP_mult_206_n1368), 
        .ZN(DP_mult_206_n2010) );
  NAND2_X1 DP_mult_206_U1598 ( .A1(DP_mult_206_n938), .A2(DP_mult_206_n1390), 
        .ZN(DP_mult_206_n2009) );
  XOR2_X1 DP_mult_206_U1597 ( .A(DP_mult_206_n938), .B(DP_mult_206_n2008), .Z(
        DP_mult_206_n909) );
  XOR2_X1 DP_mult_206_U1596 ( .A(DP_mult_206_n1390), .B(DP_mult_206_n1368), 
        .Z(DP_mult_206_n2008) );
  NOR2_X1 DP_mult_206_U1595 ( .A1(DP_mult_206_n505), .A2(DP_mult_206_n452), 
        .ZN(DP_mult_206_n450) );
  INV_X2 DP_mult_206_U1594 ( .A(DP_mult_206_n2306), .ZN(DP_mult_206_n2007) );
  XNOR2_X1 DP_mult_206_U1593 ( .A(DP_coeffs_ff_int[3]), .B(DP_mult_206_n2318), 
        .ZN(DP_mult_206_n2121) );
  XNOR2_X1 DP_mult_206_U1592 ( .A(DP_coeffs_ff_int[21]), .B(DP_mult_206_n2280), 
        .ZN(DP_mult_206_n1816) );
  INV_X2 DP_mult_206_U1591 ( .A(DP_mult_206_n2326), .ZN(DP_mult_206_n2325) );
  BUF_X4 DP_mult_206_U1590 ( .A(DP_mult_206_n251), .Z(DP_mult_206_n2270) );
  CLKBUF_X1 DP_mult_206_U1589 ( .A(DP_mult_206_n251), .Z(DP_mult_206_n2269) );
  XOR2_X1 DP_mult_206_U1588 ( .A(DP_coeffs_ff_int[19]), .B(
        DP_coeffs_ff_int[20]), .Z(DP_mult_206_n2080) );
  INV_X1 DP_mult_206_U1587 ( .A(DP_mult_206_n2199), .ZN(DP_mult_206_n2230) );
  INV_X1 DP_mult_206_U1586 ( .A(DP_mult_206_n2196), .ZN(DP_mult_206_n2024) );
  XNOR2_X1 DP_mult_206_U1585 ( .A(DP_coeffs_ff_int[13]), .B(DP_mult_206_n2301), 
        .ZN(DP_mult_206_n1812) );
  AND2_X1 DP_mult_206_U1584 ( .A1(DP_mult_206_n2062), .A2(DP_mult_206_n1814), 
        .ZN(DP_mult_206_n2005) );
  BUF_X1 DP_mult_206_U1583 ( .A(DP_mult_206_n1328), .Z(DP_mult_206_n2003) );
  NOR2_X1 DP_mult_206_U1582 ( .A1(DP_mult_206_n452), .A2(DP_mult_206_n505), 
        .ZN(DP_mult_206_n2002) );
  NAND3_X1 DP_mult_206_U1581 ( .A1(DP_mult_206_n1999), .A2(DP_mult_206_n2000), 
        .A3(DP_mult_206_n2001), .ZN(DP_mult_206_n926) );
  NAND2_X1 DP_mult_206_U1580 ( .A1(DP_mult_206_n952), .A2(DP_mult_206_n933), 
        .ZN(DP_mult_206_n2001) );
  NAND2_X1 DP_mult_206_U1579 ( .A1(DP_mult_206_n937), .A2(DP_mult_206_n933), 
        .ZN(DP_mult_206_n2000) );
  NAND2_X1 DP_mult_206_U1578 ( .A1(DP_mult_206_n937), .A2(DP_mult_206_n952), 
        .ZN(DP_mult_206_n1999) );
  NAND3_X1 DP_mult_206_U1577 ( .A1(DP_mult_206_n1996), .A2(DP_mult_206_n1997), 
        .A3(DP_mult_206_n1998), .ZN(DP_mult_206_n932) );
  NAND2_X1 DP_mult_206_U1576 ( .A1(DP_mult_206_n1435), .A2(DP_mult_206_n1413), 
        .ZN(DP_mult_206_n1998) );
  NAND2_X1 DP_mult_206_U1575 ( .A1(DP_mult_206_n1325), .A2(DP_mult_206_n1413), 
        .ZN(DP_mult_206_n1997) );
  NAND2_X1 DP_mult_206_U1574 ( .A1(DP_mult_206_n1325), .A2(DP_mult_206_n1435), 
        .ZN(DP_mult_206_n1996) );
  XOR2_X1 DP_mult_206_U1573 ( .A(DP_mult_206_n1995), .B(DP_mult_206_n933), .Z(
        DP_mult_206_n927) );
  XOR2_X1 DP_mult_206_U1572 ( .A(DP_mult_206_n937), .B(DP_mult_206_n952), .Z(
        DP_mult_206_n1995) );
  XOR2_X1 DP_mult_206_U1571 ( .A(DP_mult_206_n1994), .B(DP_mult_206_n1413), 
        .Z(DP_mult_206_n933) );
  XOR2_X1 DP_mult_206_U1570 ( .A(DP_mult_206_n1325), .B(DP_mult_206_n1435), 
        .Z(DP_mult_206_n1994) );
  INV_X1 DP_mult_206_U1569 ( .A(DP_mult_206_n2191), .ZN(DP_mult_206_n2261) );
  XNOR2_X1 DP_mult_206_U1568 ( .A(DP_mult_206_n1056), .B(DP_mult_206_n1043), 
        .ZN(DP_mult_206_n1993) );
  XNOR2_X1 DP_mult_206_U1567 ( .A(DP_mult_206_n1041), .B(DP_mult_206_n1993), 
        .ZN(DP_mult_206_n1039) );
  CLKBUF_X1 DP_mult_206_U1566 ( .A(DP_mult_206_n839), .Z(DP_mult_206_n1992) );
  INV_X1 DP_mult_206_U1565 ( .A(DP_mult_206_n2249), .ZN(DP_mult_206_n1991) );
  AOI21_X1 DP_mult_206_U1564 ( .B1(DP_mult_206_n581), .B2(DP_mult_206_n567), 
        .A(DP_mult_206_n568), .ZN(DP_mult_206_n566) );
  XOR2_X1 DP_mult_206_U1563 ( .A(DP_coeffs_ff_int[11]), .B(
        DP_coeffs_ff_int[12]), .Z(DP_mult_206_n1990) );
  INV_X2 DP_mult_206_U1562 ( .A(DP_mult_206_n2195), .ZN(DP_mult_206_n2168) );
  OR2_X2 DP_mult_206_U1561 ( .A1(DP_mult_206_n775), .A2(DP_mult_206_n788), 
        .ZN(DP_mult_206_n1989) );
  XNOR2_X1 DP_mult_206_U1560 ( .A(DP_coeffs_ff_int[5]), .B(DP_mult_206_n2317), 
        .ZN(DP_mult_206_n1808) );
  INV_X1 DP_mult_206_U1559 ( .A(DP_mult_206_n2196), .ZN(DP_mult_206_n1987) );
  INV_X1 DP_mult_206_U1558 ( .A(DP_mult_206_n2196), .ZN(DP_mult_206_n1988) );
  INV_X2 DP_mult_206_U1557 ( .A(DP_mult_206_n2323), .ZN(DP_mult_206_n2320) );
  XOR2_X1 DP_mult_206_U1556 ( .A(DP_coeffs_ff_int[3]), .B(DP_coeffs_ff_int[4]), 
        .Z(DP_mult_206_n2120) );
  INV_X2 DP_mult_206_U1555 ( .A(DP_mult_206_n2286), .ZN(DP_mult_206_n2283) );
  INV_X1 DP_mult_206_U1554 ( .A(DP_mult_206_n2281), .ZN(DP_mult_206_n1985) );
  INV_X1 DP_mult_206_U1553 ( .A(DP_mult_206_n2089), .ZN(DP_mult_206_n2252) );
  INV_X1 DP_mult_206_U1552 ( .A(DP_mult_206_n2196), .ZN(DP_mult_206_n2228) );
  INV_X2 DP_mult_206_U1551 ( .A(DP_mult_206_n2326), .ZN(DP_mult_206_n2324) );
  NOR2_X1 DP_mult_206_U1550 ( .A1(DP_mult_206_n963), .A2(DP_mult_206_n982), 
        .ZN(DP_mult_206_n558) );
  NOR2_X1 DP_mult_206_U1549 ( .A1(DP_mult_206_n963), .A2(DP_mult_206_n982), 
        .ZN(DP_mult_206_n1984) );
  AND2_X1 DP_mult_206_U1548 ( .A1(DP_mult_206_n535), .A2(DP_mult_206_n2125), 
        .ZN(DP_mult_206_n1983) );
  XNOR2_X1 DP_mult_206_U1547 ( .A(DP_mult_206_n536), .B(DP_mult_206_n1983), 
        .ZN(DP_pipe0_coeff_pipe00[3]) );
  XNOR2_X1 DP_mult_206_U1546 ( .A(DP_coeffs_ff_int[9]), .B(DP_mult_206_n2310), 
        .ZN(DP_mult_206_n1810) );
  INV_X2 DP_mult_206_U1545 ( .A(DP_mult_206_n2005), .ZN(DP_mult_206_n2235) );
  INV_X2 DP_mult_206_U1544 ( .A(DP_mult_206_n1982), .ZN(DP_mult_206_n2264) );
  INV_X1 DP_mult_206_U1543 ( .A(DP_mult_206_n2262), .ZN(DP_mult_206_n1982) );
  INV_X1 DP_mult_206_U1542 ( .A(DP_mult_206_n566), .ZN(DP_mult_206_n1981) );
  AND2_X1 DP_mult_206_U1541 ( .A1(DP_mult_206_n1978), .A2(DP_mult_206_n559), 
        .ZN(DP_mult_206_n1980) );
  XNOR2_X1 DP_mult_206_U1540 ( .A(DP_mult_206_n560), .B(DP_mult_206_n1980), 
        .ZN(DP_pipe0_coeff_pipe00[0]) );
  AND2_X1 DP_mult_206_U1539 ( .A1(DP_mult_206_n550), .A2(DP_mult_206_n674), 
        .ZN(DP_mult_206_n1979) );
  XNOR2_X1 DP_mult_206_U1538 ( .A(DP_mult_206_n551), .B(DP_mult_206_n1979), 
        .ZN(DP_pipe0_coeff_pipe00[1]) );
  OR2_X1 DP_mult_206_U1537 ( .A1(DP_mult_206_n963), .A2(DP_mult_206_n982), 
        .ZN(DP_mult_206_n1978) );
  OR2_X1 DP_mult_206_U1536 ( .A1(DP_mult_206_n1151), .A2(DP_mult_206_n1158), 
        .ZN(DP_mult_206_n1977) );
  AND2_X1 DP_mult_206_U1535 ( .A1(DP_mult_206_n1111), .A2(DP_mult_206_n1122), 
        .ZN(DP_mult_206_n1976) );
  AND2_X1 DP_mult_206_U1534 ( .A1(DP_mult_206_n1133), .A2(DP_mult_206_n1142), 
        .ZN(DP_mult_206_n1975) );
  AND2_X1 DP_mult_206_U1533 ( .A1(DP_mult_206_n1055), .A2(DP_mult_206_n1070), 
        .ZN(DP_mult_206_n1974) );
  AND2_X1 DP_mult_206_U1532 ( .A1(DP_mult_206_n1179), .A2(DP_mult_206_n1433), 
        .ZN(DP_mult_206_n1973) );
  AND2_X1 DP_mult_206_U1531 ( .A1(DP_mult_206_n1021), .A2(DP_mult_206_n1038), 
        .ZN(DP_mult_206_n1972) );
  AND2_X1 DP_mult_206_U1530 ( .A1(DP_mult_206_n1457), .A2(DP_mult_206_n1480), 
        .ZN(DP_mult_206_n1971) );
  AND2_X1 DP_mult_206_U1529 ( .A1(DP_mult_206_n1151), .A2(DP_mult_206_n1158), 
        .ZN(DP_mult_206_n1970) );
  AND2_X1 DP_mult_206_U1528 ( .A1(DP_mult_206_n1123), .A2(DP_mult_206_n1132), 
        .ZN(DP_mult_206_n1969) );
  AND2_X1 DP_mult_206_U1527 ( .A1(DP_mult_206_n1143), .A2(DP_mult_206_n1150), 
        .ZN(DP_mult_206_n1968) );
  OR2_X1 DP_mult_206_U1526 ( .A1(DP_mult_206_n1179), .A2(DP_mult_206_n1433), 
        .ZN(DP_mult_206_n1967) );
  AND2_X1 DP_mult_206_U1525 ( .A1(DP_mult_206_n1039), .A2(DP_mult_206_n1054), 
        .ZN(DP_mult_206_n1966) );
  OR2_X1 DP_mult_206_U1524 ( .A1(DP_mult_206_n1457), .A2(DP_mult_206_n1480), 
        .ZN(DP_mult_206_n1965) );
  AND2_X1 DP_mult_206_U1523 ( .A1(DP_mult_206_n1193), .A2(DP_mult_206_n1481), 
        .ZN(DP_mult_206_n1964) );
  INV_X1 DP_mult_206_U1522 ( .A(DP_mult_206_n2119), .ZN(DP_mult_206_n2127) );
  NAND3_X1 DP_mult_206_U1521 ( .A1(DP_mult_206_n2097), .A2(DP_mult_206_n2098), 
        .A3(DP_mult_206_n2099), .ZN(DP_mult_206_n954) );
  OR2_X1 DP_mult_206_U1520 ( .A1(DP_mult_206_n1055), .A2(DP_mult_206_n1070), 
        .ZN(DP_mult_206_n2175) );
  NAND3_X1 DP_mult_206_U1519 ( .A1(DP_mult_206_n2138), .A2(DP_mult_206_n2139), 
        .A3(DP_mult_206_n2140), .ZN(DP_mult_206_n994) );
  INV_X1 DP_mult_206_U1518 ( .A(DP_mult_206_n2036), .ZN(DP_mult_206_n2132) );
  INV_X2 DP_mult_206_U1517 ( .A(DP_mult_206_n2318), .ZN(DP_mult_206_n2314) );
  INV_X1 DP_mult_206_U1516 ( .A(DP_mult_206_n2200), .ZN(DP_mult_206_n2126) );
  CLKBUF_X1 DP_mult_206_U1515 ( .A(DP_mult_206_n525), .Z(DP_mult_206_n1963) );
  INV_X2 DP_mult_206_U1514 ( .A(DP_mult_206_n2136), .ZN(DP_mult_206_n2104) );
  INV_X1 DP_mult_206_U1513 ( .A(DP_mult_206_n2136), .ZN(DP_mult_206_n2220) );
  NAND3_X1 DP_mult_206_U1512 ( .A1(DP_mult_206_n1960), .A2(DP_mult_206_n1961), 
        .A3(DP_mult_206_n1962), .ZN(DP_mult_206_n818) );
  NAND2_X1 DP_mult_206_U1511 ( .A1(DP_mult_206_n1209), .A2(DP_mult_206_n1363), 
        .ZN(DP_mult_206_n1962) );
  NAND2_X1 DP_mult_206_U1510 ( .A1(DP_mult_206_n836), .A2(DP_mult_206_n1363), 
        .ZN(DP_mult_206_n1961) );
  NAND2_X1 DP_mult_206_U1509 ( .A1(DP_mult_206_n836), .A2(DP_mult_206_n1209), 
        .ZN(DP_mult_206_n1960) );
  XOR2_X1 DP_mult_206_U1508 ( .A(DP_mult_206_n836), .B(DP_mult_206_n1959), .Z(
        DP_mult_206_n819) );
  XOR2_X1 DP_mult_206_U1507 ( .A(DP_mult_206_n1209), .B(DP_mult_206_n1363), 
        .Z(DP_mult_206_n1959) );
  BUF_X2 DP_mult_206_U1506 ( .A(DP_mult_206_n2036), .Z(DP_mult_206_n2201) );
  NAND2_X1 DP_mult_206_U1505 ( .A1(DP_mult_206_n1957), .A2(DP_mult_206_n1958), 
        .ZN(DP_mult_206_n1370) );
  OR2_X1 DP_mult_206_U1504 ( .A1(DP_mult_206_n1665), .A2(DP_mult_206_n2201), 
        .ZN(DP_mult_206_n1958) );
  OR2_X1 DP_mult_206_U1503 ( .A1(DP_mult_206_n2234), .A2(DP_mult_206_n1666), 
        .ZN(DP_mult_206_n1957) );
  NAND3_X1 DP_mult_206_U1502 ( .A1(DP_mult_206_n1954), .A2(DP_mult_206_n1955), 
        .A3(DP_mult_206_n1956), .ZN(DP_mult_206_n956) );
  NAND2_X1 DP_mult_206_U1501 ( .A1(DP_mult_206_n1436), .A2(DP_mult_206_n1459), 
        .ZN(DP_mult_206_n1956) );
  NAND2_X1 DP_mult_206_U1500 ( .A1(DP_mult_206_n1370), .A2(DP_mult_206_n1459), 
        .ZN(DP_mult_206_n1955) );
  NAND2_X1 DP_mult_206_U1499 ( .A1(DP_mult_206_n1370), .A2(DP_mult_206_n1436), 
        .ZN(DP_mult_206_n1954) );
  XOR2_X1 DP_mult_206_U1498 ( .A(DP_mult_206_n1370), .B(DP_mult_206_n1953), 
        .Z(DP_mult_206_n957) );
  XOR2_X1 DP_mult_206_U1497 ( .A(DP_mult_206_n1436), .B(DP_mult_206_n1459), 
        .Z(DP_mult_206_n1953) );
  INV_X1 DP_mult_206_U1496 ( .A(DP_mult_206_n2300), .ZN(DP_mult_206_n2297) );
  INV_X1 DP_mult_206_U1495 ( .A(DP_mult_206_n1930), .ZN(DP_mult_206_n2249) );
  OAI22_X1 DP_mult_206_U1494 ( .A1(DP_mult_206_n2240), .A2(DP_mult_206_n1733), 
        .B1(DP_mult_206_n1732), .B2(DP_mult_206_n2267), .ZN(DP_mult_206_n1952)
         );
  INV_X2 DP_mult_206_U1493 ( .A(DP_mult_206_n2295), .ZN(DP_mult_206_n2292) );
  INV_X2 DP_mult_206_U1492 ( .A(DP_mult_206_n1990), .ZN(DP_mult_206_n2258) );
  INV_X2 DP_mult_206_U1491 ( .A(DP_mult_206_n2189), .ZN(DP_mult_206_n1950) );
  INV_X2 DP_mult_206_U1490 ( .A(DP_mult_206_n2189), .ZN(DP_mult_206_n1951) );
  CLKBUF_X1 DP_mult_206_U1489 ( .A(DP_mult_206_n2276), .Z(DP_mult_206_n1949)
         );
  XNOR2_X1 DP_mult_206_U1488 ( .A(DP_coeffs_ff_int[2]), .B(DP_coeffs_ff_int[1]), .ZN(DP_mult_206_n1986) );
  INV_X2 DP_mult_206_U1487 ( .A(DP_mult_206_n1948), .ZN(DP_mult_206_n2137) );
  NAND2_X2 DP_mult_206_U1486 ( .A1(DP_mult_206_n1806), .A2(DP_mult_206_n2243), 
        .ZN(DP_mult_206_n1948) );
  AND2_X1 DP_mult_206_U1485 ( .A1(DP_mult_206_n673), .A2(DP_mult_206_n543), 
        .ZN(DP_mult_206_n1947) );
  XNOR2_X1 DP_mult_206_U1484 ( .A(DP_mult_206_n544), .B(DP_mult_206_n1947), 
        .ZN(DP_pipe0_coeff_pipe00[2]) );
  INV_X1 DP_mult_206_U1483 ( .A(DP_mult_206_n2251), .ZN(DP_mult_206_n1946) );
  AOI21_X1 DP_mult_206_U1482 ( .B1(DP_mult_206_n581), .B2(DP_mult_206_n567), 
        .A(DP_mult_206_n568), .ZN(DP_mult_206_n1945) );
  AND2_X1 DP_mult_206_U1481 ( .A1(DP_mult_206_n552), .A2(DP_mult_206_n674), 
        .ZN(DP_mult_206_n545) );
  INV_X2 DP_mult_206_U1480 ( .A(DP_mult_206_n2268), .ZN(DP_mult_206_n2265) );
  INV_X1 DP_mult_206_U1479 ( .A(DP_mult_206_n2268), .ZN(DP_mult_206_n2267) );
  AND2_X1 DP_mult_206_U1478 ( .A1(DP_mult_206_n1808), .A2(DP_mult_206_n2248), 
        .ZN(DP_mult_206_n2198) );
  INV_X1 DP_mult_206_U1477 ( .A(DP_mult_206_n1943), .ZN(DP_mult_206_n1944) );
  AND2_X2 DP_mult_206_U1476 ( .A1(DP_mult_206_n1808), .A2(DP_mult_206_n2248), 
        .ZN(DP_mult_206_n1943) );
  INV_X1 DP_mult_206_U1475 ( .A(DP_mult_206_n2193), .ZN(DP_mult_206_n2234) );
  INV_X1 DP_mult_206_U1474 ( .A(DP_mult_206_n2193), .ZN(DP_mult_206_n1941) );
  INV_X1 DP_mult_206_U1473 ( .A(DP_mult_206_n2193), .ZN(DP_mult_206_n1942) );
  NAND3_X1 DP_mult_206_U1472 ( .A1(DP_mult_206_n1954), .A2(DP_mult_206_n1955), 
        .A3(DP_mult_206_n1956), .ZN(DP_mult_206_n1940) );
  NAND3_X1 DP_mult_206_U1471 ( .A1(DP_mult_206_n1937), .A2(DP_mult_206_n1938), 
        .A3(DP_mult_206_n1939), .ZN(DP_mult_206_n808) );
  NAND2_X1 DP_mult_206_U1470 ( .A1(DP_mult_206_n813), .A2(DP_mult_206_n819), 
        .ZN(DP_mult_206_n1939) );
  NAND2_X1 DP_mult_206_U1469 ( .A1(DP_mult_206_n828), .A2(DP_mult_206_n819), 
        .ZN(DP_mult_206_n1938) );
  NAND2_X1 DP_mult_206_U1468 ( .A1(DP_mult_206_n828), .A2(DP_mult_206_n813), 
        .ZN(DP_mult_206_n1937) );
  XOR2_X1 DP_mult_206_U1467 ( .A(DP_mult_206_n828), .B(DP_mult_206_n1936), .Z(
        DP_mult_206_n809) );
  XOR2_X1 DP_mult_206_U1466 ( .A(DP_mult_206_n813), .B(DP_mult_206_n819), .Z(
        DP_mult_206_n1936) );
  AND2_X2 DP_mult_206_U1465 ( .A1(DP_mult_206_n2062), .A2(DP_mult_206_n1814), 
        .ZN(DP_mult_206_n2006) );
  CLKBUF_X1 DP_mult_206_U1464 ( .A(DP_mult_206_n490), .Z(DP_mult_206_n1935) );
  CLKBUF_X1 DP_mult_206_U1463 ( .A(DP_mult_206_n886), .Z(DP_mult_206_n1934) );
  OR2_X2 DP_mult_206_U1462 ( .A1(DP_mult_206_n2236), .A2(DP_mult_206_n1683), 
        .ZN(DP_mult_206_n2029) );
  AND2_X2 DP_mult_206_U1461 ( .A1(DP_mult_206_n2029), .A2(DP_mult_206_n2030), 
        .ZN(DP_mult_206_n2004) );
  CLKBUF_X1 DP_mult_206_U1460 ( .A(DP_mult_206_n547), .Z(DP_mult_206_n1933) );
  CLKBUF_X1 DP_mult_206_U1459 ( .A(DP_mult_206_n1254), .Z(DP_mult_206_n2034)
         );
  INV_X1 DP_mult_206_U1458 ( .A(DP_mult_206_n2200), .ZN(DP_mult_206_n2222) );
  NOR2_X2 DP_mult_206_U1457 ( .A1(DP_mult_206_n919), .A2(DP_mult_206_n940), 
        .ZN(DP_mult_206_n542) );
  XNOR2_X1 DP_mult_206_U1456 ( .A(DP_coeffs_ff_int[11]), .B(
        DP_coeffs_ff_int[12]), .ZN(DP_mult_206_n1932) );
  INV_X1 DP_mult_206_U1455 ( .A(DP_mult_206_n2268), .ZN(DP_mult_206_n2266) );
  INV_X1 DP_mult_206_U1454 ( .A(DP_mult_206_n2031), .ZN(DP_mult_206_n1931) );
  BUF_X1 DP_mult_206_U1453 ( .A(DP_mult_206_n2226), .Z(DP_mult_206_n2202) );
  INV_X2 DP_mult_206_U1452 ( .A(DP_mult_206_n2195), .ZN(DP_mult_206_n2226) );
  INV_X2 DP_mult_206_U1451 ( .A(DP_mult_206_n1946), .ZN(DP_mult_206_n2253) );
  INV_X2 DP_mult_206_U1450 ( .A(DP_mult_206_n2195), .ZN(DP_mult_206_n2169) );
  XOR2_X1 DP_mult_206_U1449 ( .A(DP_coeffs_ff_int[5]), .B(DP_coeffs_ff_int[6]), 
        .Z(DP_mult_206_n1930) );
  XOR2_X1 DP_mult_206_U1448 ( .A(DP_coeffs_ff_int[5]), .B(DP_coeffs_ff_int[6]), 
        .Z(DP_mult_206_n1929) );
  HA_X1 DP_mult_206_U798 ( .A(DP_mult_206_n1456), .B(DP_mult_206_n1479), .CO(
        DP_mult_206_n1180), .S(DP_mult_206_n1181) );
  FA_X1 DP_mult_206_U797 ( .A(DP_mult_206_n1455), .B(DP_mult_206_n1478), .CI(
        DP_mult_206_n1180), .CO(DP_mult_206_n1178), .S(DP_mult_206_n1179) );
  HA_X1 DP_mult_206_U796 ( .A(DP_mult_206_n1432), .B(DP_mult_206_n1477), .CO(
        DP_mult_206_n1176), .S(DP_mult_206_n1177) );
  FA_X1 DP_mult_206_U795 ( .A(DP_mult_206_n1191), .B(DP_mult_206_n1454), .CI(
        DP_mult_206_n1177), .CO(DP_mult_206_n1174), .S(DP_mult_206_n1175) );
  FA_X1 DP_mult_206_U794 ( .A(DP_mult_206_n1476), .B(DP_mult_206_n1453), .CI(
        DP_mult_206_n1431), .CO(DP_mult_206_n1172), .S(DP_mult_206_n1173) );
  FA_X1 DP_mult_206_U793 ( .A(DP_mult_206_n1409), .B(DP_mult_206_n1176), .CI(
        DP_mult_206_n1173), .CO(DP_mult_206_n1170), .S(DP_mult_206_n1171) );
  HA_X1 DP_mult_206_U792 ( .A(DP_mult_206_n1408), .B(DP_mult_206_n1430), .CO(
        DP_mult_206_n1168), .S(DP_mult_206_n1169) );
  FA_X1 DP_mult_206_U791 ( .A(DP_mult_206_n1452), .B(DP_mult_206_n1475), .CI(
        DP_mult_206_n1190), .CO(DP_mult_206_n1166), .S(DP_mult_206_n1167) );
  FA_X1 DP_mult_206_U790 ( .A(DP_mult_206_n1172), .B(DP_mult_206_n1169), .CI(
        DP_mult_206_n1167), .CO(DP_mult_206_n1164), .S(DP_mult_206_n1165) );
  FA_X1 DP_mult_206_U789 ( .A(DP_mult_206_n1451), .B(DP_mult_206_n1474), .CI(
        DP_mult_206_n1407), .CO(DP_mult_206_n1162), .S(DP_mult_206_n1163) );
  FA_X1 DP_mult_206_U788 ( .A(DP_mult_206_n1168), .B(DP_mult_206_n1429), .CI(
        DP_mult_206_n1166), .CO(DP_mult_206_n1160), .S(DP_mult_206_n1161) );
  FA_X1 DP_mult_206_U787 ( .A(DP_mult_206_n1163), .B(DP_mult_206_n1385), .CI(
        DP_mult_206_n1164), .CO(DP_mult_206_n1158), .S(DP_mult_206_n1159) );
  HA_X1 DP_mult_206_U786 ( .A(DP_mult_206_n1384), .B(DP_mult_206_n1406), .CO(
        DP_mult_206_n1156), .S(DP_mult_206_n1157) );
  FA_X1 DP_mult_206_U785 ( .A(DP_mult_206_n1450), .B(DP_mult_206_n1428), .CI(
        DP_mult_206_n1189), .CO(DP_mult_206_n1154), .S(DP_mult_206_n1155) );
  FA_X1 DP_mult_206_U784 ( .A(DP_mult_206_n1157), .B(DP_mult_206_n1473), .CI(
        DP_mult_206_n1162), .CO(DP_mult_206_n1152), .S(DP_mult_206_n1153) );
  FA_X1 DP_mult_206_U783 ( .A(DP_mult_206_n1160), .B(DP_mult_206_n1155), .CI(
        DP_mult_206_n1153), .CO(DP_mult_206_n1150), .S(DP_mult_206_n1151) );
  FA_X1 DP_mult_206_U782 ( .A(DP_mult_206_n1383), .B(DP_mult_206_n1472), .CI(
        DP_mult_206_n1405), .CO(DP_mult_206_n1148), .S(DP_mult_206_n1149) );
  FA_X1 DP_mult_206_U781 ( .A(DP_mult_206_n1427), .B(DP_mult_206_n1449), .CI(
        DP_mult_206_n1156), .CO(DP_mult_206_n1146), .S(DP_mult_206_n1147) );
  FA_X1 DP_mult_206_U780 ( .A(DP_mult_206_n1361), .B(DP_mult_206_n1154), .CI(
        DP_mult_206_n1149), .CO(DP_mult_206_n1144), .S(DP_mult_206_n1145) );
  FA_X1 DP_mult_206_U779 ( .A(DP_mult_206_n1152), .B(DP_mult_206_n1147), .CI(
        DP_mult_206_n1145), .CO(DP_mult_206_n1142), .S(DP_mult_206_n1143) );
  HA_X1 DP_mult_206_U778 ( .A(DP_mult_206_n1360), .B(DP_mult_206_n1382), .CO(
        DP_mult_206_n1140), .S(DP_mult_206_n1141) );
  FA_X1 DP_mult_206_U777 ( .A(DP_mult_206_n1188), .B(DP_mult_206_n1471), .CI(
        DP_mult_206_n1426), .CO(DP_mult_206_n1138), .S(DP_mult_206_n1139) );
  FA_X1 DP_mult_206_U776 ( .A(DP_mult_206_n1404), .B(DP_mult_206_n1448), .CI(
        DP_mult_206_n1141), .CO(DP_mult_206_n1136), .S(DP_mult_206_n1137) );
  FA_X1 DP_mult_206_U775 ( .A(DP_mult_206_n1146), .B(DP_mult_206_n1148), .CI(
        DP_mult_206_n1139), .CO(DP_mult_206_n1134), .S(DP_mult_206_n1135) );
  FA_X1 DP_mult_206_U774 ( .A(DP_mult_206_n1144), .B(DP_mult_206_n1137), .CI(
        DP_mult_206_n1135), .CO(DP_mult_206_n1132), .S(DP_mult_206_n1133) );
  FA_X1 DP_mult_206_U773 ( .A(DP_mult_206_n1359), .B(DP_mult_206_n1470), .CI(
        DP_mult_206_n1381), .CO(DP_mult_206_n1130), .S(DP_mult_206_n1131) );
  FA_X1 DP_mult_206_U772 ( .A(DP_mult_206_n1403), .B(DP_mult_206_n1447), .CI(
        DP_mult_206_n1425), .CO(DP_mult_206_n1128), .S(DP_mult_206_n1129) );
  FA_X1 DP_mult_206_U771 ( .A(DP_mult_206_n1138), .B(DP_mult_206_n1140), .CI(
        DP_mult_206_n1337), .CO(DP_mult_206_n1126), .S(DP_mult_206_n1127) );
  FA_X1 DP_mult_206_U770 ( .A(DP_mult_206_n1131), .B(DP_mult_206_n1129), .CI(
        DP_mult_206_n1136), .CO(DP_mult_206_n1124), .S(DP_mult_206_n1125) );
  FA_X1 DP_mult_206_U769 ( .A(DP_mult_206_n1127), .B(DP_mult_206_n1134), .CI(
        DP_mult_206_n1125), .CO(DP_mult_206_n1122), .S(DP_mult_206_n1123) );
  HA_X1 DP_mult_206_U768 ( .A(DP_mult_206_n1336), .B(DP_mult_206_n1358), .CO(
        DP_mult_206_n1120), .S(DP_mult_206_n1121) );
  FA_X1 DP_mult_206_U767 ( .A(DP_mult_206_n1380), .B(DP_mult_206_n1402), .CI(
        DP_mult_206_n1187), .CO(DP_mult_206_n1118), .S(DP_mult_206_n1119) );
  FA_X1 DP_mult_206_U766 ( .A(DP_mult_206_n1424), .B(DP_mult_206_n1469), .CI(
        DP_mult_206_n1446), .CO(DP_mult_206_n1116), .S(DP_mult_206_n1117) );
  FA_X1 DP_mult_206_U765 ( .A(DP_mult_206_n1130), .B(DP_mult_206_n1121), .CI(
        DP_mult_206_n1128), .CO(DP_mult_206_n1114), .S(DP_mult_206_n1115) );
  FA_X1 DP_mult_206_U764 ( .A(DP_mult_206_n1119), .B(DP_mult_206_n1117), .CI(
        DP_mult_206_n1126), .CO(DP_mult_206_n1112), .S(DP_mult_206_n1113) );
  FA_X1 DP_mult_206_U763 ( .A(DP_mult_206_n1124), .B(DP_mult_206_n1115), .CI(
        DP_mult_206_n1113), .CO(DP_mult_206_n1110), .S(DP_mult_206_n1111) );
  FA_X1 DP_mult_206_U762 ( .A(DP_mult_206_n1335), .B(DP_mult_206_n1468), .CI(
        DP_mult_206_n1357), .CO(DP_mult_206_n1108), .S(DP_mult_206_n1109) );
  FA_X1 DP_mult_206_U761 ( .A(DP_mult_206_n1379), .B(DP_mult_206_n1445), .CI(
        DP_mult_206_n1401), .CO(DP_mult_206_n1106), .S(DP_mult_206_n1107) );
  FA_X1 DP_mult_206_U760 ( .A(DP_mult_206_n1120), .B(DP_mult_206_n1423), .CI(
        DP_mult_206_n1118), .CO(DP_mult_206_n1104), .S(DP_mult_206_n1105) );
  FA_X1 DP_mult_206_U759 ( .A(DP_mult_206_n1313), .B(DP_mult_206_n1116), .CI(
        DP_mult_206_n1107), .CO(DP_mult_206_n1102), .S(DP_mult_206_n1103) );
  FA_X1 DP_mult_206_U758 ( .A(DP_mult_206_n1114), .B(DP_mult_206_n1109), .CI(
        DP_mult_206_n1105), .CO(DP_mult_206_n1100), .S(DP_mult_206_n1101) );
  FA_X1 DP_mult_206_U757 ( .A(DP_mult_206_n1103), .B(DP_mult_206_n1112), .CI(
        DP_mult_206_n1101), .CO(DP_mult_206_n1098), .S(DP_mult_206_n1099) );
  HA_X1 DP_mult_206_U756 ( .A(DP_mult_206_n1334), .B(DP_mult_206_n1312), .CO(
        DP_mult_206_n1096), .S(DP_mult_206_n1097) );
  FA_X1 DP_mult_206_U755 ( .A(DP_mult_206_n1467), .B(DP_mult_206_n1400), .CI(
        DP_mult_206_n1186), .CO(DP_mult_206_n1094), .S(DP_mult_206_n1095) );
  FA_X1 DP_mult_206_U754 ( .A(DP_mult_206_n1378), .B(DP_mult_206_n1356), .CI(
        DP_mult_206_n1444), .CO(DP_mult_206_n1092), .S(DP_mult_206_n1093) );
  FA_X1 DP_mult_206_U753 ( .A(DP_mult_206_n1097), .B(DP_mult_206_n1422), .CI(
        DP_mult_206_n1108), .CO(DP_mult_206_n1090), .S(DP_mult_206_n1091) );
  FA_X1 DP_mult_206_U752 ( .A(DP_mult_206_n1093), .B(DP_mult_206_n1106), .CI(
        DP_mult_206_n1095), .CO(DP_mult_206_n1088), .S(DP_mult_206_n1089) );
  FA_X1 DP_mult_206_U751 ( .A(DP_mult_206_n1102), .B(DP_mult_206_n1104), .CI(
        DP_mult_206_n1091), .CO(DP_mult_206_n1086), .S(DP_mult_206_n1087) );
  FA_X1 DP_mult_206_U750 ( .A(DP_mult_206_n1100), .B(DP_mult_206_n1089), .CI(
        DP_mult_206_n1087), .CO(DP_mult_206_n1084), .S(DP_mult_206_n1085) );
  FA_X1 DP_mult_206_U749 ( .A(DP_mult_206_n1311), .B(DP_mult_206_n1466), .CI(
        DP_mult_206_n1333), .CO(DP_mult_206_n1082), .S(DP_mult_206_n1083) );
  FA_X1 DP_mult_206_U748 ( .A(DP_mult_206_n1355), .B(DP_mult_206_n1443), .CI(
        DP_mult_206_n1377), .CO(DP_mult_206_n1080), .S(DP_mult_206_n1081) );
  FA_X1 DP_mult_206_U747 ( .A(DP_mult_206_n1399), .B(DP_mult_206_n1421), .CI(
        DP_mult_206_n1096), .CO(DP_mult_206_n1078), .S(DP_mult_206_n1079) );
  FA_X1 DP_mult_206_U746 ( .A(DP_mult_206_n1092), .B(DP_mult_206_n1094), .CI(
        DP_mult_206_n1289), .CO(DP_mult_206_n1076), .S(DP_mult_206_n1077) );
  FA_X1 DP_mult_206_U745 ( .A(DP_mult_206_n1083), .B(DP_mult_206_n1081), .CI(
        DP_mult_206_n1079), .CO(DP_mult_206_n1074), .S(DP_mult_206_n1075) );
  FA_X1 DP_mult_206_U744 ( .A(DP_mult_206_n1088), .B(DP_mult_206_n1090), .CI(
        DP_mult_206_n1077), .CO(DP_mult_206_n1072), .S(DP_mult_206_n1073) );
  FA_X1 DP_mult_206_U743 ( .A(DP_mult_206_n1086), .B(DP_mult_206_n1075), .CI(
        DP_mult_206_n1073), .CO(DP_mult_206_n1070), .S(DP_mult_206_n1071) );
  HA_X1 DP_mult_206_U742 ( .A(DP_mult_206_n1288), .B(DP_mult_206_n1310), .CO(
        DP_mult_206_n1068), .S(DP_mult_206_n1069) );
  FA_X1 DP_mult_206_U741 ( .A(DP_mult_206_n1465), .B(DP_mult_206_n1376), .CI(
        DP_mult_206_n1185), .CO(DP_mult_206_n1066), .S(DP_mult_206_n1067) );
  FA_X1 DP_mult_206_U740 ( .A(DP_mult_206_n1442), .B(DP_mult_206_n1332), .CI(
        DP_mult_206_n1354), .CO(DP_mult_206_n1064), .S(DP_mult_206_n1065) );
  FA_X1 DP_mult_206_U739 ( .A(DP_mult_206_n1398), .B(DP_mult_206_n1420), .CI(
        DP_mult_206_n1069), .CO(DP_mult_206_n1062), .S(DP_mult_206_n1063) );
  FA_X1 DP_mult_206_U738 ( .A(DP_mult_206_n1080), .B(DP_mult_206_n1082), .CI(
        DP_mult_206_n1078), .CO(DP_mult_206_n1060), .S(DP_mult_206_n1061) );
  FA_X1 DP_mult_206_U737 ( .A(DP_mult_206_n1067), .B(DP_mult_206_n1065), .CI(
        DP_mult_206_n1076), .CO(DP_mult_206_n1058), .S(DP_mult_206_n1059) );
  FA_X1 DP_mult_206_U736 ( .A(DP_mult_206_n1074), .B(DP_mult_206_n1063), .CI(
        DP_mult_206_n1061), .CO(DP_mult_206_n1056), .S(DP_mult_206_n1057) );
  FA_X1 DP_mult_206_U735 ( .A(DP_mult_206_n1072), .B(DP_mult_206_n1059), .CI(
        DP_mult_206_n1057), .CO(DP_mult_206_n1054), .S(DP_mult_206_n1055) );
  FA_X1 DP_mult_206_U734 ( .A(DP_mult_206_n1309), .B(DP_mult_206_n1464), .CI(
        DP_mult_206_n1287), .CO(DP_mult_206_n1052), .S(DP_mult_206_n1053) );
  FA_X1 DP_mult_206_U733 ( .A(DP_mult_206_n1331), .B(DP_mult_206_n1353), .CI(
        DP_mult_206_n1375), .CO(DP_mult_206_n1050), .S(DP_mult_206_n1051) );
  FA_X1 DP_mult_206_U732 ( .A(DP_mult_206_n1397), .B(DP_mult_206_n1441), .CI(
        DP_mult_206_n1419), .CO(DP_mult_206_n1048), .S(DP_mult_206_n1049) );
  FA_X1 DP_mult_206_U731 ( .A(DP_mult_206_n1064), .B(DP_mult_206_n1068), .CI(
        DP_mult_206_n1066), .CO(DP_mult_206_n1046), .S(DP_mult_206_n1047) );
  FA_X1 DP_mult_206_U730 ( .A(DP_mult_206_n1049), .B(DP_mult_206_n1265), .CI(
        DP_mult_206_n1051), .CO(DP_mult_206_n1044), .S(DP_mult_206_n1045) );
  FA_X1 DP_mult_206_U729 ( .A(DP_mult_206_n1062), .B(DP_mult_206_n1053), .CI(
        DP_mult_206_n1060), .CO(DP_mult_206_n1042), .S(DP_mult_206_n1043) );
  FA_X1 DP_mult_206_U728 ( .A(DP_mult_206_n1058), .B(DP_mult_206_n1047), .CI(
        DP_mult_206_n1045), .CO(DP_mult_206_n1040), .S(DP_mult_206_n1041) );
  HA_X1 DP_mult_206_U726 ( .A(DP_mult_206_n1264), .B(DP_mult_206_n1286), .CO(
        DP_mult_206_n1036), .S(DP_mult_206_n1037) );
  FA_X1 DP_mult_206_U725 ( .A(DP_mult_206_n1308), .B(DP_mult_206_n1184), .CI(
        DP_mult_206_n1374), .CO(DP_mult_206_n1034), .S(DP_mult_206_n1035) );
  FA_X1 DP_mult_206_U724 ( .A(DP_mult_206_n1330), .B(DP_mult_206_n1396), .CI(
        DP_mult_206_n1463), .CO(DP_mult_206_n1032), .S(DP_mult_206_n1033) );
  FA_X1 DP_mult_206_U723 ( .A(DP_mult_206_n1352), .B(DP_mult_206_n1440), .CI(
        DP_mult_206_n1418), .CO(DP_mult_206_n1030), .S(DP_mult_206_n1031) );
  FA_X1 DP_mult_206_U722 ( .A(DP_mult_206_n1037), .B(DP_mult_206_n1052), .CI(
        DP_mult_206_n1050), .CO(DP_mult_206_n1028), .S(DP_mult_206_n1029) );
  FA_X1 DP_mult_206_U721 ( .A(DP_mult_206_n1031), .B(DP_mult_206_n1048), .CI(
        DP_mult_206_n1033), .CO(DP_mult_206_n1026), .S(DP_mult_206_n1027) );
  FA_X1 DP_mult_206_U720 ( .A(DP_mult_206_n1046), .B(DP_mult_206_n1035), .CI(
        DP_mult_206_n1029), .CO(DP_mult_206_n1024), .S(DP_mult_206_n1025) );
  FA_X1 DP_mult_206_U716 ( .A(DP_mult_206_n1373), .B(DP_mult_206_n1307), .CI(
        DP_mult_206_n1329), .CO(DP_mult_206_n1016), .S(DP_mult_206_n1017) );
  FA_X1 DP_mult_206_U715 ( .A(DP_mult_206_n1395), .B(DP_mult_206_n1462), .CI(
        DP_mult_206_n1417), .CO(DP_mult_206_n1014), .S(DP_mult_206_n1015) );
  FA_X1 DP_mult_206_U714 ( .A(DP_mult_206_n1036), .B(DP_mult_206_n1439), .CI(
        DP_mult_206_n1032), .CO(DP_mult_206_n1012), .S(DP_mult_206_n1013) );
  FA_X1 DP_mult_206_U713 ( .A(DP_mult_206_n1241), .B(DP_mult_206_n1034), .CI(
        DP_mult_206_n1030), .CO(DP_mult_206_n1010), .S(DP_mult_206_n1011) );
  FA_X1 DP_mult_206_U712 ( .A(DP_mult_206_n1017), .B(DP_mult_206_n1015), .CI(
        DP_mult_206_n1019), .CO(DP_mult_206_n1008), .S(DP_mult_206_n1009) );
  FA_X1 DP_mult_206_U711 ( .A(DP_mult_206_n1013), .B(DP_mult_206_n1028), .CI(
        DP_mult_206_n1026), .CO(DP_mult_206_n1006), .S(DP_mult_206_n1007) );
  FA_X1 DP_mult_206_U710 ( .A(DP_mult_206_n1009), .B(DP_mult_206_n1011), .CI(
        DP_mult_206_n1024), .CO(DP_mult_206_n1004), .S(DP_mult_206_n1005) );
  FA_X1 DP_mult_206_U709 ( .A(DP_mult_206_n1022), .B(DP_mult_206_n1007), .CI(
        DP_mult_206_n1005), .CO(DP_mult_206_n1002), .S(DP_mult_206_n1003) );
  HA_X1 DP_mult_206_U708 ( .A(DP_mult_206_n1262), .B(DP_mult_206_n1240), .CO(
        DP_mult_206_n1000), .S(DP_mult_206_n1001) );
  FA_X1 DP_mult_206_U707 ( .A(DP_mult_206_n1461), .B(DP_mult_206_n1350), .CI(
        DP_mult_206_n1183), .CO(DP_mult_206_n998), .S(DP_mult_206_n999) );
  FA_X1 DP_mult_206_U706 ( .A(DP_mult_206_n1284), .B(DP_mult_206_n1438), .CI(
        DP_mult_206_n1372), .CO(DP_mult_206_n996), .S(DP_mult_206_n997) );
  FA_X1 DP_mult_206_U703 ( .A(DP_mult_206_n1014), .B(DP_mult_206_n1016), .CI(
        DP_mult_206_n995), .CO(DP_mult_206_n990), .S(DP_mult_206_n991) );
  FA_X1 DP_mult_206_U702 ( .A(DP_mult_206_n999), .B(DP_mult_206_n997), .CI(
        DP_mult_206_n1012), .CO(DP_mult_206_n988), .S(DP_mult_206_n989) );
  FA_X1 DP_mult_206_U701 ( .A(DP_mult_206_n993), .B(DP_mult_206_n1010), .CI(
        DP_mult_206_n1008), .CO(DP_mult_206_n986), .S(DP_mult_206_n987) );
  FA_X1 DP_mult_206_U700 ( .A(DP_mult_206_n989), .B(DP_mult_206_n991), .CI(
        DP_mult_206_n1006), .CO(DP_mult_206_n984), .S(DP_mult_206_n985) );
  FA_X1 DP_mult_206_U699 ( .A(DP_mult_206_n1004), .B(DP_mult_206_n987), .CI(
        DP_mult_206_n985), .CO(DP_mult_206_n982), .S(DP_mult_206_n983) );
  FA_X1 DP_mult_206_U698 ( .A(DP_mult_206_n1261), .B(DP_mult_206_n1349), .CI(
        DP_mult_206_n1239), .CO(DP_mult_206_n980), .S(DP_mult_206_n981) );
  FA_X1 DP_mult_206_U697 ( .A(DP_mult_206_n1460), .B(DP_mult_206_n1371), .CI(
        DP_mult_206_n1283), .CO(DP_mult_206_n978), .S(DP_mult_206_n979) );
  FA_X1 DP_mult_206_U696 ( .A(DP_mult_206_n1305), .B(DP_mult_206_n1327), .CI(
        DP_mult_206_n1437), .CO(DP_mult_206_n976), .S(DP_mult_206_n977) );
  FA_X1 DP_mult_206_U693 ( .A(DP_mult_206_n977), .B(DP_mult_206_n998), .CI(
        DP_mult_206_n979), .CO(DP_mult_206_n970), .S(DP_mult_206_n971) );
  FA_X1 DP_mult_206_U692 ( .A(DP_mult_206_n975), .B(DP_mult_206_n981), .CI(
        DP_mult_206_n992), .CO(DP_mult_206_n968), .S(DP_mult_206_n969) );
  FA_X1 DP_mult_206_U691 ( .A(DP_mult_206_n973), .B(DP_mult_206_n990), .CI(
        DP_mult_206_n988), .CO(DP_mult_206_n966), .S(DP_mult_206_n967) );
  FA_X1 DP_mult_206_U690 ( .A(DP_mult_206_n969), .B(DP_mult_206_n971), .CI(
        DP_mult_206_n986), .CO(DP_mult_206_n964), .S(DP_mult_206_n965) );
  FA_X1 DP_mult_206_U689 ( .A(DP_mult_206_n984), .B(DP_mult_206_n967), .CI(
        DP_mult_206_n965), .CO(DP_mult_206_n962), .S(DP_mult_206_n963) );
  HA_X1 DP_mult_206_U688 ( .A(DP_mult_206_n1238), .B(DP_mult_206_n1216), .CO(
        DP_mult_206_n960), .S(DP_mult_206_n961) );
  FA_X1 DP_mult_206_U684 ( .A(DP_mult_206_n1326), .B(DP_mult_206_n1392), .CI(
        DP_mult_206_n961), .CO(DP_mult_206_n952), .S(DP_mult_206_n953) );
  FA_X1 DP_mult_206_U683 ( .A(DP_mult_206_n976), .B(DP_mult_206_n980), .CI(
        DP_mult_206_n978), .CO(DP_mult_206_n950), .S(DP_mult_206_n951) );
  FA_X1 DP_mult_206_U682 ( .A(DP_mult_206_n955), .B(DP_mult_206_n974), .CI(
        DP_mult_206_n957), .CO(DP_mult_206_n948), .S(DP_mult_206_n949) );
  FA_X1 DP_mult_206_U681 ( .A(DP_mult_206_n972), .B(DP_mult_206_n959), .CI(
        DP_mult_206_n953), .CO(DP_mult_206_n946), .S(DP_mult_206_n947) );
  FA_X1 DP_mult_206_U680 ( .A(DP_mult_206_n951), .B(DP_mult_206_n970), .CI(
        DP_mult_206_n968), .CO(DP_mult_206_n944), .S(DP_mult_206_n945) );
  FA_X1 DP_mult_206_U679 ( .A(DP_mult_206_n947), .B(DP_mult_206_n949), .CI(
        DP_mult_206_n966), .CO(DP_mult_206_n942), .S(DP_mult_206_n943) );
  FA_X1 DP_mult_206_U678 ( .A(DP_mult_206_n964), .B(DP_mult_206_n945), .CI(
        DP_mult_206_n943), .CO(DP_mult_206_n940), .S(DP_mult_206_n941) );
  FA_X1 DP_mult_206_U675 ( .A(DP_mult_206_n1259), .B(DP_mult_206_n1347), .CI(
        DP_mult_206_n1303), .CO(DP_mult_206_n936), .S(DP_mult_206_n937) );
  FA_X1 DP_mult_206_U674 ( .A(DP_mult_206_n1281), .B(DP_mult_206_n1369), .CI(
        DP_mult_206_n1391), .CO(DP_mult_206_n934), .S(DP_mult_206_n935) );
  FA_X1 DP_mult_206_U672 ( .A(DP_mult_206_n1458), .B(DP_mult_206_n960), .CI(
        DP_mult_206_n939), .CO(DP_mult_206_n930), .S(DP_mult_206_n931) );
  FA_X1 DP_mult_206_U669 ( .A(DP_mult_206_n950), .B(DP_mult_206_n935), .CI(
        DP_mult_206_n931), .CO(DP_mult_206_n924), .S(DP_mult_206_n925) );
  FA_X1 DP_mult_206_U668 ( .A(DP_mult_206_n929), .B(DP_mult_206_n948), .CI(
        DP_mult_206_n946), .CO(DP_mult_206_n922), .S(DP_mult_206_n923) );
  FA_X1 DP_mult_206_U667 ( .A(DP_mult_206_n925), .B(DP_mult_206_n927), .CI(
        DP_mult_206_n944), .CO(DP_mult_206_n920), .S(DP_mult_206_n921) );
  FA_X1 DP_mult_206_U664 ( .A(DP_mult_206_n1214), .B(DP_mult_206_n1302), .CI(
        DP_mult_206_n917), .CO(DP_mult_206_n914), .S(DP_mult_206_n915) );
  FA_X1 DP_mult_206_U663 ( .A(DP_mult_206_n1236), .B(DP_mult_206_n1412), .CI(
        DP_mult_206_n1258), .CO(DP_mult_206_n912), .S(DP_mult_206_n913) );
  FA_X1 DP_mult_206_U662 ( .A(DP_mult_206_n1346), .B(DP_mult_206_n1324), .CI(
        DP_mult_206_n1280), .CO(DP_mult_206_n910), .S(DP_mult_206_n911) );
  FA_X1 DP_mult_206_U660 ( .A(DP_mult_206_n932), .B(DP_mult_206_n936), .CI(
        DP_mult_206_n934), .CO(DP_mult_206_n906), .S(DP_mult_206_n907) );
  FA_X1 DP_mult_206_U659 ( .A(DP_mult_206_n911), .B(DP_mult_206_n913), .CI(
        DP_mult_206_n915), .CO(DP_mult_206_n904), .S(DP_mult_206_n905) );
  FA_X1 DP_mult_206_U658 ( .A(DP_mult_206_n909), .B(DP_mult_206_n930), .CI(
        DP_mult_206_n928), .CO(DP_mult_206_n902), .S(DP_mult_206_n903) );
  FA_X1 DP_mult_206_U657 ( .A(DP_mult_206_n907), .B(DP_mult_206_n926), .CI(
        DP_mult_206_n905), .CO(DP_mult_206_n900), .S(DP_mult_206_n901) );
  FA_X1 DP_mult_206_U654 ( .A(DP_mult_206_n1235), .B(DP_mult_206_n1213), .CI(
        DP_mult_206_n1411), .CO(DP_mult_206_n894), .S(DP_mult_206_n895) );
  FA_X1 DP_mult_206_U653 ( .A(DP_mult_206_n2050), .B(DP_mult_206_n1323), .CI(
        DP_mult_206_n1279), .CO(DP_mult_206_n892), .S(DP_mult_206_n893) );
  FA_X1 DP_mult_206_U652 ( .A(DP_mult_206_n1257), .B(DP_mult_206_n1301), .CI(
        DP_mult_206_n1345), .CO(DP_mult_206_n890), .S(DP_mult_206_n891) );
  FA_X1 DP_mult_206_U651 ( .A(DP_mult_206_n1367), .B(DP_mult_206_n1389), .CI(
        DP_mult_206_n1434), .CO(DP_mult_206_n888), .S(DP_mult_206_n889) );
  FA_X1 DP_mult_206_U650 ( .A(DP_mult_206_n910), .B(DP_mult_206_n912), .CI(
        DP_mult_206_n914), .CO(DP_mult_206_n886), .S(DP_mult_206_n887) );
  FA_X1 DP_mult_206_U647 ( .A(DP_mult_206_n887), .B(DP_mult_206_n904), .CI(
        DP_mult_206_n902), .CO(DP_mult_206_n880), .S(DP_mult_206_n881) );
  FA_X1 DP_mult_206_U646 ( .A(DP_mult_206_n883), .B(DP_mult_206_n885), .CI(
        DP_mult_206_n900), .CO(DP_mult_206_n878), .S(DP_mult_206_n879) );
  FA_X1 DP_mult_206_U645 ( .A(DP_mult_206_n898), .B(DP_mult_206_n881), .CI(
        DP_mult_206_n879), .CO(DP_mult_206_n876), .S(DP_mult_206_n877) );
  FA_X1 DP_mult_206_U643 ( .A(DP_mult_206_n1388), .B(DP_mult_206_n1278), .CI(
        DP_mult_206_n875), .CO(DP_mult_206_n872), .S(DP_mult_206_n873) );
  FA_X1 DP_mult_206_U642 ( .A(DP_mult_206_n1366), .B(DP_mult_206_n1212), .CI(
        DP_mult_206_n1344), .CO(DP_mult_206_n870), .S(DP_mult_206_n871) );
  FA_X1 DP_mult_206_U641 ( .A(DP_mult_206_n1234), .B(DP_mult_206_n1322), .CI(
        DP_mult_206_n1256), .CO(DP_mult_206_n868), .S(DP_mult_206_n869) );
  FA_X1 DP_mult_206_U640 ( .A(DP_mult_206_n1300), .B(DP_mult_206_n894), .CI(
        DP_mult_206_n892), .CO(DP_mult_206_n866), .S(DP_mult_206_n867) );
  FA_X1 DP_mult_206_U639 ( .A(DP_mult_206_n890), .B(DP_mult_206_n869), .CI(
        DP_mult_206_n871), .CO(DP_mult_206_n864), .S(DP_mult_206_n865) );
  FA_X1 DP_mult_206_U637 ( .A(DP_mult_206_n867), .B(DP_mult_206_n884), .CI(
        DP_mult_206_n865), .CO(DP_mult_206_n860), .S(DP_mult_206_n861) );
  FA_X1 DP_mult_206_U636 ( .A(DP_mult_206_n863), .B(DP_mult_206_n882), .CI(
        DP_mult_206_n880), .CO(DP_mult_206_n858), .S(DP_mult_206_n859) );
  FA_X1 DP_mult_206_U635 ( .A(DP_mult_206_n878), .B(DP_mult_206_n861), .CI(
        DP_mult_206_n859), .CO(DP_mult_206_n856), .S(DP_mult_206_n857) );
  FA_X1 DP_mult_206_U634 ( .A(DP_mult_206_n1387), .B(DP_mult_206_n1233), .CI(
        DP_mult_206_n1211), .CO(DP_mult_206_n854), .S(DP_mult_206_n855) );
  FA_X1 DP_mult_206_U633 ( .A(DP_mult_206_n1255), .B(DP_mult_206_n1321), .CI(
        DP_mult_206_n874), .CO(DP_mult_206_n852), .S(DP_mult_206_n853) );
  FA_X1 DP_mult_206_U632 ( .A(DP_mult_206_n1277), .B(DP_mult_206_n1343), .CI(
        DP_mult_206_n1299), .CO(DP_mult_206_n850), .S(DP_mult_206_n851) );
  FA_X1 DP_mult_206_U629 ( .A(DP_mult_206_n855), .B(DP_mult_206_n853), .CI(
        DP_mult_206_n866), .CO(DP_mult_206_n844), .S(DP_mult_206_n845) );
  FA_X1 DP_mult_206_U627 ( .A(DP_mult_206_n845), .B(DP_mult_206_n847), .CI(
        DP_mult_206_n860), .CO(DP_mult_206_n840), .S(DP_mult_206_n841) );
  FA_X1 DP_mult_206_U626 ( .A(DP_mult_206_n858), .B(DP_mult_206_n843), .CI(
        DP_mult_206_n841), .CO(DP_mult_206_n838), .S(DP_mult_206_n839) );
  FA_X1 DP_mult_206_U623 ( .A(DP_mult_206_n1232), .B(DP_mult_206_n1364), .CI(
        DP_mult_206_n1342), .CO(DP_mult_206_n832), .S(DP_mult_206_n833) );
  FA_X1 DP_mult_206_U621 ( .A(DP_mult_206_n850), .B(DP_mult_206_n854), .CI(
        DP_mult_206_n852), .CO(DP_mult_206_n828), .S(DP_mult_206_n829) );
  FA_X1 DP_mult_206_U620 ( .A(DP_mult_206_n835), .B(DP_mult_206_n831), .CI(
        DP_mult_206_n833), .CO(DP_mult_206_n826), .S(DP_mult_206_n827) );
  FA_X1 DP_mult_206_U617 ( .A(DP_mult_206_n840), .B(DP_mult_206_n825), .CI(
        DP_mult_206_n823), .CO(DP_mult_206_n820), .S(DP_mult_206_n821) );
  FA_X1 DP_mult_206_U615 ( .A(DP_mult_206_n1231), .B(DP_mult_206_n1297), .CI(
        DP_mult_206_n1275), .CO(DP_mult_206_n816), .S(DP_mult_206_n817) );
  FA_X1 DP_mult_206_U614 ( .A(DP_mult_206_n1319), .B(DP_mult_206_n1253), .CI(
        DP_mult_206_n1341), .CO(DP_mult_206_n814), .S(DP_mult_206_n815) );
  FA_X1 DP_mult_206_U613 ( .A(DP_mult_206_n1386), .B(DP_mult_206_n830), .CI(
        DP_mult_206_n834), .CO(DP_mult_206_n812), .S(DP_mult_206_n813) );
  FA_X1 DP_mult_206_U612 ( .A(DP_mult_206_n815), .B(DP_mult_206_n832), .CI(
        DP_mult_206_n817), .CO(DP_mult_206_n810), .S(DP_mult_206_n811) );
  FA_X1 DP_mult_206_U610 ( .A(DP_mult_206_n811), .B(DP_mult_206_n826), .CI(
        DP_mult_206_n824), .CO(DP_mult_206_n806), .S(DP_mult_206_n807) );
  FA_X1 DP_mult_206_U609 ( .A(DP_mult_206_n822), .B(DP_mult_206_n809), .CI(
        DP_mult_206_n807), .CO(DP_mult_206_n804), .S(DP_mult_206_n805) );
  FA_X1 DP_mult_206_U607 ( .A(DP_mult_206_n1340), .B(DP_mult_206_n1252), .CI(
        DP_mult_206_n803), .CO(DP_mult_206_n800), .S(DP_mult_206_n801) );
  FA_X1 DP_mult_206_U606 ( .A(DP_mult_206_n1208), .B(DP_mult_206_n1318), .CI(
        DP_mult_206_n1230), .CO(DP_mult_206_n798), .S(DP_mult_206_n799) );
  FA_X1 DP_mult_206_U604 ( .A(DP_mult_206_n814), .B(DP_mult_206_n816), .CI(
        DP_mult_206_n799), .CO(DP_mult_206_n794), .S(DP_mult_206_n795) );
  FA_X1 DP_mult_206_U603 ( .A(DP_mult_206_n797), .B(DP_mult_206_n801), .CI(
        DP_mult_206_n812), .CO(DP_mult_206_n792), .S(DP_mult_206_n793) );
  FA_X1 DP_mult_206_U601 ( .A(DP_mult_206_n806), .B(DP_mult_206_n793), .CI(
        DP_mult_206_n791), .CO(DP_mult_206_n788), .S(DP_mult_206_n789) );
  FA_X1 DP_mult_206_U600 ( .A(DP_mult_206_n1251), .B(DP_mult_206_n1207), .CI(
        DP_mult_206_n802), .CO(DP_mult_206_n786), .S(DP_mult_206_n787) );
  FA_X1 DP_mult_206_U599 ( .A(DP_mult_206_n1273), .B(DP_mult_206_n1317), .CI(
        DP_mult_206_n1295), .CO(DP_mult_206_n784), .S(DP_mult_206_n785) );
  FA_X1 DP_mult_206_U598 ( .A(DP_mult_206_n1339), .B(DP_mult_206_n1229), .CI(
        DP_mult_206_n1362), .CO(DP_mult_206_n782), .S(DP_mult_206_n783) );
  FA_X1 DP_mult_206_U597 ( .A(DP_mult_206_n798), .B(DP_mult_206_n800), .CI(
        DP_mult_206_n785), .CO(DP_mult_206_n780), .S(DP_mult_206_n781) );
  FA_X1 DP_mult_206_U596 ( .A(DP_mult_206_n783), .B(DP_mult_206_n787), .CI(
        DP_mult_206_n796), .CO(DP_mult_206_n778), .S(DP_mult_206_n779) );
  FA_X1 DP_mult_206_U595 ( .A(DP_mult_206_n781), .B(DP_mult_206_n794), .CI(
        DP_mult_206_n792), .CO(DP_mult_206_n776), .S(DP_mult_206_n777) );
  FA_X1 DP_mult_206_U594 ( .A(DP_mult_206_n790), .B(DP_mult_206_n779), .CI(
        DP_mult_206_n777), .CO(DP_mult_206_n774), .S(DP_mult_206_n775) );
  FA_X1 DP_mult_206_U592 ( .A(DP_mult_206_n1316), .B(DP_mult_206_n1250), .CI(
        DP_mult_206_n773), .CO(DP_mult_206_n770), .S(DP_mult_206_n771) );
  FA_X1 DP_mult_206_U591 ( .A(DP_mult_206_n1294), .B(DP_mult_206_n1206), .CI(
        DP_mult_206_n1272), .CO(DP_mult_206_n768), .S(DP_mult_206_n769) );
  FA_X1 DP_mult_206_U590 ( .A(DP_mult_206_n786), .B(DP_mult_206_n1228), .CI(
        DP_mult_206_n784), .CO(DP_mult_206_n766), .S(DP_mult_206_n767) );
  FA_X1 DP_mult_206_U589 ( .A(DP_mult_206_n771), .B(DP_mult_206_n769), .CI(
        DP_mult_206_n782), .CO(DP_mult_206_n764), .S(DP_mult_206_n765) );
  FA_X1 DP_mult_206_U588 ( .A(DP_mult_206_n767), .B(DP_mult_206_n780), .CI(
        DP_mult_206_n778), .CO(DP_mult_206_n762), .S(DP_mult_206_n763) );
  FA_X1 DP_mult_206_U587 ( .A(DP_mult_206_n776), .B(DP_mult_206_n765), .CI(
        DP_mult_206_n763), .CO(DP_mult_206_n760), .S(DP_mult_206_n761) );
  FA_X1 DP_mult_206_U586 ( .A(DP_mult_206_n772), .B(DP_mult_206_n1205), .CI(
        DP_mult_206_n1227), .CO(DP_mult_206_n758), .S(DP_mult_206_n759) );
  FA_X1 DP_mult_206_U585 ( .A(DP_mult_206_n1249), .B(DP_mult_206_n1293), .CI(
        DP_mult_206_n1315), .CO(DP_mult_206_n756), .S(DP_mult_206_n757) );
  FA_X1 DP_mult_206_U584 ( .A(DP_mult_206_n1338), .B(DP_mult_206_n1271), .CI(
        DP_mult_206_n770), .CO(DP_mult_206_n754), .S(DP_mult_206_n755) );
  FA_X1 DP_mult_206_U583 ( .A(DP_mult_206_n757), .B(DP_mult_206_n768), .CI(
        DP_mult_206_n759), .CO(DP_mult_206_n752), .S(DP_mult_206_n753) );
  FA_X1 DP_mult_206_U582 ( .A(DP_mult_206_n755), .B(DP_mult_206_n766), .CI(
        DP_mult_206_n764), .CO(DP_mult_206_n750), .S(DP_mult_206_n751) );
  FA_X1 DP_mult_206_U581 ( .A(DP_mult_206_n762), .B(DP_mult_206_n753), .CI(
        DP_mult_206_n751), .CO(DP_mult_206_n748), .S(DP_mult_206_n749) );
  FA_X1 DP_mult_206_U579 ( .A(DP_mult_206_n1292), .B(DP_mult_206_n1248), .CI(
        DP_mult_206_n747), .CO(DP_mult_206_n744), .S(DP_mult_206_n745) );
  FA_X1 DP_mult_206_U578 ( .A(DP_mult_206_n1226), .B(DP_mult_206_n1204), .CI(
        DP_mult_206_n1270), .CO(DP_mult_206_n742), .S(DP_mult_206_n743) );
  FA_X1 DP_mult_206_U577 ( .A(DP_mult_206_n756), .B(DP_mult_206_n758), .CI(
        DP_mult_206_n743), .CO(DP_mult_206_n740), .S(DP_mult_206_n741) );
  FA_X1 DP_mult_206_U576 ( .A(DP_mult_206_n754), .B(DP_mult_206_n745), .CI(
        DP_mult_206_n752), .CO(DP_mult_206_n738), .S(DP_mult_206_n739) );
  FA_X1 DP_mult_206_U575 ( .A(DP_mult_206_n750), .B(DP_mult_206_n741), .CI(
        DP_mult_206_n739), .CO(DP_mult_206_n736), .S(DP_mult_206_n737) );
  FA_X1 DP_mult_206_U574 ( .A(DP_mult_206_n746), .B(DP_mult_206_n1203), .CI(
        DP_mult_206_n1247), .CO(DP_mult_206_n734), .S(DP_mult_206_n735) );
  FA_X1 DP_mult_206_U573 ( .A(DP_mult_206_n1225), .B(DP_mult_206_n1291), .CI(
        DP_mult_206_n1269), .CO(DP_mult_206_n732), .S(DP_mult_206_n733) );
  FA_X1 DP_mult_206_U572 ( .A(DP_mult_206_n744), .B(DP_mult_206_n1314), .CI(
        DP_mult_206_n742), .CO(DP_mult_206_n730), .S(DP_mult_206_n731) );
  FA_X1 DP_mult_206_U571 ( .A(DP_mult_206_n735), .B(DP_mult_206_n733), .CI(
        DP_mult_206_n740), .CO(DP_mult_206_n728), .S(DP_mult_206_n729) );
  FA_X1 DP_mult_206_U570 ( .A(DP_mult_206_n738), .B(DP_mult_206_n731), .CI(
        DP_mult_206_n729), .CO(DP_mult_206_n726), .S(DP_mult_206_n727) );
  FA_X1 DP_mult_206_U568 ( .A(DP_mult_206_n1268), .B(DP_mult_206_n1224), .CI(
        DP_mult_206_n725), .CO(DP_mult_206_n722), .S(DP_mult_206_n723) );
  FA_X1 DP_mult_206_U567 ( .A(DP_mult_206_n1202), .B(DP_mult_206_n1246), .CI(
        DP_mult_206_n734), .CO(DP_mult_206_n720), .S(DP_mult_206_n721) );
  FA_X1 DP_mult_206_U566 ( .A(DP_mult_206_n723), .B(DP_mult_206_n732), .CI(
        DP_mult_206_n730), .CO(DP_mult_206_n718), .S(DP_mult_206_n719) );
  FA_X1 DP_mult_206_U565 ( .A(DP_mult_206_n728), .B(DP_mult_206_n721), .CI(
        DP_mult_206_n719), .CO(DP_mult_206_n716), .S(DP_mult_206_n717) );
  FA_X1 DP_mult_206_U564 ( .A(DP_mult_206_n1267), .B(DP_mult_206_n1201), .CI(
        DP_mult_206_n724), .CO(DP_mult_206_n714), .S(DP_mult_206_n715) );
  FA_X1 DP_mult_206_U563 ( .A(DP_mult_206_n1245), .B(DP_mult_206_n1223), .CI(
        DP_mult_206_n1290), .CO(DP_mult_206_n712), .S(DP_mult_206_n713) );
  FA_X1 DP_mult_206_U562 ( .A(DP_mult_206_n715), .B(DP_mult_206_n722), .CI(
        DP_mult_206_n720), .CO(DP_mult_206_n710), .S(DP_mult_206_n711) );
  FA_X1 DP_mult_206_U561 ( .A(DP_mult_206_n718), .B(DP_mult_206_n713), .CI(
        DP_mult_206_n711), .CO(DP_mult_206_n708), .S(DP_mult_206_n709) );
  FA_X1 DP_mult_206_U559 ( .A(DP_mult_206_n1222), .B(DP_mult_206_n1200), .CI(
        DP_mult_206_n707), .CO(DP_mult_206_n704), .S(DP_mult_206_n705) );
  FA_X1 DP_mult_206_U558 ( .A(DP_mult_206_n714), .B(DP_mult_206_n1244), .CI(
        DP_mult_206_n705), .CO(DP_mult_206_n702), .S(DP_mult_206_n703) );
  FA_X1 DP_mult_206_U557 ( .A(DP_mult_206_n710), .B(DP_mult_206_n712), .CI(
        DP_mult_206_n703), .CO(DP_mult_206_n700), .S(DP_mult_206_n701) );
  FA_X1 DP_mult_206_U556 ( .A(DP_mult_206_n1221), .B(DP_mult_206_n1199), .CI(
        DP_mult_206_n706), .CO(DP_mult_206_n698), .S(DP_mult_206_n699) );
  FA_X1 DP_mult_206_U555 ( .A(DP_mult_206_n1266), .B(DP_mult_206_n1243), .CI(
        DP_mult_206_n704), .CO(DP_mult_206_n696), .S(DP_mult_206_n697) );
  FA_X1 DP_mult_206_U554 ( .A(DP_mult_206_n702), .B(DP_mult_206_n699), .CI(
        DP_mult_206_n697), .CO(DP_mult_206_n694), .S(DP_mult_206_n695) );
  FA_X1 DP_mult_206_U552 ( .A(DP_mult_206_n1198), .B(DP_mult_206_n1220), .CI(
        DP_mult_206_n693), .CO(DP_mult_206_n690), .S(DP_mult_206_n691) );
  FA_X1 DP_mult_206_U551 ( .A(DP_mult_206_n691), .B(DP_mult_206_n698), .CI(
        DP_mult_206_n696), .CO(DP_mult_206_n688), .S(DP_mult_206_n689) );
  FA_X1 DP_mult_206_U550 ( .A(DP_mult_206_n1219), .B(DP_mult_206_n692), .CI(
        DP_mult_206_n1197), .CO(DP_mult_206_n686), .S(DP_mult_206_n687) );
  FA_X1 DP_mult_206_U549 ( .A(DP_mult_206_n690), .B(DP_mult_206_n1242), .CI(
        DP_mult_206_n687), .CO(DP_mult_206_n684), .S(DP_mult_206_n685) );
  FA_X1 DP_mult_206_U547 ( .A(DP_mult_206_n683), .B(DP_mult_206_n1196), .CI(
        DP_mult_206_n686), .CO(DP_mult_206_n680), .S(DP_mult_206_n681) );
  FA_X1 DP_mult_206_U546 ( .A(DP_mult_206_n1195), .B(DP_mult_206_n682), .CI(
        DP_mult_206_n1218), .CO(DP_mult_206_n678), .S(DP_mult_206_n679) );
  INV_X1 DP_mult_207_U2807 ( .A(DP_coeffs_ff_int[26]), .ZN(DP_mult_207_n2316)
         );
  INV_X1 DP_mult_207_U2806 ( .A(DP_coeffs_ff_int[26]), .ZN(DP_mult_207_n2315)
         );
  INV_X1 DP_mult_207_U2805 ( .A(DP_mult_207_n2316), .ZN(DP_mult_207_n2314) );
  INV_X1 DP_mult_207_U2804 ( .A(DP_coeffs_ff_int[28]), .ZN(DP_mult_207_n2310)
         );
  INV_X1 DP_mult_207_U2803 ( .A(DP_mult_207_n2310), .ZN(DP_mult_207_n2309) );
  INV_X1 DP_mult_207_U2802 ( .A(DP_mult_207_n1939), .ZN(DP_mult_207_n2306) );
  INV_X1 DP_mult_207_U2801 ( .A(DP_coeffs_ff_int[30]), .ZN(DP_mult_207_n2305)
         );
  INV_X1 DP_mult_207_U2800 ( .A(DP_mult_207_n2306), .ZN(DP_mult_207_n2304) );
  INV_X1 DP_mult_207_U2799 ( .A(DP_coeffs_ff_int[32]), .ZN(DP_mult_207_n2302)
         );
  INV_X1 DP_mult_207_U2798 ( .A(DP_coeffs_ff_int[32]), .ZN(DP_mult_207_n2301)
         );
  INV_X1 DP_mult_207_U2797 ( .A(DP_mult_207_n2302), .ZN(DP_mult_207_n2300) );
  INV_X1 DP_mult_207_U2796 ( .A(DP_coeffs_ff_int[34]), .ZN(DP_mult_207_n2297)
         );
  INV_X1 DP_mult_207_U2795 ( .A(DP_coeffs_ff_int[34]), .ZN(DP_mult_207_n2296)
         );
  INV_X1 DP_mult_207_U2794 ( .A(DP_mult_207_n2297), .ZN(DP_mult_207_n2295) );
  INV_X1 DP_mult_207_U2793 ( .A(DP_coeffs_ff_int[36]), .ZN(DP_mult_207_n2292)
         );
  INV_X1 DP_mult_207_U2792 ( .A(DP_coeffs_ff_int[36]), .ZN(DP_mult_207_n2291)
         );
  INV_X1 DP_mult_207_U2791 ( .A(DP_mult_207_n2292), .ZN(DP_mult_207_n2290) );
  INV_X1 DP_mult_207_U2790 ( .A(DP_coeffs_ff_int[38]), .ZN(DP_mult_207_n2289)
         );
  INV_X1 DP_mult_207_U2789 ( .A(DP_coeffs_ff_int[38]), .ZN(DP_mult_207_n2288)
         );
  INV_X1 DP_mult_207_U2788 ( .A(DP_mult_207_n2288), .ZN(DP_mult_207_n2287) );
  INV_X1 DP_mult_207_U2787 ( .A(DP_coeffs_ff_int[40]), .ZN(DP_mult_207_n2284)
         );
  INV_X1 DP_mult_207_U2786 ( .A(DP_coeffs_ff_int[40]), .ZN(DP_mult_207_n2283)
         );
  INV_X1 DP_mult_207_U2785 ( .A(DP_mult_207_n2284), .ZN(DP_mult_207_n2282) );
  INV_X1 DP_mult_207_U2784 ( .A(DP_coeffs_ff_int[42]), .ZN(DP_mult_207_n2279)
         );
  INV_X1 DP_mult_207_U2783 ( .A(DP_coeffs_ff_int[42]), .ZN(DP_mult_207_n2278)
         );
  INV_X1 DP_mult_207_U2782 ( .A(DP_mult_207_n2279), .ZN(DP_mult_207_n2277) );
  INV_X1 DP_mult_207_U2781 ( .A(DP_coeffs_ff_int[44]), .ZN(DP_mult_207_n2274)
         );
  INV_X1 DP_mult_207_U2780 ( .A(DP_coeffs_ff_int[44]), .ZN(DP_mult_207_n2273)
         );
  INV_X1 DP_mult_207_U2779 ( .A(DP_mult_207_n2274), .ZN(DP_mult_207_n2272) );
  INV_X1 DP_mult_207_U2778 ( .A(DP_coeffs_ff_int[46]), .ZN(DP_mult_207_n2268)
         );
  INV_X1 DP_mult_207_U2777 ( .A(DP_coeffs_ff_int[46]), .ZN(DP_mult_207_n2267)
         );
  INV_X1 DP_mult_207_U2776 ( .A(DP_mult_207_n2268), .ZN(DP_mult_207_n2266) );
  INV_X1 DP_mult_207_U2775 ( .A(DP_mult_207_n2084), .ZN(DP_mult_207_n2260) );
  INV_X1 DP_mult_207_U2774 ( .A(DP_mult_207_n2082), .ZN(DP_mult_207_n2256) );
  INV_X1 DP_mult_207_U2773 ( .A(DP_mult_207_n2254), .ZN(DP_mult_207_n2253) );
  INV_X2 DP_mult_207_U2772 ( .A(DP_mult_207_n2274), .ZN(DP_mult_207_n2271) );
  INV_X2 DP_mult_207_U2771 ( .A(DP_mult_207_n2187), .ZN(DP_mult_207_n2220) );
  XNOR2_X1 DP_mult_207_U2770 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1713) );
  XNOR2_X1 DP_mult_207_U2769 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1711) );
  XNOR2_X1 DP_mult_207_U2768 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1719) );
  XNOR2_X1 DP_mult_207_U2767 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1715) );
  XNOR2_X1 DP_mult_207_U2766 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1709) );
  OAI22_X1 DP_mult_207_U2765 ( .A1(DP_mult_207_n2230), .A2(DP_mult_207_n1683), 
        .B1(DP_mult_207_n1682), .B2(DP_mult_207_n2256), .ZN(DP_mult_207_n836)
         );
  XNOR2_X1 DP_mult_207_U2764 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1717) );
  OAI22_X1 DP_mult_207_U2763 ( .A1(DP_mult_207_n2229), .A2(DP_mult_207_n1693), 
        .B1(DP_mult_207_n1692), .B2(DP_mult_207_n2255), .ZN(DP_mult_207_n1396)
         );
  OAI22_X1 DP_mult_207_U2762 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n2283), 
        .B1(DP_mult_207_n1706), .B2(DP_mult_207_n2255), .ZN(DP_mult_207_n1190)
         );
  OAI22_X1 DP_mult_207_U2761 ( .A1(DP_mult_207_n2196), .A2(DP_mult_207_n1684), 
        .B1(DP_mult_207_n2255), .B2(DP_mult_207_n1683), .ZN(DP_mult_207_n1387)
         );
  INV_X1 DP_mult_207_U2760 ( .A(DP_mult_207_n836), .ZN(DP_mult_207_n837) );
  OAI22_X1 DP_mult_207_U2759 ( .A1(DP_mult_207_n2196), .A2(DP_mult_207_n1688), 
        .B1(DP_mult_207_n1958), .B2(DP_mult_207_n1687), .ZN(DP_mult_207_n1391)
         );
  OAI22_X1 DP_mult_207_U2758 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1685), 
        .B1(DP_mult_207_n1684), .B2(DP_mult_207_n2255), .ZN(DP_mult_207_n1388)
         );
  OAI22_X1 DP_mult_207_U2757 ( .A1(DP_mult_207_n2229), .A2(DP_mult_207_n1692), 
        .B1(DP_mult_207_n2256), .B2(DP_mult_207_n1691), .ZN(DP_mult_207_n1395)
         );
  OAI22_X1 DP_mult_207_U2756 ( .A1(DP_mult_207_n2196), .A2(DP_mult_207_n1687), 
        .B1(DP_mult_207_n1686), .B2(DP_mult_207_n2256), .ZN(DP_mult_207_n1390)
         );
  OAI22_X1 DP_mult_207_U2755 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1690), 
        .B1(DP_mult_207_n2255), .B2(DP_mult_207_n1689), .ZN(DP_mult_207_n1393)
         );
  OAI22_X1 DP_mult_207_U2754 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1689), 
        .B1(DP_mult_207_n1688), .B2(DP_mult_207_n2256), .ZN(DP_mult_207_n1392)
         );
  OAI22_X1 DP_mult_207_U2753 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1686), 
        .B1(DP_mult_207_n2255), .B2(DP_mult_207_n1685), .ZN(DP_mult_207_n1389)
         );
  OAI22_X1 DP_mult_207_U2752 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1691), 
        .B1(DP_mult_207_n1690), .B2(DP_mult_207_n2255), .ZN(DP_mult_207_n1394)
         );
  NAND2_X1 DP_mult_207_U2751 ( .A1(DP_mult_207_n775), .A2(DP_mult_207_n788), 
        .ZN(DP_mult_207_n474) );
  OAI21_X1 DP_mult_207_U2750 ( .B1(DP_mult_207_n2104), .B2(DP_mult_207_n398), 
        .A(DP_mult_207_n399), .ZN(DP_mult_207_n397) );
  OAI21_X1 DP_mult_207_U2749 ( .B1(DP_mult_207_n2104), .B2(DP_mult_207_n389), 
        .A(DP_mult_207_n390), .ZN(DP_mult_207_n388) );
  OAI21_X1 DP_mult_207_U2748 ( .B1(DP_mult_207_n2103), .B2(DP_mult_207_n431), 
        .A(DP_mult_207_n432), .ZN(DP_mult_207_n430) );
  OAI21_X1 DP_mult_207_U2747 ( .B1(DP_mult_207_n2212), .B2(DP_mult_207_n411), 
        .A(DP_mult_207_n412), .ZN(DP_mult_207_n410) );
  OAI21_X1 DP_mult_207_U2746 ( .B1(DP_mult_207_n301), .B2(DP_mult_207_n420), 
        .A(DP_mult_207_n421), .ZN(DP_mult_207_n419) );
  OAI21_X1 DP_mult_207_U2745 ( .B1(DP_mult_207_n2103), .B2(DP_mult_207_n343), 
        .A(DP_mult_207_n344), .ZN(DP_mult_207_n342) );
  OAI21_X1 DP_mult_207_U2744 ( .B1(DP_mult_207_n2212), .B2(DP_mult_207_n380), 
        .A(DP_mult_207_n381), .ZN(DP_mult_207_n379) );
  OAI21_X1 DP_mult_207_U2743 ( .B1(DP_mult_207_n2103), .B2(DP_mult_207_n371), 
        .A(DP_mult_207_n372), .ZN(DP_mult_207_n370) );
  OAI21_X1 DP_mult_207_U2742 ( .B1(DP_mult_207_n2104), .B2(DP_mult_207_n354), 
        .A(DP_mult_207_n355), .ZN(DP_mult_207_n353) );
  OAI21_X1 DP_mult_207_U2741 ( .B1(DP_mult_207_n301), .B2(DP_mult_207_n438), 
        .A(DP_mult_207_n439), .ZN(DP_mult_207_n437) );
  OAI21_X1 DP_mult_207_U2740 ( .B1(DP_mult_207_n301), .B2(DP_mult_207_n326), 
        .A(DP_mult_207_n327), .ZN(DP_mult_207_n325) );
  XNOR2_X1 DP_mult_207_U2739 ( .A(DP_mult_207_n437), .B(DP_mult_207_n311), 
        .ZN(DP_pipe0_coeff_pipe01[13]) );
  XNOR2_X1 DP_mult_207_U2738 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1584) );
  XNOR2_X1 DP_mult_207_U2737 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1586) );
  XNOR2_X1 DP_mult_207_U2736 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1594) );
  OAI22_X1 DP_mult_207_U2735 ( .A1(DP_mult_207_n2144), .A2(DP_mult_207_n1558), 
        .B1(DP_mult_207_n1557), .B2(DP_mult_207_n2008), .ZN(DP_mult_207_n706)
         );
  XNOR2_X1 DP_mult_207_U2734 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1590) );
  XNOR2_X1 DP_mult_207_U2733 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1592) );
  XNOR2_X1 DP_mult_207_U2732 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1588) );
  OAI22_X1 DP_mult_207_U2731 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1562), 
        .B1(DP_mult_207_n1561), .B2(DP_mult_207_n2008), .ZN(DP_mult_207_n1270)
         );
  OAI22_X1 DP_mult_207_U2730 ( .A1(DP_mult_207_n2219), .A2(DP_mult_207_n1568), 
        .B1(DP_mult_207_n1567), .B2(DP_mult_207_n2241), .ZN(DP_mult_207_n1276)
         );
  OAI22_X1 DP_mult_207_U2729 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n2305), 
        .B1(DP_mult_207_n1581), .B2(DP_mult_207_n2008), .ZN(DP_mult_207_n1185)
         );
  OAI22_X1 DP_mult_207_U2728 ( .A1(DP_mult_207_n2144), .A2(DP_mult_207_n1559), 
        .B1(DP_mult_207_n2008), .B2(DP_mult_207_n1558), .ZN(DP_mult_207_n1267)
         );
  OAI22_X1 DP_mult_207_U2727 ( .A1(DP_mult_207_n2144), .A2(DP_mult_207_n1560), 
        .B1(DP_mult_207_n1559), .B2(DP_mult_207_n2241), .ZN(DP_mult_207_n1268)
         );
  OAI22_X1 DP_mult_207_U2726 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1565), 
        .B1(DP_mult_207_n2241), .B2(DP_mult_207_n1564), .ZN(DP_mult_207_n1273)
         );
  OAI22_X1 DP_mult_207_U2725 ( .A1(DP_mult_207_n2144), .A2(DP_mult_207_n1561), 
        .B1(DP_mult_207_n2008), .B2(DP_mult_207_n1560), .ZN(DP_mult_207_n1269)
         );
  OAI22_X1 DP_mult_207_U2724 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1564), 
        .B1(DP_mult_207_n1563), .B2(DP_mult_207_n2241), .ZN(DP_mult_207_n1272)
         );
  OAI22_X1 DP_mult_207_U2723 ( .A1(DP_mult_207_n2144), .A2(DP_mult_207_n1566), 
        .B1(DP_mult_207_n1565), .B2(DP_mult_207_n2008), .ZN(DP_mult_207_n1274)
         );
  OAI22_X1 DP_mult_207_U2722 ( .A1(DP_mult_207_n2144), .A2(DP_mult_207_n1567), 
        .B1(DP_mult_207_n2241), .B2(DP_mult_207_n1566), .ZN(DP_mult_207_n1275)
         );
  OAI22_X1 DP_mult_207_U2721 ( .A1(DP_mult_207_n2144), .A2(DP_mult_207_n1563), 
        .B1(DP_mult_207_n2008), .B2(DP_mult_207_n1562), .ZN(DP_mult_207_n1271)
         );
  NAND2_X1 DP_mult_207_U2720 ( .A1(DP_mult_207_n694), .A2(DP_mult_207_n689), 
        .ZN(DP_mult_207_n378) );
  NAND2_X1 DP_mult_207_U2719 ( .A1(DP_mult_207_n2178), .A2(DP_mult_207_n2180), 
        .ZN(DP_mult_207_n364) );
  NAND2_X1 DP_mult_207_U2718 ( .A1(DP_mult_207_n382), .A2(DP_mult_207_n2178), 
        .ZN(DP_mult_207_n371) );
  AOI21_X1 DP_mult_207_U2717 ( .B1(DP_mult_207_n383), .B2(DP_mult_207_n2178), 
        .A(DP_mult_207_n376), .ZN(DP_mult_207_n372) );
  NAND2_X1 DP_mult_207_U2716 ( .A1(DP_mult_207_n2178), .A2(DP_mult_207_n378), 
        .ZN(DP_mult_207_n305) );
  INV_X1 DP_mult_207_U2715 ( .A(DP_mult_207_n325), .ZN(
        DP_pipe0_coeff_pipe01[23]) );
  XNOR2_X1 DP_mult_207_U2714 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1742) );
  XNOR2_X1 DP_mult_207_U2713 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1738) );
  XNOR2_X1 DP_mult_207_U2712 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1744) );
  XNOR2_X1 DP_mult_207_U2711 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1736) );
  XNOR2_X1 DP_mult_207_U2710 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1740) );
  OAI22_X1 DP_mult_207_U2709 ( .A1(DP_mult_207_n2231), .A2(DP_mult_207_n1724), 
        .B1(DP_mult_207_n1723), .B2(DP_mult_207_n2258), .ZN(DP_mult_207_n1426)
         );
  XNOR2_X1 DP_mult_207_U2708 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1734) );
  OAI22_X1 DP_mult_207_U2707 ( .A1(DP_mult_207_n2232), .A2(DP_mult_207_n1714), 
        .B1(DP_mult_207_n1713), .B2(DP_mult_207_n2257), .ZN(DP_mult_207_n1416)
         );
  OAI22_X1 DP_mult_207_U2706 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1719), 
        .B1(DP_mult_207_n2257), .B2(DP_mult_207_n1718), .ZN(DP_mult_207_n1421)
         );
  OAI22_X1 DP_mult_207_U2705 ( .A1(DP_mult_207_n2150), .A2(DP_mult_207_n1716), 
        .B1(DP_mult_207_n1715), .B2(DP_mult_207_n2258), .ZN(DP_mult_207_n1418)
         );
  OAI22_X1 DP_mult_207_U2704 ( .A1(DP_mult_207_n2231), .A2(DP_mult_207_n1712), 
        .B1(DP_mult_207_n1711), .B2(DP_mult_207_n2257), .ZN(DP_mult_207_n1414)
         );
  OAI22_X1 DP_mult_207_U2703 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1722), 
        .B1(DP_mult_207_n1721), .B2(DP_mult_207_n2257), .ZN(DP_mult_207_n1424)
         );
  OAI22_X1 DP_mult_207_U2702 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1729), 
        .B1(DP_mult_207_n2257), .B2(DP_mult_207_n1728), .ZN(DP_mult_207_n1431)
         );
  OAI22_X1 DP_mult_207_U2701 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1728), 
        .B1(DP_mult_207_n1727), .B2(DP_mult_207_n2257), .ZN(DP_mult_207_n1430)
         );
  OAI22_X1 DP_mult_207_U2700 ( .A1(DP_mult_207_n2151), .A2(DP_mult_207_n1710), 
        .B1(DP_mult_207_n1709), .B2(DP_mult_207_n2258), .ZN(DP_mult_207_n1412)
         );
  OAI22_X1 DP_mult_207_U2699 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1723), 
        .B1(DP_mult_207_n2258), .B2(DP_mult_207_n1722), .ZN(DP_mult_207_n1425)
         );
  OAI22_X1 DP_mult_207_U2698 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1725), 
        .B1(DP_mult_207_n2258), .B2(DP_mult_207_n1724), .ZN(DP_mult_207_n1427)
         );
  OAI22_X1 DP_mult_207_U2697 ( .A1(DP_mult_207_n2151), .A2(DP_mult_207_n1708), 
        .B1(DP_mult_207_n1707), .B2(DP_mult_207_n2257), .ZN(DP_mult_207_n874)
         );
  OAI22_X1 DP_mult_207_U2696 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1730), 
        .B1(DP_mult_207_n1729), .B2(DP_mult_207_n2258), .ZN(DP_mult_207_n1432)
         );
  OAI22_X1 DP_mult_207_U2695 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1726), 
        .B1(DP_mult_207_n1725), .B2(DP_mult_207_n2257), .ZN(DP_mult_207_n1428)
         );
  OAI22_X1 DP_mult_207_U2694 ( .A1(DP_mult_207_n2151), .A2(DP_mult_207_n1718), 
        .B1(DP_mult_207_n1717), .B2(DP_mult_207_n2257), .ZN(DP_mult_207_n1420)
         );
  OAI22_X1 DP_mult_207_U2693 ( .A1(DP_mult_207_n2150), .A2(DP_mult_207_n2278), 
        .B1(DP_mult_207_n1731), .B2(DP_mult_207_n2258), .ZN(DP_mult_207_n1191)
         );
  OAI22_X1 DP_mult_207_U2692 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1721), 
        .B1(DP_mult_207_n2258), .B2(DP_mult_207_n1720), .ZN(DP_mult_207_n1423)
         );
  OAI22_X1 DP_mult_207_U2691 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1720), 
        .B1(DP_mult_207_n1719), .B2(DP_mult_207_n2258), .ZN(DP_mult_207_n1422)
         );
  OAI22_X1 DP_mult_207_U2690 ( .A1(DP_mult_207_n2203), .A2(DP_mult_207_n1727), 
        .B1(DP_mult_207_n2257), .B2(DP_mult_207_n1726), .ZN(DP_mult_207_n1429)
         );
  OAI21_X1 DP_mult_207_U2689 ( .B1(DP_mult_207_n536), .B2(DP_mult_207_n498), 
        .A(DP_mult_207_n499), .ZN(DP_mult_207_n497) );
  OAI21_X1 DP_mult_207_U2688 ( .B1(DP_mult_207_n536), .B2(DP_mult_207_n487), 
        .A(DP_mult_207_n488), .ZN(DP_mult_207_n486) );
  OAI21_X1 DP_mult_207_U2687 ( .B1(DP_mult_207_n536), .B2(DP_mult_207_n476), 
        .A(DP_mult_207_n477), .ZN(DP_mult_207_n475) );
  OAI21_X1 DP_mult_207_U2686 ( .B1(DP_mult_207_n536), .B2(DP_mult_207_n523), 
        .A(DP_mult_207_n524), .ZN(DP_mult_207_n522) );
  OAI21_X1 DP_mult_207_U2685 ( .B1(DP_mult_207_n536), .B2(DP_mult_207_n463), 
        .A(DP_mult_207_n464), .ZN(DP_mult_207_n462) );
  OAI21_X1 DP_mult_207_U2684 ( .B1(DP_mult_207_n536), .B2(DP_mult_207_n2208), 
        .A(DP_mult_207_n535), .ZN(DP_mult_207_n533) );
  OAI21_X1 DP_mult_207_U2683 ( .B1(DP_mult_207_n536), .B2(DP_mult_207_n516), 
        .A(DP_mult_207_n517), .ZN(DP_mult_207_n515) );
  OAI21_X1 DP_mult_207_U2682 ( .B1(DP_mult_207_n536), .B2(DP_mult_207_n505), 
        .A(DP_mult_207_n2211), .ZN(DP_mult_207_n504) );
  XNOR2_X1 DP_mult_207_U2681 ( .A(DP_mult_207_n533), .B(DP_mult_207_n320), 
        .ZN(DP_pipe0_coeff_pipe01[4]) );
  XNOR2_X1 DP_mult_207_U2680 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2290), .ZN(
        DP_mult_207_n1642) );
  XNOR2_X1 DP_mult_207_U2679 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2290), .ZN(
        DP_mult_207_n1640) );
  XNOR2_X1 DP_mult_207_U2678 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2016), .ZN(
        DP_mult_207_n1638) );
  XNOR2_X1 DP_mult_207_U2677 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2290), .ZN(
        DP_mult_207_n1644) );
  OAI22_X1 DP_mult_207_U2676 ( .A1(DP_mult_207_n1993), .A2(DP_mult_207_n1608), 
        .B1(DP_mult_207_n1607), .B2(DP_mult_207_n2247), .ZN(DP_mult_207_n746)
         );
  XNOR2_X1 DP_mult_207_U2675 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2016), .ZN(
        DP_mult_207_n1634) );
  XNOR2_X1 DP_mult_207_U2674 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2290), .ZN(
        DP_mult_207_n1636) );
  OAI22_X1 DP_mult_207_U2673 ( .A1(DP_mult_207_n2224), .A2(DP_mult_207_n1614), 
        .B1(DP_mult_207_n1613), .B2(DP_mult_207_n2246), .ZN(DP_mult_207_n1320)
         );
  OAI22_X1 DP_mult_207_U2672 ( .A1(DP_mult_207_n2224), .A2(DP_mult_207_n1618), 
        .B1(DP_mult_207_n1617), .B2(DP_mult_207_n2246), .ZN(DP_mult_207_n1324)
         );
  OAI22_X1 DP_mult_207_U2671 ( .A1(DP_mult_207_n1993), .A2(DP_mult_207_n1609), 
        .B1(DP_mult_207_n2247), .B2(DP_mult_207_n1608), .ZN(DP_mult_207_n1315)
         );
  OAI22_X1 DP_mult_207_U2670 ( .A1(DP_mult_207_n2224), .A2(DP_mult_207_n1616), 
        .B1(DP_mult_207_n1615), .B2(DP_mult_207_n2247), .ZN(DP_mult_207_n1322)
         );
  INV_X1 DP_mult_207_U2669 ( .A(DP_mult_207_n746), .ZN(DP_mult_207_n747) );
  OAI22_X1 DP_mult_207_U2668 ( .A1(DP_mult_207_n2198), .A2(DP_mult_207_n1615), 
        .B1(DP_mult_207_n2246), .B2(DP_mult_207_n1614), .ZN(DP_mult_207_n1321)
         );
  OAI22_X1 DP_mult_207_U2667 ( .A1(DP_mult_207_n2224), .A2(DP_mult_207_n1611), 
        .B1(DP_mult_207_n2246), .B2(DP_mult_207_n1610), .ZN(DP_mult_207_n1317)
         );
  OAI22_X1 DP_mult_207_U2666 ( .A1(DP_mult_207_n1993), .A2(DP_mult_207_n2296), 
        .B1(DP_mult_207_n1631), .B2(DP_mult_207_n2246), .ZN(DP_mult_207_n1187)
         );
  OAI22_X1 DP_mult_207_U2665 ( .A1(DP_mult_207_n2224), .A2(DP_mult_207_n1617), 
        .B1(DP_mult_207_n2247), .B2(DP_mult_207_n1616), .ZN(DP_mult_207_n1323)
         );
  OAI22_X1 DP_mult_207_U2664 ( .A1(DP_mult_207_n1993), .A2(DP_mult_207_n1612), 
        .B1(DP_mult_207_n1611), .B2(DP_mult_207_n2246), .ZN(DP_mult_207_n1318)
         );
  OAI22_X1 DP_mult_207_U2663 ( .A1(DP_mult_207_n1993), .A2(DP_mult_207_n1613), 
        .B1(DP_mult_207_n2247), .B2(DP_mult_207_n1612), .ZN(DP_mult_207_n1319)
         );
  OAI22_X1 DP_mult_207_U2662 ( .A1(DP_mult_207_n1993), .A2(DP_mult_207_n1610), 
        .B1(DP_mult_207_n1609), .B2(DP_mult_207_n2247), .ZN(DP_mult_207_n1316)
         );
  NAND2_X1 DP_mult_207_U2661 ( .A1(DP_mult_207_n717), .A2(DP_mult_207_n726), 
        .ZN(DP_mult_207_n418) );
  AOI21_X1 DP_mult_207_U2660 ( .B1(DP_mult_207_n346), .B2(DP_mult_207_n2182), 
        .A(DP_mult_207_n339), .ZN(DP_mult_207_n337) );
  INV_X1 DP_mult_207_U2659 ( .A(DP_mult_207_n346), .ZN(DP_mult_207_n344) );
  OAI21_X1 DP_mult_207_U2658 ( .B1(DP_mult_207_n2165), .B2(DP_mult_207_n452), 
        .A(DP_mult_207_n453), .ZN(DP_mult_207_n451) );
  OAI22_X1 DP_mult_207_U2657 ( .A1(DP_mult_207_n2234), .A2(DP_mult_207_n1733), 
        .B1(DP_mult_207_n1732), .B2(DP_mult_207_n2259), .ZN(DP_mult_207_n916)
         );
  OAI22_X1 DP_mult_207_U2656 ( .A1(DP_mult_207_n2022), .A2(DP_mult_207_n1605), 
        .B1(DP_mult_207_n1604), .B2(DP_mult_207_n2243), .ZN(DP_mult_207_n1312)
         );
  NAND2_X1 DP_mult_207_U2655 ( .A1(DP_mult_207_n454), .A2(DP_mult_207_n2042), 
        .ZN(DP_mult_207_n452) );
  AOI21_X1 DP_mult_207_U2654 ( .B1(DP_mult_207_n454), .B2(DP_mult_207_n490), 
        .A(DP_mult_207_n455), .ZN(DP_mult_207_n453) );
  AOI21_X1 DP_mult_207_U2653 ( .B1(DP_mult_207_n553), .B2(DP_mult_207_n2126), 
        .A(DP_mult_207_n541), .ZN(DP_mult_207_n539) );
  XNOR2_X1 DP_mult_207_U2652 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2285), .ZN(
        DP_mult_207_n1667) );
  XNOR2_X1 DP_mult_207_U2651 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2092), .ZN(
        DP_mult_207_n1659) );
  XNOR2_X1 DP_mult_207_U2650 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2285), .ZN(
        DP_mult_207_n1665) );
  XNOR2_X1 DP_mult_207_U2649 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2285), .ZN(
        DP_mult_207_n1661) );
  XNOR2_X1 DP_mult_207_U2648 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2285), .ZN(
        DP_mult_207_n1669) );
  XNOR2_X1 DP_mult_207_U2647 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2092), .ZN(
        DP_mult_207_n1663) );
  OAI22_X1 DP_mult_207_U2646 ( .A1(DP_mult_207_n2225), .A2(DP_mult_207_n1650), 
        .B1(DP_mult_207_n2250), .B2(DP_mult_207_n1649), .ZN(DP_mult_207_n1355)
         );
  OAI22_X1 DP_mult_207_U2645 ( .A1(DP_mult_207_n2225), .A2(DP_mult_207_n1651), 
        .B1(DP_mult_207_n1650), .B2(DP_mult_207_n2249), .ZN(DP_mult_207_n1356)
         );
  OAI22_X1 DP_mult_207_U2644 ( .A1(DP_mult_207_n2081), .A2(DP_mult_207_n1646), 
        .B1(DP_mult_207_n2250), .B2(DP_mult_207_n1645), .ZN(DP_mult_207_n1351)
         );
  OAI22_X1 DP_mult_207_U2643 ( .A1(DP_mult_207_n2080), .A2(DP_mult_207_n1647), 
        .B1(DP_mult_207_n1646), .B2(DP_mult_207_n2250), .ZN(DP_mult_207_n1352)
         );
  OAI22_X1 DP_mult_207_U2642 ( .A1(DP_mult_207_n2017), .A2(DP_mult_207_n1655), 
        .B1(DP_mult_207_n1654), .B2(DP_mult_207_n2249), .ZN(DP_mult_207_n1360)
         );
  OAI22_X1 DP_mult_207_U2641 ( .A1(DP_mult_207_n2017), .A2(DP_mult_207_n1654), 
        .B1(DP_mult_207_n2249), .B2(DP_mult_207_n1653), .ZN(DP_mult_207_n1359)
         );
  OAI22_X1 DP_mult_207_U2640 ( .A1(DP_mult_207_n2225), .A2(DP_mult_207_n1644), 
        .B1(DP_mult_207_n2250), .B2(DP_mult_207_n1643), .ZN(DP_mult_207_n1349)
         );
  OAI22_X1 DP_mult_207_U2639 ( .A1(DP_mult_207_n2017), .A2(DP_mult_207_n1648), 
        .B1(DP_mult_207_n2250), .B2(DP_mult_207_n1647), .ZN(DP_mult_207_n1353)
         );
  OAI22_X1 DP_mult_207_U2638 ( .A1(DP_mult_207_n2225), .A2(DP_mult_207_n1653), 
        .B1(DP_mult_207_n1652), .B2(DP_mult_207_n2249), .ZN(DP_mult_207_n1358)
         );
  OAI22_X1 DP_mult_207_U2637 ( .A1(DP_mult_207_n2080), .A2(DP_mult_207_n1645), 
        .B1(DP_mult_207_n1644), .B2(DP_mult_207_n2249), .ZN(DP_mult_207_n1350)
         );
  OAI22_X1 DP_mult_207_U2636 ( .A1(DP_mult_207_n2226), .A2(DP_mult_207_n1649), 
        .B1(DP_mult_207_n1648), .B2(DP_mult_207_n2250), .ZN(DP_mult_207_n1354)
         );
  OAI22_X1 DP_mult_207_U2635 ( .A1(DP_mult_207_n2226), .A2(DP_mult_207_n1652), 
        .B1(DP_mult_207_n2249), .B2(DP_mult_207_n1651), .ZN(DP_mult_207_n1357)
         );
  OAI22_X1 DP_mult_207_U2634 ( .A1(DP_mult_207_n2095), .A2(DP_mult_207_n1504), 
        .B1(DP_mult_207_n2237), .B2(DP_mult_207_n1503), .ZN(DP_mult_207_n1215)
         );
  OAI22_X1 DP_mult_207_U2633 ( .A1(DP_mult_207_n2053), .A2(DP_mult_207_n1498), 
        .B1(DP_mult_207_n2237), .B2(DP_mult_207_n1497), .ZN(DP_mult_207_n1209)
         );
  OAI22_X1 DP_mult_207_U2632 ( .A1(DP_mult_207_n2215), .A2(DP_mult_207_n1505), 
        .B1(DP_mult_207_n1504), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n1216)
         );
  OAI22_X1 DP_mult_207_U2631 ( .A1(DP_mult_207_n2053), .A2(DP_mult_207_n1499), 
        .B1(DP_mult_207_n1498), .B2(DP_mult_207_n2237), .ZN(DP_mult_207_n1210)
         );
  OAI22_X1 DP_mult_207_U2630 ( .A1(DP_mult_207_n2215), .A2(DP_mult_207_n1503), 
        .B1(DP_mult_207_n1502), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n1214)
         );
  OAI22_X1 DP_mult_207_U2629 ( .A1(DP_mult_207_n2053), .A2(DP_mult_207_n1494), 
        .B1(DP_mult_207_n2238), .B2(DP_mult_207_n1493), .ZN(DP_mult_207_n1205)
         );
  OAI22_X1 DP_mult_207_U2628 ( .A1(DP_mult_207_n2053), .A2(DP_mult_207_n1500), 
        .B1(DP_mult_207_n2238), .B2(DP_mult_207_n1499), .ZN(DP_mult_207_n1211)
         );
  OAI22_X1 DP_mult_207_U2627 ( .A1(DP_mult_207_n2094), .A2(DP_mult_207_n1501), 
        .B1(DP_mult_207_n1500), .B2(DP_mult_207_n2237), .ZN(DP_mult_207_n1212)
         );
  OAI22_X1 DP_mult_207_U2626 ( .A1(DP_mult_207_n2094), .A2(DP_mult_207_n1502), 
        .B1(DP_mult_207_n2237), .B2(DP_mult_207_n1501), .ZN(DP_mult_207_n1213)
         );
  OAI22_X1 DP_mult_207_U2625 ( .A1(DP_mult_207_n2053), .A2(DP_mult_207_n1495), 
        .B1(DP_mult_207_n1494), .B2(DP_mult_207_n2238), .ZN(DP_mult_207_n1206)
         );
  OAI22_X1 DP_mult_207_U2624 ( .A1(DP_mult_207_n2095), .A2(DP_mult_207_n1496), 
        .B1(DP_mult_207_n2238), .B2(DP_mult_207_n1495), .ZN(DP_mult_207_n1207)
         );
  OAI22_X1 DP_mult_207_U2623 ( .A1(DP_mult_207_n2096), .A2(DP_mult_207_n1497), 
        .B1(DP_mult_207_n1496), .B2(DP_mult_207_n2238), .ZN(DP_mult_207_n1208)
         );
  XNOR2_X1 DP_mult_207_U2622 ( .A(DP_mult_207_n430), .B(DP_mult_207_n310), 
        .ZN(DP_pipe0_coeff_pipe01[14]) );
  XNOR2_X1 DP_mult_207_U2621 ( .A(DP_coeffs_ff_int[40]), .B(
        DP_coeffs_ff_int[39]), .ZN(DP_mult_207_n259) );
  XNOR2_X1 DP_mult_207_U2620 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2282), .ZN(
        DP_mult_207_n1692) );
  XNOR2_X1 DP_mult_207_U2619 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2281), .ZN(
        DP_mult_207_n1694) );
  XNOR2_X1 DP_mult_207_U2618 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2281), .ZN(
        DP_mult_207_n1684) );
  XNOR2_X1 DP_mult_207_U2617 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2281), .ZN(
        DP_mult_207_n1690) );
  XNOR2_X1 DP_mult_207_U2616 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2282), .ZN(
        DP_mult_207_n1686) );
  XNOR2_X1 DP_mult_207_U2615 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2281), .ZN(
        DP_mult_207_n1688) );
  OAI22_X1 DP_mult_207_U2614 ( .A1(DP_mult_207_n2045), .A2(DP_mult_207_n1668), 
        .B1(DP_mult_207_n1667), .B2(DP_mult_207_n2252), .ZN(DP_mult_207_n1372)
         );
  OAI22_X1 DP_mult_207_U2613 ( .A1(DP_mult_207_n2227), .A2(DP_mult_207_n1659), 
        .B1(DP_mult_207_n2253), .B2(DP_mult_207_n1658), .ZN(DP_mult_207_n1363)
         );
  OAI22_X1 DP_mult_207_U2612 ( .A1(DP_mult_207_n2227), .A2(DP_mult_207_n1662), 
        .B1(DP_mult_207_n1661), .B2(DP_mult_207_n2252), .ZN(DP_mult_207_n1366)
         );
  OAI22_X1 DP_mult_207_U2611 ( .A1(DP_mult_207_n2045), .A2(DP_mult_207_n1665), 
        .B1(DP_mult_207_n2252), .B2(DP_mult_207_n1664), .ZN(DP_mult_207_n1369)
         );
  OAI22_X1 DP_mult_207_U2610 ( .A1(DP_mult_207_n2228), .A2(DP_mult_207_n1658), 
        .B1(DP_mult_207_n1657), .B2(DP_mult_207_n2253), .ZN(DP_mult_207_n802)
         );
  OAI22_X1 DP_mult_207_U2609 ( .A1(DP_mult_207_n2228), .A2(DP_mult_207_n1667), 
        .B1(DP_mult_207_n2253), .B2(DP_mult_207_n1666), .ZN(DP_mult_207_n1371)
         );
  OAI22_X1 DP_mult_207_U2608 ( .A1(DP_mult_207_n2044), .A2(DP_mult_207_n1664), 
        .B1(DP_mult_207_n1663), .B2(DP_mult_207_n2253), .ZN(DP_mult_207_n1368)
         );
  OAI22_X1 DP_mult_207_U2607 ( .A1(DP_mult_207_n2044), .A2(DP_mult_207_n2288), 
        .B1(DP_mult_207_n1681), .B2(DP_mult_207_n2252), .ZN(DP_mult_207_n1189)
         );
  OAI22_X1 DP_mult_207_U2606 ( .A1(DP_mult_207_n2044), .A2(DP_mult_207_n1663), 
        .B1(DP_mult_207_n2253), .B2(DP_mult_207_n1662), .ZN(DP_mult_207_n1367)
         );
  OAI22_X1 DP_mult_207_U2605 ( .A1(DP_mult_207_n2228), .A2(DP_mult_207_n1660), 
        .B1(DP_mult_207_n1659), .B2(DP_mult_207_n2252), .ZN(DP_mult_207_n1364)
         );
  OAI22_X1 DP_mult_207_U2604 ( .A1(DP_mult_207_n2228), .A2(DP_mult_207_n1661), 
        .B1(DP_mult_207_n2252), .B2(DP_mult_207_n1660), .ZN(DP_mult_207_n1365)
         );
  OAI22_X1 DP_mult_207_U2603 ( .A1(DP_mult_207_n2096), .A2(DP_mult_207_n1492), 
        .B1(DP_mult_207_n2238), .B2(DP_mult_207_n1491), .ZN(DP_mult_207_n1203)
         );
  NAND2_X1 DP_mult_207_U2602 ( .A1(DP_mult_207_n362), .A2(DP_mult_207_n2172), 
        .ZN(DP_mult_207_n360) );
  NAND2_X1 DP_mult_207_U2601 ( .A1(DP_mult_207_n356), .A2(DP_mult_207_n2181), 
        .ZN(DP_mult_207_n347) );
  OAI22_X1 DP_mult_207_U2600 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1739), 
        .B1(DP_mult_207_n1738), .B2(DP_mult_207_n2259), .ZN(DP_mult_207_n1440)
         );
  OAI22_X1 DP_mult_207_U2599 ( .A1(DP_mult_207_n2234), .A2(DP_mult_207_n1737), 
        .B1(DP_mult_207_n1736), .B2(DP_mult_207_n2259), .ZN(DP_mult_207_n1438)
         );
  OAI22_X1 DP_mult_207_U2598 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1743), 
        .B1(DP_mult_207_n1742), .B2(DP_mult_207_n1943), .ZN(DP_mult_207_n1444)
         );
  OAI22_X1 DP_mult_207_U2597 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1742), 
        .B1(DP_mult_207_n2259), .B2(DP_mult_207_n1741), .ZN(DP_mult_207_n1443)
         );
  XNOR2_X1 DP_mult_207_U2596 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1765) );
  XNOR2_X1 DP_mult_207_U2595 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1769) );
  XNOR2_X1 DP_mult_207_U2594 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1761) );
  OAI22_X1 DP_mult_207_U2593 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1755), 
        .B1(DP_mult_207_n1754), .B2(DP_mult_207_n1943), .ZN(DP_mult_207_n1456)
         );
  XNOR2_X1 DP_mult_207_U2592 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1759) );
  XNOR2_X1 DP_mult_207_U2591 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1763) );
  XNOR2_X1 DP_mult_207_U2590 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1767) );
  OAI22_X1 DP_mult_207_U2589 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1741), 
        .B1(DP_mult_207_n1740), .B2(DP_mult_207_n2259), .ZN(DP_mult_207_n1442)
         );
  INV_X1 DP_mult_207_U2588 ( .A(DP_mult_207_n2089), .ZN(DP_mult_207_n917) );
  OAI22_X1 DP_mult_207_U2587 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1753), 
        .B1(DP_mult_207_n1752), .B2(DP_mult_207_n2260), .ZN(DP_mult_207_n1454)
         );
  OAI22_X1 DP_mult_207_U2586 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n2274), 
        .B1(DP_mult_207_n1756), .B2(DP_mult_207_n1943), .ZN(DP_mult_207_n1192)
         );
  NAND2_X1 DP_mult_207_U2585 ( .A1(DP_mult_207_n805), .A2(DP_mult_207_n820), 
        .ZN(DP_mult_207_n496) );
  XNOR2_X1 DP_mult_207_U2584 ( .A(DP_mult_207_n419), .B(DP_mult_207_n309), 
        .ZN(DP_pipe0_coeff_pipe01[15]) );
  OAI21_X1 DP_mult_207_U2583 ( .B1(DP_mult_207_n566), .B2(DP_mult_207_n538), 
        .A(DP_mult_207_n539), .ZN(DP_mult_207_n537) );
  OAI22_X1 DP_mult_207_U2582 ( .A1(DP_mult_207_n2222), .A2(DP_mult_207_n1604), 
        .B1(DP_mult_207_n1991), .B2(DP_mult_207_n1603), .ZN(DP_mult_207_n1311)
         );
  OAI22_X1 DP_mult_207_U2581 ( .A1(DP_mult_207_n2003), .A2(DP_mult_207_n1599), 
        .B1(DP_mult_207_n1598), .B2(DP_mult_207_n2242), .ZN(DP_mult_207_n1306)
         );
  OAI22_X1 DP_mult_207_U2580 ( .A1(DP_mult_207_n2222), .A2(DP_mult_207_n2302), 
        .B1(DP_mult_207_n1606), .B2(DP_mult_207_n1991), .ZN(DP_mult_207_n1186)
         );
  OAI22_X1 DP_mult_207_U2579 ( .A1(DP_mult_207_n2003), .A2(DP_mult_207_n1603), 
        .B1(DP_mult_207_n1602), .B2(DP_mult_207_n1991), .ZN(DP_mult_207_n1310)
         );
  OAI22_X1 DP_mult_207_U2578 ( .A1(DP_mult_207_n2221), .A2(DP_mult_207_n1598), 
        .B1(DP_mult_207_n2242), .B2(DP_mult_207_n1597), .ZN(DP_mult_207_n1305)
         );
  OAI22_X1 DP_mult_207_U2577 ( .A1(DP_mult_207_n2221), .A2(DP_mult_207_n1597), 
        .B1(DP_mult_207_n1596), .B2(DP_mult_207_n2243), .ZN(DP_mult_207_n1304)
         );
  OAI22_X1 DP_mult_207_U2576 ( .A1(DP_mult_207_n2023), .A2(DP_mult_207_n1595), 
        .B1(DP_mult_207_n1594), .B2(DP_mult_207_n2243), .ZN(DP_mult_207_n1302)
         );
  OAI22_X1 DP_mult_207_U2575 ( .A1(DP_mult_207_n2222), .A2(DP_mult_207_n1585), 
        .B1(DP_mult_207_n1584), .B2(DP_mult_207_n2242), .ZN(DP_mult_207_n1292)
         );
  OAI22_X1 DP_mult_207_U2574 ( .A1(DP_mult_207_n2023), .A2(DP_mult_207_n1591), 
        .B1(DP_mult_207_n1590), .B2(DP_mult_207_n2242), .ZN(DP_mult_207_n1298)
         );
  OAI22_X1 DP_mult_207_U2573 ( .A1(DP_mult_207_n2222), .A2(DP_mult_207_n1594), 
        .B1(DP_mult_207_n2243), .B2(DP_mult_207_n1593), .ZN(DP_mult_207_n1301)
         );
  OAI22_X1 DP_mult_207_U2572 ( .A1(DP_mult_207_n2022), .A2(DP_mult_207_n1596), 
        .B1(DP_mult_207_n2243), .B2(DP_mult_207_n1595), .ZN(DP_mult_207_n1303)
         );
  OAI22_X1 DP_mult_207_U2571 ( .A1(DP_mult_207_n2222), .A2(DP_mult_207_n1601), 
        .B1(DP_mult_207_n1600), .B2(DP_mult_207_n2242), .ZN(DP_mult_207_n1308)
         );
  OAI22_X1 DP_mult_207_U2570 ( .A1(DP_mult_207_n2023), .A2(DP_mult_207_n1587), 
        .B1(DP_mult_207_n1586), .B2(DP_mult_207_n2242), .ZN(DP_mult_207_n1294)
         );
  OAI22_X1 DP_mult_207_U2569 ( .A1(DP_mult_207_n2003), .A2(DP_mult_207_n1600), 
        .B1(DP_mult_207_n2243), .B2(DP_mult_207_n1599), .ZN(DP_mult_207_n1307)
         );
  OAI22_X1 DP_mult_207_U2568 ( .A1(DP_mult_207_n2023), .A2(DP_mult_207_n1583), 
        .B1(DP_mult_207_n1582), .B2(DP_mult_207_n1991), .ZN(DP_mult_207_n724)
         );
  OAI22_X1 DP_mult_207_U2567 ( .A1(DP_mult_207_n2022), .A2(DP_mult_207_n1602), 
        .B1(DP_mult_207_n2242), .B2(DP_mult_207_n1601), .ZN(DP_mult_207_n1309)
         );
  OAI22_X1 DP_mult_207_U2566 ( .A1(DP_mult_207_n2221), .A2(DP_mult_207_n1589), 
        .B1(DP_mult_207_n1588), .B2(DP_mult_207_n2242), .ZN(DP_mult_207_n1296)
         );
  OAI22_X1 DP_mult_207_U2565 ( .A1(DP_mult_207_n2022), .A2(DP_mult_207_n1593), 
        .B1(DP_mult_207_n1592), .B2(DP_mult_207_n2242), .ZN(DP_mult_207_n1300)
         );
  OAI22_X1 DP_mult_207_U2564 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1527), 
        .B1(DP_mult_207_n2240), .B2(DP_mult_207_n1526), .ZN(DP_mult_207_n1237)
         );
  OAI22_X1 DP_mult_207_U2563 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1530), 
        .B1(DP_mult_207_n1529), .B2(DP_mult_207_n2240), .ZN(DP_mult_207_n1240)
         );
  OAI22_X1 DP_mult_207_U2562 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1528), 
        .B1(DP_mult_207_n1527), .B2(DP_mult_207_n2240), .ZN(DP_mult_207_n1238)
         );
  OAI22_X1 DP_mult_207_U2561 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1529), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1528), .ZN(DP_mult_207_n1239)
         );
  OAI22_X1 DP_mult_207_U2560 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1516), 
        .B1(DP_mult_207_n1515), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n1226)
         );
  OAI22_X1 DP_mult_207_U2559 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1524), 
        .B1(DP_mult_207_n1523), .B2(DP_mult_207_n2240), .ZN(DP_mult_207_n1234)
         );
  OAI22_X1 DP_mult_207_U2558 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n2316), 
        .B1(DP_mult_207_n1531), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n1183)
         );
  OAI22_X1 DP_mult_207_U2557 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1526), 
        .B1(DP_mult_207_n1525), .B2(DP_mult_207_n2240), .ZN(DP_mult_207_n1236)
         );
  OAI22_X1 DP_mult_207_U2556 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1523), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1522), .ZN(DP_mult_207_n1233)
         );
  OAI22_X1 DP_mult_207_U2555 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1525), 
        .B1(DP_mult_207_n2240), .B2(DP_mult_207_n1524), .ZN(DP_mult_207_n1235)
         );
  OAI22_X1 DP_mult_207_U2554 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1512), 
        .B1(DP_mult_207_n1511), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n1222)
         );
  OAI22_X1 DP_mult_207_U2553 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1514), 
        .B1(DP_mult_207_n1513), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n1224)
         );
  OAI22_X1 DP_mult_207_U2552 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1519), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1518), .ZN(DP_mult_207_n1229)
         );
  OAI22_X1 DP_mult_207_U2551 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1510), 
        .B1(DP_mult_207_n1509), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n1220)
         );
  OAI22_X1 DP_mult_207_U2550 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1520), 
        .B1(DP_mult_207_n1519), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n1230)
         );
  OAI22_X1 DP_mult_207_U2549 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1521), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1520), .ZN(DP_mult_207_n1231)
         );
  OAI22_X1 DP_mult_207_U2548 ( .A1(DP_mult_207_n2046), .A2(DP_mult_207_n1522), 
        .B1(DP_mult_207_n1521), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n1232)
         );
  OAI22_X1 DP_mult_207_U2547 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1518), 
        .B1(DP_mult_207_n1517), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n1228)
         );
  OAI22_X1 DP_mult_207_U2546 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1508), 
        .B1(DP_mult_207_n1507), .B2(DP_mult_207_n2239), .ZN(DP_mult_207_n682)
         );
  OAI22_X1 DP_mult_207_U2545 ( .A1(DP_mult_207_n2201), .A2(DP_mult_207_n1551), 
        .B1(DP_mult_207_n1550), .B2(DP_mult_207_n2077), .ZN(DP_mult_207_n1260)
         );
  OAI22_X1 DP_mult_207_U2544 ( .A1(DP_mult_207_n2202), .A2(DP_mult_207_n1553), 
        .B1(DP_mult_207_n1552), .B2(DP_mult_207_n2140), .ZN(DP_mult_207_n1262)
         );
  OAI22_X1 DP_mult_207_U2543 ( .A1(DP_mult_207_n2201), .A2(DP_mult_207_n1554), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1553), .ZN(DP_mult_207_n1263)
         );
  OAI22_X1 DP_mult_207_U2542 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1539), 
        .B1(DP_mult_207_n1538), .B2(DP_mult_207_n2077), .ZN(DP_mult_207_n1248)
         );
  OAI22_X1 DP_mult_207_U2541 ( .A1(DP_mult_207_n2202), .A2(DP_mult_207_n1545), 
        .B1(DP_mult_207_n1544), .B2(DP_mult_207_n2140), .ZN(DP_mult_207_n1254)
         );
  OAI22_X1 DP_mult_207_U2540 ( .A1(DP_mult_207_n2202), .A2(DP_mult_207_n1550), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1549), .ZN(DP_mult_207_n1259)
         );
  OAI22_X1 DP_mult_207_U2539 ( .A1(DP_mult_207_n2201), .A2(DP_mult_207_n1555), 
        .B1(DP_mult_207_n1554), .B2(DP_mult_207_n2077), .ZN(DP_mult_207_n1264)
         );
  OAI22_X1 DP_mult_207_U2538 ( .A1(DP_mult_207_n2202), .A2(DP_mult_207_n1547), 
        .B1(DP_mult_207_n1546), .B2(DP_mult_207_n2140), .ZN(DP_mult_207_n1256)
         );
  OAI22_X1 DP_mult_207_U2537 ( .A1(DP_mult_207_n2202), .A2(DP_mult_207_n1548), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1547), .ZN(DP_mult_207_n1257)
         );
  OAI22_X1 DP_mult_207_U2536 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1533), 
        .B1(DP_mult_207_n1532), .B2(DP_mult_207_n2140), .ZN(DP_mult_207_n692)
         );
  OAI22_X1 DP_mult_207_U2535 ( .A1(DP_mult_207_n2202), .A2(DP_mult_207_n1549), 
        .B1(DP_mult_207_n1548), .B2(DP_mult_207_n2140), .ZN(DP_mult_207_n1258)
         );
  OAI22_X1 DP_mult_207_U2534 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1541), 
        .B1(DP_mult_207_n1540), .B2(DP_mult_207_n2077), .ZN(DP_mult_207_n1250)
         );
  OAI22_X1 DP_mult_207_U2533 ( .A1(DP_mult_207_n2201), .A2(DP_mult_207_n1546), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1545), .ZN(DP_mult_207_n1255)
         );
  OAI22_X1 DP_mult_207_U2532 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n2310), 
        .B1(DP_mult_207_n1556), .B2(DP_mult_207_n2140), .ZN(DP_mult_207_n1184)
         );
  OAI22_X1 DP_mult_207_U2531 ( .A1(DP_mult_207_n2201), .A2(DP_mult_207_n1552), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1551), .ZN(DP_mult_207_n1261)
         );
  OAI22_X1 DP_mult_207_U2530 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1543), 
        .B1(DP_mult_207_n1542), .B2(DP_mult_207_n2077), .ZN(DP_mult_207_n1252)
         );
  OAI22_X1 DP_mult_207_U2529 ( .A1(DP_mult_207_n2201), .A2(DP_mult_207_n1544), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1543), .ZN(DP_mult_207_n1253)
         );
  OAI22_X1 DP_mult_207_U2528 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1537), 
        .B1(DP_mult_207_n1536), .B2(DP_mult_207_n2140), .ZN(DP_mult_207_n1246)
         );
  OAI22_X1 DP_mult_207_U2527 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1535), 
        .B1(DP_mult_207_n1534), .B2(DP_mult_207_n2077), .ZN(DP_mult_207_n1244)
         );
  OAI22_X1 DP_mult_207_U2526 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1703), 
        .B1(DP_mult_207_n1702), .B2(DP_mult_207_n2021), .ZN(DP_mult_207_n1406)
         );
  OAI22_X1 DP_mult_207_U2525 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1705), 
        .B1(DP_mult_207_n1704), .B2(DP_mult_207_n2078), .ZN(DP_mult_207_n1408)
         );
  NAND2_X1 DP_mult_207_U2524 ( .A1(DP_mult_207_n761), .A2(DP_mult_207_n774), 
        .ZN(DP_mult_207_n461) );
  XNOR2_X1 DP_mult_207_U2523 ( .A(DP_mult_207_n410), .B(DP_mult_207_n308), 
        .ZN(DP_pipe0_coeff_pipe01[16]) );
  XNOR2_X1 DP_mult_207_U2522 ( .A(DP_mult_207_n1237), .B(DP_mult_207_n2093), 
        .ZN(DP_mult_207_n939) );
  OR2_X1 DP_mult_207_U2521 ( .A1(DP_mult_207_n1215), .A2(DP_mult_207_n1237), 
        .ZN(DP_mult_207_n938) );
  OAI22_X1 DP_mult_207_U2520 ( .A1(DP_mult_207_n2198), .A2(DP_mult_207_n1628), 
        .B1(DP_mult_207_n1627), .B2(DP_mult_207_n2247), .ZN(DP_mult_207_n1334)
         );
  XNOR2_X1 DP_mult_207_U2519 ( .A(DP_mult_207_n397), .B(DP_mult_207_n307), 
        .ZN(DP_pipe0_coeff_pipe01[17]) );
  OAI21_X1 DP_mult_207_U2518 ( .B1(DP_mult_207_n421), .B2(DP_mult_207_n347), 
        .A(DP_mult_207_n348), .ZN(DP_mult_207_n346) );
  INV_X1 DP_mult_207_U2517 ( .A(DP_mult_207_n421), .ZN(DP_mult_207_n423) );
  OAI21_X1 DP_mult_207_U2516 ( .B1(DP_mult_207_n390), .B2(DP_mult_207_n384), 
        .A(DP_mult_207_n387), .ZN(DP_mult_207_n383) );
  XNOR2_X1 DP_mult_207_U2515 ( .A(DP_mult_207_n370), .B(DP_mult_207_n304), 
        .ZN(DP_pipe0_coeff_pipe01[20]) );
  OAI21_X1 DP_mult_207_U2514 ( .B1(DP_mult_207_n555), .B2(DP_mult_207_n1940), 
        .A(DP_mult_207_n550), .ZN(DP_mult_207_n546) );
  NOR2_X1 DP_mult_207_U2513 ( .A1(DP_mult_207_n1942), .A2(DP_mult_207_n1940), 
        .ZN(DP_mult_207_n545) );
  NOR2_X1 DP_mult_207_U2512 ( .A1(DP_mult_207_n542), .A2(DP_mult_207_n547), 
        .ZN(DP_mult_207_n540) );
  NAND2_X1 DP_mult_207_U2511 ( .A1(DP_mult_207_n839), .A2(DP_mult_207_n856), 
        .ZN(DP_mult_207_n514) );
  OAI22_X1 DP_mult_207_U2510 ( .A1(DP_mult_207_n2096), .A2(DP_mult_207_n1931), 
        .B1(DP_mult_207_n1506), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n1182)
         );
  OAI22_X1 DP_mult_207_U2509 ( .A1(DP_mult_207_n2080), .A2(DP_mult_207_n2291), 
        .B1(DP_mult_207_n1656), .B2(DP_mult_207_n2249), .ZN(DP_mult_207_n1188)
         );
  OAI22_X1 DP_mult_207_U2508 ( .A1(DP_mult_207_n2081), .A2(DP_mult_207_n1641), 
        .B1(DP_mult_207_n1640), .B2(DP_mult_207_n2250), .ZN(DP_mult_207_n1346)
         );
  OAI22_X1 DP_mult_207_U2507 ( .A1(DP_mult_207_n2081), .A2(DP_mult_207_n1643), 
        .B1(DP_mult_207_n1642), .B2(DP_mult_207_n2249), .ZN(DP_mult_207_n1348)
         );
  OAI22_X1 DP_mult_207_U2506 ( .A1(DP_mult_207_n2080), .A2(DP_mult_207_n1642), 
        .B1(DP_mult_207_n2249), .B2(DP_mult_207_n1641), .ZN(DP_mult_207_n1347)
         );
  OAI22_X1 DP_mult_207_U2505 ( .A1(DP_mult_207_n2017), .A2(DP_mult_207_n1633), 
        .B1(DP_mult_207_n1632), .B2(DP_mult_207_n2249), .ZN(DP_mult_207_n772)
         );
  OAI22_X1 DP_mult_207_U2504 ( .A1(DP_mult_207_n2225), .A2(DP_mult_207_n1638), 
        .B1(DP_mult_207_n2249), .B2(DP_mult_207_n1637), .ZN(DP_mult_207_n1343)
         );
  OAI22_X1 DP_mult_207_U2503 ( .A1(DP_mult_207_n2081), .A2(DP_mult_207_n1640), 
        .B1(DP_mult_207_n2249), .B2(DP_mult_207_n1639), .ZN(DP_mult_207_n1345)
         );
  OAI22_X1 DP_mult_207_U2502 ( .A1(DP_mult_207_n2226), .A2(DP_mult_207_n1639), 
        .B1(DP_mult_207_n1638), .B2(DP_mult_207_n2250), .ZN(DP_mult_207_n1344)
         );
  OAI22_X1 DP_mult_207_U2501 ( .A1(DP_mult_207_n2226), .A2(DP_mult_207_n1635), 
        .B1(DP_mult_207_n1634), .B2(DP_mult_207_n2250), .ZN(DP_mult_207_n1340)
         );
  OAI22_X1 DP_mult_207_U2500 ( .A1(DP_mult_207_n2017), .A2(DP_mult_207_n1634), 
        .B1(DP_mult_207_n2250), .B2(DP_mult_207_n1633), .ZN(DP_mult_207_n1339)
         );
  OAI22_X1 DP_mult_207_U2499 ( .A1(DP_mult_207_n2226), .A2(DP_mult_207_n1636), 
        .B1(DP_mult_207_n2250), .B2(DP_mult_207_n1635), .ZN(DP_mult_207_n1341)
         );
  OAI22_X1 DP_mult_207_U2498 ( .A1(DP_mult_207_n2080), .A2(DP_mult_207_n1637), 
        .B1(DP_mult_207_n1636), .B2(DP_mult_207_n2249), .ZN(DP_mult_207_n1342)
         );
  OAI22_X1 DP_mult_207_U2497 ( .A1(DP_mult_207_n2219), .A2(DP_mult_207_n1576), 
        .B1(DP_mult_207_n1575), .B2(DP_mult_207_n2241), .ZN(DP_mult_207_n1284)
         );
  OAI22_X1 DP_mult_207_U2496 ( .A1(DP_mult_207_n2219), .A2(DP_mult_207_n1572), 
        .B1(DP_mult_207_n1571), .B2(DP_mult_207_n2241), .ZN(DP_mult_207_n1280)
         );
  OAI22_X1 DP_mult_207_U2495 ( .A1(DP_mult_207_n2219), .A2(DP_mult_207_n1574), 
        .B1(DP_mult_207_n1573), .B2(DP_mult_207_n2241), .ZN(DP_mult_207_n1282)
         );
  OAI22_X1 DP_mult_207_U2494 ( .A1(DP_mult_207_n2219), .A2(DP_mult_207_n1577), 
        .B1(DP_mult_207_n2241), .B2(DP_mult_207_n1576), .ZN(DP_mult_207_n1285)
         );
  OAI22_X1 DP_mult_207_U2493 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1579), 
        .B1(DP_mult_207_n2241), .B2(DP_mult_207_n1578), .ZN(DP_mult_207_n1287)
         );
  OAI22_X1 DP_mult_207_U2492 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1569), 
        .B1(DP_mult_207_n2008), .B2(DP_mult_207_n1568), .ZN(DP_mult_207_n1277)
         );
  OAI22_X1 DP_mult_207_U2491 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1573), 
        .B1(DP_mult_207_n2241), .B2(DP_mult_207_n1572), .ZN(DP_mult_207_n1281)
         );
  OAI22_X1 DP_mult_207_U2490 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1580), 
        .B1(DP_mult_207_n1579), .B2(DP_mult_207_n2008), .ZN(DP_mult_207_n1288)
         );
  OAI22_X1 DP_mult_207_U2489 ( .A1(DP_mult_207_n2219), .A2(DP_mult_207_n1578), 
        .B1(DP_mult_207_n1577), .B2(DP_mult_207_n2008), .ZN(DP_mult_207_n1286)
         );
  OAI22_X1 DP_mult_207_U2488 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1575), 
        .B1(DP_mult_207_n2241), .B2(DP_mult_207_n1574), .ZN(DP_mult_207_n1283)
         );
  OAI22_X1 DP_mult_207_U2487 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1570), 
        .B1(DP_mult_207_n1569), .B2(DP_mult_207_n2241), .ZN(DP_mult_207_n1278)
         );
  OAI22_X1 DP_mult_207_U2486 ( .A1(DP_mult_207_n2220), .A2(DP_mult_207_n1571), 
        .B1(DP_mult_207_n2008), .B2(DP_mult_207_n1570), .ZN(DP_mult_207_n1279)
         );
  XNOR2_X1 DP_mult_207_U2485 ( .A(DP_mult_207_n388), .B(DP_mult_207_n306), 
        .ZN(DP_pipe0_coeff_pipe01[18]) );
  OAI22_X1 DP_mult_207_U2484 ( .A1(DP_mult_207_n2228), .A2(DP_mult_207_n1670), 
        .B1(DP_mult_207_n1669), .B2(DP_mult_207_n2252), .ZN(DP_mult_207_n1374)
         );
  OAI22_X1 DP_mult_207_U2483 ( .A1(DP_mult_207_n2045), .A2(DP_mult_207_n1676), 
        .B1(DP_mult_207_n1675), .B2(DP_mult_207_n2252), .ZN(DP_mult_207_n1380)
         );
  OAI22_X1 DP_mult_207_U2482 ( .A1(DP_mult_207_n1678), .A2(DP_mult_207_n2044), 
        .B1(DP_mult_207_n1677), .B2(DP_mult_207_n2253), .ZN(DP_mult_207_n1382)
         );
  OAI22_X1 DP_mult_207_U2481 ( .A1(DP_mult_207_n1674), .A2(DP_mult_207_n2227), 
        .B1(DP_mult_207_n1673), .B2(DP_mult_207_n2252), .ZN(DP_mult_207_n1378)
         );
  OAI22_X1 DP_mult_207_U2480 ( .A1(DP_mult_207_n2228), .A2(DP_mult_207_n1680), 
        .B1(DP_mult_207_n1679), .B2(DP_mult_207_n2252), .ZN(DP_mult_207_n1384)
         );
  OAI22_X1 DP_mult_207_U2479 ( .A1(DP_mult_207_n2045), .A2(DP_mult_207_n1679), 
        .B1(DP_mult_207_n2253), .B2(DP_mult_207_n1678), .ZN(DP_mult_207_n1383)
         );
  OAI22_X1 DP_mult_207_U2478 ( .A1(DP_mult_207_n2228), .A2(DP_mult_207_n1671), 
        .B1(DP_mult_207_n2252), .B2(DP_mult_207_n1670), .ZN(DP_mult_207_n1375)
         );
  OAI22_X1 DP_mult_207_U2477 ( .A1(DP_mult_207_n2044), .A2(DP_mult_207_n1675), 
        .B1(DP_mult_207_n2253), .B2(DP_mult_207_n1674), .ZN(DP_mult_207_n1379)
         );
  OAI22_X1 DP_mult_207_U2476 ( .A1(DP_mult_207_n2044), .A2(DP_mult_207_n1669), 
        .B1(DP_mult_207_n2253), .B2(DP_mult_207_n1668), .ZN(DP_mult_207_n1373)
         );
  OAI22_X1 DP_mult_207_U2475 ( .A1(DP_mult_207_n2045), .A2(DP_mult_207_n1673), 
        .B1(DP_mult_207_n2252), .B2(DP_mult_207_n1672), .ZN(DP_mult_207_n1377)
         );
  OAI22_X1 DP_mult_207_U2474 ( .A1(DP_mult_207_n2045), .A2(DP_mult_207_n1677), 
        .B1(DP_mult_207_n2253), .B2(DP_mult_207_n1676), .ZN(DP_mult_207_n1381)
         );
  OAI22_X1 DP_mult_207_U2473 ( .A1(DP_mult_207_n2045), .A2(DP_mult_207_n1672), 
        .B1(DP_mult_207_n1671), .B2(DP_mult_207_n2253), .ZN(DP_mult_207_n1376)
         );
  NOR2_X1 DP_mult_207_U2472 ( .A1(DP_mult_207_n531), .A2(DP_mult_207_n534), 
        .ZN(DP_mult_207_n525) );
  NAND2_X1 DP_mult_207_U2471 ( .A1(DP_mult_207_n525), .A2(DP_mult_207_n511), 
        .ZN(DP_mult_207_n505) );
  INV_X1 DP_mult_207_U2470 ( .A(DP_mult_207_n534), .ZN(DP_mult_207_n672) );
  NAND2_X1 DP_mult_207_U2469 ( .A1(DP_mult_207_n2088), .A2(DP_mult_207_n670), 
        .ZN(DP_mult_207_n516) );
  INV_X1 DP_mult_207_U2468 ( .A(DP_mult_207_n2088), .ZN(DP_mult_207_n523) );
  XNOR2_X1 DP_mult_207_U2467 ( .A(DP_mult_207_n379), .B(DP_mult_207_n305), 
        .ZN(DP_pipe0_coeff_pipe01[19]) );
  AOI21_X1 DP_mult_207_U2466 ( .B1(DP_mult_207_n2160), .B2(DP_mult_207_n670), 
        .A(DP_mult_207_n519), .ZN(DP_mult_207_n517) );
  INV_X1 DP_mult_207_U2465 ( .A(DP_mult_207_n2160), .ZN(DP_mult_207_n524) );
  INV_X1 DP_mult_207_U2464 ( .A(DP_mult_207_n474), .ZN(DP_mult_207_n472) );
  NAND2_X1 DP_mult_207_U2463 ( .A1(DP_mult_207_n1992), .A2(DP_mult_207_n474), 
        .ZN(DP_mult_207_n314) );
  XNOR2_X1 DP_mult_207_U2462 ( .A(DP_mult_207_n353), .B(DP_mult_207_n303), 
        .ZN(DP_pipe0_coeff_pipe01[21]) );
  OAI21_X1 DP_mult_207_U2461 ( .B1(DP_mult_207_n2209), .B2(DP_mult_207_n2210), 
        .A(DP_mult_207_n2331), .ZN(DP_mult_207_n1194) );
  OAI21_X1 DP_mult_207_U2460 ( .B1(DP_mult_207_n2162), .B2(DP_mult_207_n521), 
        .A(DP_mult_207_n514), .ZN(DP_mult_207_n512) );
  INV_X1 DP_mult_207_U2459 ( .A(DP_mult_207_n521), .ZN(DP_mult_207_n519) );
  NAND2_X1 DP_mult_207_U2458 ( .A1(DP_mult_207_n670), .A2(DP_mult_207_n1953), 
        .ZN(DP_mult_207_n319) );
  XNOR2_X1 DP_mult_207_U2457 ( .A(DP_mult_207_n342), .B(DP_mult_207_n302), 
        .ZN(DP_pipe0_coeff_pipe01[22]) );
  AOI21_X1 DP_mult_207_U2456 ( .B1(DP_mult_207_n508), .B2(DP_mult_207_n2115), 
        .A(DP_mult_207_n2163), .ZN(DP_mult_207_n488) );
  NAND2_X1 DP_mult_207_U2455 ( .A1(DP_mult_207_n2207), .A2(DP_mult_207_n2115), 
        .ZN(DP_mult_207_n487) );
  XNOR2_X1 DP_mult_207_U2454 ( .A(DP_mult_207_n475), .B(DP_mult_207_n314), 
        .ZN(DP_pipe0_coeff_pipe01[10]) );
  OAI22_X1 DP_mult_207_U2453 ( .A1(DP_mult_207_n2095), .A2(DP_mult_207_n1493), 
        .B1(DP_mult_207_n1492), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n1204)
         );
  NAND2_X1 DP_mult_207_U2452 ( .A1(DP_mult_207_n1071), .A2(DP_mult_207_n1084), 
        .ZN(DP_mult_207_n591) );
  NAND2_X1 DP_mult_207_U2451 ( .A1(DP_mult_207_n345), .A2(DP_mult_207_n2182), 
        .ZN(DP_mult_207_n336) );
  AOI21_X1 DP_mult_207_U2450 ( .B1(DP_mult_207_n423), .B2(DP_mult_207_n356), 
        .A(DP_mult_207_n359), .ZN(DP_mult_207_n355) );
  NAND2_X1 DP_mult_207_U2449 ( .A1(DP_mult_207_n422), .A2(DP_mult_207_n356), 
        .ZN(DP_mult_207_n354) );
  INV_X1 DP_mult_207_U2448 ( .A(DP_mult_207_n345), .ZN(DP_mult_207_n343) );
  NAND2_X1 DP_mult_207_U2447 ( .A1(DP_mult_207_n2177), .A2(DP_mult_207_n409), 
        .ZN(DP_mult_207_n308) );
  INV_X1 DP_mult_207_U2446 ( .A(DP_mult_207_n2149), .ZN(DP_mult_207_n670) );
  NOR2_X1 DP_mult_207_U2445 ( .A1(DP_mult_207_n520), .A2(DP_mult_207_n513), 
        .ZN(DP_mult_207_n511) );
  NOR2_X1 DP_mult_207_U2444 ( .A1(DP_mult_207_n857), .A2(DP_mult_207_n876), 
        .ZN(DP_mult_207_n520) );
  NAND2_X1 DP_mult_207_U2443 ( .A1(DP_mult_207_n749), .A2(DP_mult_207_n760), 
        .ZN(DP_mult_207_n439) );
  NOR2_X1 DP_mult_207_U2442 ( .A1(DP_mult_207_n749), .A2(DP_mult_207_n760), 
        .ZN(DP_mult_207_n438) );
  NAND2_X1 DP_mult_207_U2441 ( .A1(DP_mult_207_n1992), .A2(DP_mult_207_n666), 
        .ZN(DP_mult_207_n467) );
  AOI21_X1 DP_mult_207_U2440 ( .B1(DP_mult_207_n1992), .B2(DP_mult_207_n483), 
        .A(DP_mult_207_n472), .ZN(DP_mult_207_n468) );
  NAND2_X1 DP_mult_207_U2439 ( .A1(DP_mult_207_n2167), .A2(DP_mult_207_n2168), 
        .ZN(DP_mult_207_n456) );
  OAI22_X1 DP_mult_207_U2438 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1746), 
        .B1(DP_mult_207_n1943), .B2(DP_mult_207_n1745), .ZN(DP_mult_207_n1447)
         );
  OAI22_X1 DP_mult_207_U2437 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1752), 
        .B1(DP_mult_207_n2259), .B2(DP_mult_207_n1751), .ZN(DP_mult_207_n1453)
         );
  OAI22_X1 DP_mult_207_U2436 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1751), 
        .B1(DP_mult_207_n1750), .B2(DP_mult_207_n2260), .ZN(DP_mult_207_n1452)
         );
  OAI21_X1 DP_mult_207_U2435 ( .B1(DP_mult_207_n2085), .B2(DP_mult_207_n503), 
        .A(DP_mult_207_n496), .ZN(DP_mult_207_n490) );
  XNOR2_X1 DP_mult_207_U2434 ( .A(DP_mult_207_n462), .B(DP_mult_207_n313), 
        .ZN(DP_pipe0_coeff_pipe01[11]) );
  NAND2_X1 DP_mult_207_U2433 ( .A1(DP_mult_207_n540), .A2(DP_mult_207_n552), 
        .ZN(DP_mult_207_n538) );
  NOR2_X1 DP_mult_207_U2432 ( .A1(DP_mult_207_n633), .A2(DP_mult_207_n631), 
        .ZN(DP_mult_207_n629) );
  OAI21_X1 DP_mult_207_U2431 ( .B1(DP_mult_207_n638), .B2(DP_mult_207_n636), 
        .A(DP_mult_207_n637), .ZN(DP_mult_207_n635) );
  NAND2_X1 DP_mult_207_U2430 ( .A1(DP_mult_207_n737), .A2(DP_mult_207_n748), 
        .ZN(DP_mult_207_n436) );
  NOR2_X1 DP_mult_207_U2429 ( .A1(DP_mult_207_n737), .A2(DP_mult_207_n748), 
        .ZN(DP_mult_207_n435) );
  INV_X1 DP_mult_207_U2428 ( .A(DP_mult_207_n772), .ZN(DP_mult_207_n773) );
  OAI21_X1 DP_mult_207_U2427 ( .B1(DP_mult_207_n2155), .B2(DP_mult_207_n550), 
        .A(DP_mult_207_n543), .ZN(DP_mult_207_n541) );
  INV_X1 DP_mult_207_U2426 ( .A(DP_mult_207_n382), .ZN(DP_mult_207_n380) );
  NOR2_X1 DP_mult_207_U2425 ( .A1(DP_mult_207_n505), .A2(DP_mult_207_n452), 
        .ZN(DP_mult_207_n450) );
  INV_X1 DP_mult_207_U2424 ( .A(DP_mult_207_n451), .ZN(DP_mult_207_n2214) );
  NAND2_X1 DP_mult_207_U2423 ( .A1(DP_mult_207_n450), .A2(DP_mult_207_n537), 
        .ZN(DP_mult_207_n2213) );
  INV_X1 DP_mult_207_U2422 ( .A(DP_mult_207_n2165), .ZN(DP_mult_207_n508) );
  XNOR2_X1 DP_mult_207_U2421 ( .A(DP_mult_207_n497), .B(DP_mult_207_n316), 
        .ZN(DP_pipe0_coeff_pipe01[8]) );
  AOI21_X1 DP_mult_207_U2420 ( .B1(DP_mult_207_n359), .B2(DP_mult_207_n2181), 
        .A(DP_mult_207_n350), .ZN(DP_mult_207_n348) );
  OAI21_X1 DP_mult_207_U2419 ( .B1(DP_mult_207_n428), .B2(DP_mult_207_n436), 
        .A(DP_mult_207_n429), .ZN(DP_mult_207_n427) );
  INV_X1 DP_mult_207_U2418 ( .A(DP_mult_207_n428), .ZN(DP_mult_207_n661) );
  AOI21_X1 DP_mult_207_U2417 ( .B1(DP_mult_207_n508), .B2(DP_mult_207_n465), 
        .A(DP_mult_207_n466), .ZN(DP_mult_207_n464) );
  AOI21_X1 DP_mult_207_U2416 ( .B1(DP_mult_207_n508), .B2(DP_mult_207_n478), 
        .A(DP_mult_207_n479), .ZN(DP_mult_207_n477) );
  AOI21_X1 DP_mult_207_U2415 ( .B1(DP_mult_207_n508), .B2(DP_mult_207_n668), 
        .A(DP_mult_207_n501), .ZN(DP_mult_207_n499) );
  NAND2_X1 DP_mult_207_U2414 ( .A1(DP_mult_207_n701), .A2(DP_mult_207_n708), 
        .ZN(DP_mult_207_n396) );
  OAI21_X1 DP_mult_207_U2413 ( .B1(DP_mult_207_n405), .B2(DP_mult_207_n360), 
        .A(DP_mult_207_n361), .ZN(DP_mult_207_n359) );
  XNOR2_X1 DP_mult_207_U2412 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1617) );
  XNOR2_X1 DP_mult_207_U2411 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1613) );
  XNOR2_X1 DP_mult_207_U2410 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1615) );
  XNOR2_X1 DP_mult_207_U2409 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1619) );
  XNOR2_X1 DP_mult_207_U2408 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1611) );
  XNOR2_X1 DP_mult_207_U2407 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1609) );
  XNOR2_X1 DP_mult_207_U2406 ( .A(DP_mult_207_n522), .B(DP_mult_207_n319), 
        .ZN(DP_pipe0_coeff_pipe01[5]) );
  XNOR2_X1 DP_mult_207_U2405 ( .A(DP_mult_207_n515), .B(DP_mult_207_n318), 
        .ZN(DP_pipe0_coeff_pipe01[6]) );
  OAI21_X1 DP_mult_207_U2404 ( .B1(DP_mult_207_n2188), .B2(DP_mult_207_n2087), 
        .A(DP_mult_207_n2325), .ZN(DP_mult_207_n1338) );
  XNOR2_X1 DP_mult_207_U2403 ( .A(DP_mult_207_n504), .B(DP_mult_207_n317), 
        .ZN(DP_pipe0_coeff_pipe01[7]) );
  OAI22_X1 DP_mult_207_U2402 ( .A1(DP_mult_207_n2199), .A2(DP_mult_207_n1627), 
        .B1(DP_mult_207_n2247), .B2(DP_mult_207_n1626), .ZN(DP_mult_207_n1333)
         );
  OAI22_X1 DP_mult_207_U2401 ( .A1(DP_mult_207_n2200), .A2(DP_mult_207_n1630), 
        .B1(DP_mult_207_n1629), .B2(DP_mult_207_n2247), .ZN(DP_mult_207_n1336)
         );
  OAI22_X1 DP_mult_207_U2400 ( .A1(DP_mult_207_n2200), .A2(DP_mult_207_n1622), 
        .B1(DP_mult_207_n1621), .B2(DP_mult_207_n2246), .ZN(DP_mult_207_n1328)
         );
  OAI22_X1 DP_mult_207_U2399 ( .A1(DP_mult_207_n2200), .A2(DP_mult_207_n1629), 
        .B1(DP_mult_207_n2247), .B2(DP_mult_207_n1628), .ZN(DP_mult_207_n1335)
         );
  OAI22_X1 DP_mult_207_U2398 ( .A1(DP_mult_207_n2200), .A2(DP_mult_207_n1625), 
        .B1(DP_mult_207_n2246), .B2(DP_mult_207_n1624), .ZN(DP_mult_207_n1331)
         );
  OAI22_X1 DP_mult_207_U2397 ( .A1(DP_mult_207_n2199), .A2(DP_mult_207_n1624), 
        .B1(DP_mult_207_n1623), .B2(DP_mult_207_n2247), .ZN(DP_mult_207_n1330)
         );
  OAI22_X1 DP_mult_207_U2396 ( .A1(DP_mult_207_n2200), .A2(DP_mult_207_n1623), 
        .B1(DP_mult_207_n2247), .B2(DP_mult_207_n1622), .ZN(DP_mult_207_n1329)
         );
  OAI22_X1 DP_mult_207_U2395 ( .A1(DP_mult_207_n2199), .A2(DP_mult_207_n1626), 
        .B1(DP_mult_207_n1625), .B2(DP_mult_207_n2246), .ZN(DP_mult_207_n1332)
         );
  OAI22_X1 DP_mult_207_U2394 ( .A1(DP_mult_207_n2199), .A2(DP_mult_207_n1621), 
        .B1(DP_mult_207_n2246), .B2(DP_mult_207_n1620), .ZN(DP_mult_207_n1327)
         );
  OAI22_X1 DP_mult_207_U2393 ( .A1(DP_mult_207_n2199), .A2(DP_mult_207_n1619), 
        .B1(DP_mult_207_n2247), .B2(DP_mult_207_n1618), .ZN(DP_mult_207_n1325)
         );
  OAI22_X1 DP_mult_207_U2392 ( .A1(DP_mult_207_n2199), .A2(DP_mult_207_n1620), 
        .B1(DP_mult_207_n1619), .B2(DP_mult_207_n2246), .ZN(DP_mult_207_n1326)
         );
  XNOR2_X1 DP_mult_207_U2391 ( .A(DP_mult_207_n486), .B(DP_mult_207_n315), 
        .ZN(DP_pipe0_coeff_pipe01[9]) );
  OAI22_X1 DP_mult_207_U2390 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1740), 
        .B1(DP_mult_207_n1943), .B2(DP_mult_207_n1739), .ZN(DP_mult_207_n1441)
         );
  OAI22_X1 DP_mult_207_U2389 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1736), 
        .B1(DP_mult_207_n2260), .B2(DP_mult_207_n1735), .ZN(DP_mult_207_n1437)
         );
  OAI22_X1 DP_mult_207_U2388 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1734), 
        .B1(DP_mult_207_n2260), .B2(DP_mult_207_n1733), .ZN(DP_mult_207_n1435)
         );
  OAI22_X1 DP_mult_207_U2387 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1738), 
        .B1(DP_mult_207_n2259), .B2(DP_mult_207_n1737), .ZN(DP_mult_207_n1439)
         );
  INV_X1 DP_mult_207_U2386 ( .A(DP_mult_207_n480), .ZN(DP_mult_207_n666) );
  NOR2_X1 DP_mult_207_U2385 ( .A1(DP_mult_207_n456), .A2(DP_mult_207_n480), 
        .ZN(DP_mult_207_n454) );
  NOR2_X1 DP_mult_207_U2384 ( .A1(DP_mult_207_n491), .A2(DP_mult_207_n467), 
        .ZN(DP_mult_207_n465) );
  OAI21_X1 DP_mult_207_U2383 ( .B1(DP_mult_207_n492), .B2(DP_mult_207_n480), 
        .A(DP_mult_207_n481), .ZN(DP_mult_207_n479) );
  NOR2_X1 DP_mult_207_U2382 ( .A1(DP_mult_207_n491), .A2(DP_mult_207_n480), 
        .ZN(DP_mult_207_n478) );
  OAI21_X1 DP_mult_207_U2381 ( .B1(DP_mult_207_n492), .B2(DP_mult_207_n467), 
        .A(DP_mult_207_n468), .ZN(DP_mult_207_n466) );
  OAI22_X1 DP_mult_207_U2380 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1744), 
        .B1(DP_mult_207_n2260), .B2(DP_mult_207_n1743), .ZN(DP_mult_207_n1445)
         );
  OAI21_X1 DP_mult_207_U2379 ( .B1(DP_mult_207_n631), .B2(DP_mult_207_n634), 
        .A(DP_mult_207_n632), .ZN(DP_mult_207_n630) );
  AOI21_X1 DP_mult_207_U2378 ( .B1(DP_mult_207_n629), .B2(DP_mult_207_n635), 
        .A(DP_mult_207_n630), .ZN(DP_mult_207_n628) );
  OAI21_X1 DP_mult_207_U2377 ( .B1(DP_mult_207_n594), .B2(DP_mult_207_n582), 
        .A(DP_mult_207_n583), .ZN(DP_mult_207_n581) );
  AOI21_X1 DP_mult_207_U2376 ( .B1(DP_mult_207_n581), .B2(DP_mult_207_n567), 
        .A(DP_mult_207_n568), .ZN(DP_mult_207_n566) );
  NOR2_X1 DP_mult_207_U2375 ( .A1(DP_mult_207_n336), .A2(DP_mult_207_n334), 
        .ZN(DP_mult_207_n332) );
  NAND2_X1 DP_mult_207_U2374 ( .A1(DP_mult_207_n963), .A2(DP_mult_207_n982), 
        .ZN(DP_mult_207_n559) );
  NAND2_X1 DP_mult_207_U2373 ( .A1(DP_mult_207_n1003), .A2(DP_mult_207_n1020), 
        .ZN(DP_mult_207_n570) );
  INV_X1 DP_mult_207_U2372 ( .A(DP_mult_207_n2148), .ZN(DP_mult_207_n565) );
  OAI21_X1 DP_mult_207_U2371 ( .B1(DP_mult_207_n456), .B2(DP_mult_207_n481), 
        .A(DP_mult_207_n457), .ZN(DP_mult_207_n455) );
  INV_X1 DP_mult_207_U2370 ( .A(DP_mult_207_n508), .ZN(DP_mult_207_n2211) );
  OAI21_X1 DP_mult_207_U2369 ( .B1(DP_mult_207_n572), .B2(DP_mult_207_n1950), 
        .A(DP_mult_207_n570), .ZN(DP_mult_207_n568) );
  OAI22_X1 DP_mult_207_U2368 ( .A1(DP_mult_207_n2114), .A2(DP_mult_207_n1697), 
        .B1(DP_mult_207_n1696), .B2(DP_mult_207_n2255), .ZN(DP_mult_207_n1400)
         );
  INV_X1 DP_mult_207_U2367 ( .A(DP_mult_207_n490), .ZN(DP_mult_207_n492) );
  NAND2_X1 DP_mult_207_U2366 ( .A1(DP_mult_207_n918), .A2(DP_mult_207_n897), 
        .ZN(DP_mult_207_n535) );
  NOR2_X1 DP_mult_207_U2365 ( .A1(DP_mult_207_n918), .A2(DP_mult_207_n897), 
        .ZN(DP_mult_207_n534) );
  XNOR2_X1 DP_mult_207_U2364 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2304), .ZN(
        DP_mult_207_n1567) );
  XNOR2_X1 DP_mult_207_U2363 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2304), .ZN(
        DP_mult_207_n1561) );
  XNOR2_X1 DP_mult_207_U2362 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2304), .ZN(
        DP_mult_207_n1569) );
  XNOR2_X1 DP_mult_207_U2361 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2304), .ZN(
        DP_mult_207_n1563) );
  XNOR2_X1 DP_mult_207_U2360 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2304), .ZN(
        DP_mult_207_n1565) );
  XNOR2_X1 DP_mult_207_U2359 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2304), .ZN(
        DP_mult_207_n1559) );
  OAI22_X1 DP_mult_207_U2358 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n2267), 
        .B1(DP_mult_207_n1781), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1193)
         );
  INV_X1 DP_mult_207_U2357 ( .A(DP_mult_207_n2042), .ZN(DP_mult_207_n491) );
  INV_X1 DP_mult_207_U2356 ( .A(DP_mult_207_n502), .ZN(DP_mult_207_n668) );
  NAND2_X1 DP_mult_207_U2355 ( .A1(DP_mult_207_n1099), .A2(DP_mult_207_n1110), 
        .ZN(DP_mult_207_n598) );
  XNOR2_X1 DP_mult_207_U2354 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2308), .ZN(
        DP_mult_207_n1538) );
  XNOR2_X1 DP_mult_207_U2353 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2309), .ZN(
        DP_mult_207_n1540) );
  XNOR2_X1 DP_mult_207_U2352 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2308), .ZN(
        DP_mult_207_n1544) );
  XNOR2_X1 DP_mult_207_U2351 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2308), .ZN(
        DP_mult_207_n1542) );
  XNOR2_X1 DP_mult_207_U2350 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2309), .ZN(
        DP_mult_207_n1536) );
  XNOR2_X1 DP_mult_207_U2349 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2308), .ZN(
        DP_mult_207_n1534) );
  OAI21_X1 DP_mult_207_U2348 ( .B1(DP_mult_207_n2090), .B2(DP_mult_207_n535), 
        .A(DP_mult_207_n532), .ZN(DP_mult_207_n526) );
  NOR2_X1 DP_mult_207_U2347 ( .A1(DP_mult_207_n1085), .A2(DP_mult_207_n1098), 
        .ZN(DP_mult_207_n592) );
  NAND2_X1 DP_mult_207_U2346 ( .A1(DP_mult_207_n1085), .A2(DP_mult_207_n1098), 
        .ZN(DP_mult_207_n593) );
  INV_X1 DP_mult_207_U2345 ( .A(DP_mult_207_n706), .ZN(DP_mult_207_n707) );
  NAND2_X1 DP_mult_207_U2344 ( .A1(DP_mult_207_n685), .A2(DP_mult_207_n688), 
        .ZN(DP_mult_207_n369) );
  OAI21_X1 DP_mult_207_U2343 ( .B1(DP_mult_207_n337), .B2(DP_mult_207_n334), 
        .A(DP_mult_207_n335), .ZN(DP_mult_207_n333) );
  OAI22_X1 DP_mult_207_U2342 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1754), 
        .B1(DP_mult_207_n2259), .B2(DP_mult_207_n1753), .ZN(DP_mult_207_n1455)
         );
  OAI22_X1 DP_mult_207_U2341 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1749), 
        .B1(DP_mult_207_n1748), .B2(DP_mult_207_n2259), .ZN(DP_mult_207_n1450)
         );
  OAI22_X1 DP_mult_207_U2340 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1750), 
        .B1(DP_mult_207_n2260), .B2(DP_mult_207_n1749), .ZN(DP_mult_207_n1451)
         );
  OAI22_X1 DP_mult_207_U2339 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1745), 
        .B1(DP_mult_207_n1744), .B2(DP_mult_207_n2259), .ZN(DP_mult_207_n1446)
         );
  OAI22_X1 DP_mult_207_U2338 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1748), 
        .B1(DP_mult_207_n1943), .B2(DP_mult_207_n1747), .ZN(DP_mult_207_n1449)
         );
  OAI22_X1 DP_mult_207_U2337 ( .A1(DP_mult_207_n2233), .A2(DP_mult_207_n1747), 
        .B1(DP_mult_207_n1746), .B2(DP_mult_207_n2259), .ZN(DP_mult_207_n1448)
         );
  INV_X1 DP_mult_207_U2336 ( .A(DP_mult_207_n672), .ZN(DP_mult_207_n2208) );
  INV_X1 DP_mult_207_U2335 ( .A(DP_mult_207_n2083), .ZN(DP_mult_207_n2259) );
  OAI21_X1 DP_mult_207_U2334 ( .B1(DP_mult_207_n2195), .B2(DP_mult_207_n2084), 
        .A(DP_mult_207_n2321), .ZN(DP_mult_207_n1434) );
  OAI21_X1 DP_mult_207_U2333 ( .B1(DP_mult_207_n2193), .B2(DP_mult_207_n1945), 
        .A(DP_mult_207_n2324), .ZN(DP_mult_207_n1362) );
  AOI21_X1 DP_mult_207_U2332 ( .B1(DP_mult_207_n333), .B2(DP_mult_207_n2183), 
        .A(DP_mult_207_n2179), .ZN(DP_mult_207_n327) );
  NAND2_X1 DP_mult_207_U2331 ( .A1(DP_mult_207_n877), .A2(DP_mult_207_n896), 
        .ZN(DP_mult_207_n532) );
  NAND3_X1 DP_mult_207_U2330 ( .A1(DP_mult_207_n2204), .A2(DP_mult_207_n2205), 
        .A3(DP_mult_207_n2206), .ZN(DP_mult_207_n896) );
  NAND2_X1 DP_mult_207_U2329 ( .A1(DP_mult_207_n1995), .A2(DP_mult_207_n901), 
        .ZN(DP_mult_207_n2206) );
  NAND2_X1 DP_mult_207_U2328 ( .A1(DP_mult_207_n899), .A2(DP_mult_207_n901), 
        .ZN(DP_mult_207_n2205) );
  NAND2_X1 DP_mult_207_U2327 ( .A1(DP_mult_207_n899), .A2(DP_mult_207_n1995), 
        .ZN(DP_mult_207_n2204) );
  INV_X1 DP_mult_207_U2326 ( .A(DP_mult_207_n2191), .ZN(DP_mult_207_n2230) );
  OAI21_X1 DP_mult_207_U2325 ( .B1(DP_mult_207_n2097), .B2(DP_mult_207_n564), 
        .A(DP_mult_207_n559), .ZN(DP_mult_207_n553) );
  INV_X1 DP_mult_207_U2324 ( .A(DP_mult_207_n553), .ZN(DP_mult_207_n555) );
  AOI21_X1 DP_mult_207_U2323 ( .B1(DP_mult_207_n565), .B2(DP_mult_207_n1985), 
        .A(DP_mult_207_n2075), .ZN(DP_mult_207_n551) );
  NAND2_X1 DP_mult_207_U2322 ( .A1(DP_mult_207_n332), .A2(DP_mult_207_n2183), 
        .ZN(DP_mult_207_n326) );
  INV_X1 DP_mult_207_U2321 ( .A(DP_mult_207_n2195), .ZN(DP_mult_207_n2234) );
  NOR2_X1 DP_mult_207_U2320 ( .A1(DP_mult_207_n571), .A2(DP_mult_207_n569), 
        .ZN(DP_mult_207_n567) );
  INV_X1 DP_mult_207_U2319 ( .A(DP_mult_207_n1988), .ZN(DP_mult_207_n2246) );
  AOI21_X1 DP_mult_207_U2318 ( .B1(DP_mult_207_n2169), .B2(DP_mult_207_n1966), 
        .A(DP_mult_207_n1973), .ZN(DP_mult_207_n572) );
  NAND2_X1 DP_mult_207_U2317 ( .A1(DP_mult_207_n2169), .A2(DP_mult_207_n2170), 
        .ZN(DP_mult_207_n571) );
  NAND2_X1 DP_mult_207_U2316 ( .A1(DP_mult_207_n2176), .A2(DP_mult_207_n2174), 
        .ZN(DP_mult_207_n599) );
  OAI22_X1 DP_mult_207_U2315 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1702), 
        .B1(DP_mult_207_n2078), .B2(DP_mult_207_n1701), .ZN(DP_mult_207_n1405)
         );
  OAI22_X1 DP_mult_207_U2314 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1700), 
        .B1(DP_mult_207_n2021), .B2(DP_mult_207_n1699), .ZN(DP_mult_207_n1403)
         );
  OAI22_X1 DP_mult_207_U2313 ( .A1(DP_mult_207_n2196), .A2(DP_mult_207_n1694), 
        .B1(DP_mult_207_n1958), .B2(DP_mult_207_n1693), .ZN(DP_mult_207_n1397)
         );
  OAI22_X1 DP_mult_207_U2312 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1698), 
        .B1(DP_mult_207_n1958), .B2(DP_mult_207_n1697), .ZN(DP_mult_207_n1401)
         );
  OAI22_X1 DP_mult_207_U2311 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1704), 
        .B1(DP_mult_207_n2078), .B2(DP_mult_207_n1703), .ZN(DP_mult_207_n1407)
         );
  OAI22_X1 DP_mult_207_U2310 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1701), 
        .B1(DP_mult_207_n1700), .B2(DP_mult_207_n2078), .ZN(DP_mult_207_n1404)
         );
  OAI22_X1 DP_mult_207_U2309 ( .A1(DP_mult_207_n2197), .A2(DP_mult_207_n1695), 
        .B1(DP_mult_207_n1694), .B2(DP_mult_207_n2255), .ZN(DP_mult_207_n1398)
         );
  INV_X1 DP_mult_207_U2308 ( .A(DP_mult_207_n2192), .ZN(DP_mult_207_n2223) );
  OAI21_X1 DP_mult_207_U2307 ( .B1(DP_mult_207_n2192), .B2(DP_mult_207_n2005), 
        .A(DP_mult_207_n2326), .ZN(DP_mult_207_n1314) );
  AOI21_X1 DP_mult_207_U2306 ( .B1(DP_mult_207_n2168), .B2(DP_mult_207_n472), 
        .A(DP_mult_207_n459), .ZN(DP_mult_207_n457) );
  NOR2_X1 DP_mult_207_U2305 ( .A1(DP_mult_207_n839), .A2(DP_mult_207_n856), 
        .ZN(DP_mult_207_n513) );
  NAND2_X1 DP_mult_207_U2304 ( .A1(DP_mult_207_n1941), .A2(DP_mult_207_n940), 
        .ZN(DP_mult_207_n543) );
  NAND2_X1 DP_mult_207_U2303 ( .A1(DP_mult_207_n426), .A2(DP_mult_207_n663), 
        .ZN(DP_mult_207_n420) );
  NOR2_X1 DP_mult_207_U2302 ( .A1(DP_mult_207_n420), .A2(DP_mult_207_n347), 
        .ZN(DP_mult_207_n345) );
  INV_X1 DP_mult_207_U2301 ( .A(DP_mult_207_n420), .ZN(DP_mult_207_n422) );
  NOR2_X1 DP_mult_207_U2300 ( .A1(DP_mult_207_n821), .A2(DP_mult_207_n838), 
        .ZN(DP_mult_207_n502) );
  NOR2_X1 DP_mult_207_U2299 ( .A1(DP_mult_207_n805), .A2(DP_mult_207_n820), 
        .ZN(DP_mult_207_n495) );
  INV_X1 DP_mult_207_U2298 ( .A(DP_mult_207_n439), .ZN(DP_mult_207_n445) );
  INV_X1 DP_mult_207_U2297 ( .A(DP_mult_207_n383), .ZN(DP_mult_207_n381) );
  INV_X1 DP_mult_207_U2296 ( .A(DP_mult_207_n2267), .ZN(DP_mult_207_n2263) );
  INV_X1 DP_mult_207_U2295 ( .A(DP_mult_207_n2190), .ZN(DP_mult_207_n2231) );
  INV_X1 DP_mult_207_U2294 ( .A(DP_mult_207_n1984), .ZN(DP_mult_207_n2217) );
  OAI22_X1 DP_mult_207_U2293 ( .A1(DP_mult_207_n2151), .A2(DP_mult_207_n1715), 
        .B1(DP_mult_207_n2258), .B2(DP_mult_207_n1714), .ZN(DP_mult_207_n1417)
         );
  OAI22_X1 DP_mult_207_U2292 ( .A1(DP_mult_207_n2150), .A2(DP_mult_207_n1711), 
        .B1(DP_mult_207_n2257), .B2(DP_mult_207_n1710), .ZN(DP_mult_207_n1413)
         );
  OAI22_X1 DP_mult_207_U2291 ( .A1(DP_mult_207_n2231), .A2(DP_mult_207_n1709), 
        .B1(DP_mult_207_n2258), .B2(DP_mult_207_n1708), .ZN(DP_mult_207_n1411)
         );
  OAI22_X1 DP_mult_207_U2290 ( .A1(DP_mult_207_n2150), .A2(DP_mult_207_n1717), 
        .B1(DP_mult_207_n2257), .B2(DP_mult_207_n1716), .ZN(DP_mult_207_n1419)
         );
  OAI22_X1 DP_mult_207_U2289 ( .A1(DP_mult_207_n2231), .A2(DP_mult_207_n1713), 
        .B1(DP_mult_207_n2258), .B2(DP_mult_207_n1712), .ZN(DP_mult_207_n1415)
         );
  INV_X1 DP_mult_207_U2288 ( .A(DP_mult_207_n2191), .ZN(DP_mult_207_n2229) );
  OAI22_X1 DP_mult_207_U2287 ( .A1(DP_mult_207_n2003), .A2(DP_mult_207_n1586), 
        .B1(DP_mult_207_n1991), .B2(DP_mult_207_n1585), .ZN(DP_mult_207_n1293)
         );
  OAI22_X1 DP_mult_207_U2286 ( .A1(DP_mult_207_n2221), .A2(DP_mult_207_n1592), 
        .B1(DP_mult_207_n2242), .B2(DP_mult_207_n1591), .ZN(DP_mult_207_n1299)
         );
  OAI22_X1 DP_mult_207_U2285 ( .A1(DP_mult_207_n2023), .A2(DP_mult_207_n1588), 
        .B1(DP_mult_207_n1991), .B2(DP_mult_207_n1587), .ZN(DP_mult_207_n1295)
         );
  OAI22_X1 DP_mult_207_U2284 ( .A1(DP_mult_207_n2022), .A2(DP_mult_207_n1590), 
        .B1(DP_mult_207_n2242), .B2(DP_mult_207_n1589), .ZN(DP_mult_207_n1297)
         );
  OAI22_X1 DP_mult_207_U2283 ( .A1(DP_mult_207_n2221), .A2(DP_mult_207_n1584), 
        .B1(DP_mult_207_n1991), .B2(DP_mult_207_n1583), .ZN(DP_mult_207_n1291)
         );
  OAI21_X1 DP_mult_207_U2282 ( .B1(DP_mult_207_n2067), .B2(DP_mult_207_n1944), 
        .A(DP_mult_207_n2330), .ZN(DP_mult_207_n1218) );
  XNOR2_X1 DP_mult_207_U2281 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1482) );
  INV_X1 DP_mult_207_U2280 ( .A(DP_coeffs_ff_int[47]), .ZN(DP_mult_207_n251)
         );
  XNOR2_X1 DP_mult_207_U2279 ( .A(DP_mult_207_n2272), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1755) );
  OAI22_X1 DP_mult_207_U2278 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1778), 
        .B1(DP_mult_207_n1777), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1479)
         );
  XNOR2_X1 DP_mult_207_U2277 ( .A(DP_mult_207_n2300), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1605) );
  AND2_X2 DP_mult_207_U2276 ( .A1(DP_mult_207_n1816), .A2(DP_mult_207_n1954), 
        .ZN(DP_mult_207_n2195) );
  XNOR2_X1 DP_mult_207_U2275 ( .A(DP_mult_207_n2266), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1780) );
  OAI22_X1 DP_mult_207_U2274 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1780), 
        .B1(DP_mult_207_n1779), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1481)
         );
  XNOR2_X1 DP_mult_207_U2273 ( .A(DP_mult_207_n2295), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1630) );
  INV_X1 DP_mult_207_U2272 ( .A(DP_mult_207_n259), .ZN(DP_mult_207_n2254) );
  INV_X1 DP_mult_207_U2271 ( .A(DP_mult_207_n1757), .ZN(DP_mult_207_n2320) );
  OAI21_X1 DP_mult_207_U2270 ( .B1(DP_coeffs_ff_int[47]), .B2(
        DP_mult_207_n1971), .A(DP_mult_207_n2320), .ZN(DP_mult_207_n1458) );
  NAND2_X1 DP_mult_207_U2269 ( .A1(DP_mult_207_n2168), .A2(DP_mult_207_n461), 
        .ZN(DP_mult_207_n313) );
  NAND2_X1 DP_mult_207_U2268 ( .A1(DP_mult_207_n666), .A2(DP_mult_207_n481), 
        .ZN(DP_mult_207_n315) );
  NAND2_X1 DP_mult_207_U2267 ( .A1(DP_mult_207_n2164), .A2(DP_mult_207_n496), 
        .ZN(DP_mult_207_n316) );
  NAND2_X1 DP_mult_207_U2266 ( .A1(DP_mult_207_n668), .A2(DP_mult_207_n503), 
        .ZN(DP_mult_207_n317) );
  NAND2_X1 DP_mult_207_U2265 ( .A1(DP_mult_207_n514), .A2(DP_mult_207_n2091), 
        .ZN(DP_mult_207_n318) );
  NAND2_X1 DP_mult_207_U2264 ( .A1(DP_mult_207_n2161), .A2(DP_mult_207_n1952), 
        .ZN(DP_mult_207_n320) );
  INV_X1 DP_mult_207_U2263 ( .A(DP_mult_207_n265), .ZN(DP_mult_207_n2244) );
  AND2_X2 DP_mult_207_U2262 ( .A1(DP_mult_207_n1810), .A2(DP_mult_207_n265), 
        .ZN(DP_mult_207_n2189) );
  XNOR2_X1 DP_mult_207_U2261 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1492) );
  XNOR2_X1 DP_mult_207_U2260 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2311), .ZN(
        DP_mult_207_n1519) );
  XNOR2_X1 DP_mult_207_U2259 ( .A(DP_pipe01[11]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1494) );
  XNOR2_X1 DP_mult_207_U2258 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2311), .ZN(
        DP_mult_207_n1509) );
  XNOR2_X1 DP_mult_207_U2257 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2311), .ZN(
        DP_mult_207_n1513) );
  XNOR2_X1 DP_mult_207_U2256 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2311), .ZN(
        DP_mult_207_n1511) );
  XNOR2_X1 DP_mult_207_U2255 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2311), .ZN(
        DP_mult_207_n1515) );
  XNOR2_X1 DP_mult_207_U2254 ( .A(DP_pipe01[13]), .B(DP_mult_207_n2311), .ZN(
        DP_mult_207_n1517) );
  XOR2_X1 DP_mult_207_U2253 ( .A(DP_coeffs_ff_int[47]), .B(DP_mult_207_n2263), 
        .Z(DP_mult_207_n1817) );
  XNOR2_X1 DP_mult_207_U2252 ( .A(DP_mult_207_n2318), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1505) );
  XNOR2_X1 DP_mult_207_U2251 ( .A(DP_mult_207_n2290), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1655) );
  XNOR2_X1 DP_mult_207_U2250 ( .A(DP_mult_207_n2277), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1730) );
  OAI22_X1 DP_mult_207_U2249 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1776), 
        .B1(DP_mult_207_n1775), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1477)
         );
  XNOR2_X1 DP_mult_207_U2248 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1729) );
  XNOR2_X1 DP_mult_207_U2247 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1629) );
  XNOR2_X1 DP_mult_207_U2246 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2307), .ZN(
        DP_mult_207_n1548) );
  XNOR2_X1 DP_mult_207_U2245 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1752) );
  XNOR2_X1 DP_mult_207_U2244 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2015), .ZN(
        DP_mult_207_n1652) );
  XNOR2_X1 DP_mult_207_U2243 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1754) );
  XNOR2_X1 DP_mult_207_U2242 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2312), .ZN(
        DP_mult_207_n1525) );
  XNOR2_X1 DP_mult_207_U2241 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2318), .ZN(
        DP_mult_207_n1502) );
  XNOR2_X1 DP_mult_207_U2240 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2057), .ZN(
        DP_mult_207_n1571) );
  XNOR2_X1 DP_mult_207_U2239 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1500) );
  XNOR2_X1 DP_mult_207_U2238 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2312), .ZN(
        DP_mult_207_n1523) );
  XNOR2_X1 DP_mult_207_U2237 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1750) );
  XNOR2_X1 DP_mult_207_U2236 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2280), .ZN(
        DP_mult_207_n1704) );
  XNOR2_X1 DP_mult_207_U2235 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2307), .ZN(
        DP_mult_207_n1546) );
  XNOR2_X1 DP_mult_207_U2234 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2318), .ZN(
        DP_mult_207_n1504) );
  XNOR2_X1 DP_mult_207_U2233 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2312), .ZN(
        DP_mult_207_n1527) );
  XNOR2_X1 DP_mult_207_U2232 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1723) );
  XNOR2_X1 DP_mult_207_U2231 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2092), .ZN(
        DP_mult_207_n1679) );
  XNOR2_X1 DP_mult_207_U2230 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2280), .ZN(
        DP_mult_207_n1702) );
  XNOR2_X1 DP_mult_207_U2229 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2318), .ZN(
        DP_mult_207_n1498) );
  XNOR2_X1 DP_mult_207_U2228 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2312), .ZN(
        DP_mult_207_n1521) );
  XNOR2_X1 DP_mult_207_U2227 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2092), .ZN(
        DP_mult_207_n1677) );
  XNOR2_X1 DP_mult_207_U2226 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2016), .ZN(
        DP_mult_207_n1654) );
  XNOR2_X1 DP_mult_207_U2225 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1727) );
  XNOR2_X1 DP_mult_207_U2224 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2092), .ZN(
        DP_mult_207_n1675) );
  XNOR2_X1 DP_mult_207_U2223 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1725) );
  XNOR2_X1 DP_mult_207_U2222 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1748) );
  XNOR2_X1 DP_mult_207_U2221 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2308), .ZN(
        DP_mult_207_n1550) );
  XNOR2_X1 DP_mult_207_U2220 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1596) );
  XNOR2_X1 DP_mult_207_U2219 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2280), .ZN(
        DP_mult_207_n1700) );
  XNOR2_X1 DP_mult_207_U2218 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1746) );
  XNOR2_X1 DP_mult_207_U2217 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2057), .ZN(
        DP_mult_207_n1573) );
  XNOR2_X1 DP_mult_207_U2216 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1721) );
  XNOR2_X1 DP_mult_207_U2215 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1496) );
  XNOR2_X1 DP_mult_207_U2214 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2312), .ZN(
        DP_mult_207_n1529) );
  XNOR2_X1 DP_mult_207_U2213 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2307), .ZN(
        DP_mult_207_n1552) );
  XNOR2_X1 DP_mult_207_U2212 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2057), .ZN(
        DP_mult_207_n1575) );
  XNOR2_X1 DP_mult_207_U2211 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1621) );
  XNOR2_X1 DP_mult_207_U2210 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1598) );
  XNOR2_X1 DP_mult_207_U2209 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2057), .ZN(
        DP_mult_207_n1577) );
  XNOR2_X1 DP_mult_207_U2208 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2016), .ZN(
        DP_mult_207_n1646) );
  XNOR2_X1 DP_mult_207_U2207 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2307), .ZN(
        DP_mult_207_n1554) );
  XNOR2_X1 DP_mult_207_U2206 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1623) );
  XNOR2_X1 DP_mult_207_U2205 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2285), .ZN(
        DP_mult_207_n1673) );
  XNOR2_X1 DP_mult_207_U2204 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2015), .ZN(
        DP_mult_207_n1650) );
  XNOR2_X1 DP_mult_207_U2203 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1602) );
  XNOR2_X1 DP_mult_207_U2202 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2057), .ZN(
        DP_mult_207_n1579) );
  XNOR2_X1 DP_mult_207_U2201 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1600) );
  XNOR2_X1 DP_mult_207_U2200 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2092), .ZN(
        DP_mult_207_n1671) );
  XNOR2_X1 DP_mult_207_U2199 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1625) );
  XNOR2_X1 DP_mult_207_U2198 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2015), .ZN(
        DP_mult_207_n1648) );
  XNOR2_X1 DP_mult_207_U2197 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1604) );
  XNOR2_X1 DP_mult_207_U2196 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1627) );
  XNOR2_X1 DP_mult_207_U2195 ( .A(DP_pipe01[21]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1484) );
  XNOR2_X1 DP_mult_207_U2194 ( .A(DP_pipe01[19]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1486) );
  XNOR2_X1 DP_mult_207_U2193 ( .A(DP_pipe01[17]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1488) );
  XNOR2_X1 DP_mult_207_U2192 ( .A(DP_pipe01[15]), .B(DP_mult_207_n2317), .ZN(
        DP_mult_207_n1490) );
  XNOR2_X1 DP_mult_207_U2191 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2280), .ZN(
        DP_mult_207_n1698) );
  XNOR2_X1 DP_mult_207_U2190 ( .A(DP_mult_207_n2281), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1705) );
  XNOR2_X1 DP_mult_207_U2189 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2312), .ZN(
        DP_mult_207_n1507) );
  XNOR2_X1 DP_mult_207_U2188 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2309), .ZN(
        DP_mult_207_n1532) );
  XNOR2_X1 DP_mult_207_U2187 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2298), .ZN(
        DP_mult_207_n1582) );
  XNOR2_X1 DP_mult_207_U2186 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2057), .ZN(
        DP_mult_207_n1557) );
  XNOR2_X1 DP_mult_207_U2185 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2293), .ZN(
        DP_mult_207_n1607) );
  XNOR2_X1 DP_mult_207_U2184 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2270), .ZN(
        DP_mult_207_n1732) );
  XNOR2_X1 DP_mult_207_U2183 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2275), .ZN(
        DP_mult_207_n1707) );
  XNOR2_X1 DP_mult_207_U2182 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2280), .ZN(
        DP_mult_207_n1682) );
  XNOR2_X1 DP_mult_207_U2181 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2285), .ZN(
        DP_mult_207_n1657) );
  XNOR2_X1 DP_mult_207_U2180 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2016), .ZN(
        DP_mult_207_n1632) );
  XNOR2_X1 DP_mult_207_U2179 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2280), .ZN(
        DP_mult_207_n1696) );
  XNOR2_X1 DP_mult_207_U2178 ( .A(DP_mult_207_n2314), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1530) );
  XNOR2_X1 DP_mult_207_U2177 ( .A(DP_pipe01[23]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1757) );
  XNOR2_X1 DP_mult_207_U2176 ( .A(DP_pipe01[1]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1779) );
  XNOR2_X1 DP_mult_207_U2175 ( .A(DP_pipe01[5]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1775) );
  XNOR2_X1 DP_mult_207_U2174 ( .A(DP_pipe01[3]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1777) );
  XNOR2_X1 DP_mult_207_U2173 ( .A(DP_pipe01[7]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1773) );
  XNOR2_X1 DP_mult_207_U2172 ( .A(DP_pipe01[9]), .B(DP_mult_207_n2264), .ZN(
        DP_mult_207_n1771) );
  XNOR2_X1 DP_mult_207_U2171 ( .A(DP_mult_207_n2304), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1560) );
  XNOR2_X1 DP_mult_207_U2170 ( .A(DP_mult_207_n2300), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1583) );
  XNOR2_X1 DP_mult_207_U2169 ( .A(DP_mult_207_n2304), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1558) );
  XNOR2_X1 DP_mult_207_U2168 ( .A(DP_mult_207_n2303), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1570) );
  XNOR2_X1 DP_mult_207_U2167 ( .A(DP_mult_207_n2281), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1685) );
  XNOR2_X1 DP_mult_207_U2166 ( .A(DP_mult_207_n2290), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1639) );
  XNOR2_X1 DP_mult_207_U2165 ( .A(DP_mult_207_n2307), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1547) );
  XNOR2_X1 DP_mult_207_U2164 ( .A(DP_mult_207_n2277), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1708) );
  XNOR2_X1 DP_mult_207_U2163 ( .A(DP_mult_207_n2286), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1662) );
  XNOR2_X1 DP_mult_207_U2162 ( .A(DP_mult_207_n2313), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1524) );
  XNOR2_X1 DP_mult_207_U2161 ( .A(DP_mult_207_n2294), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1616) );
  XNOR2_X1 DP_mult_207_U2160 ( .A(DP_mult_207_n2299), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1591) );
  XNOR2_X1 DP_mult_207_U2159 ( .A(DP_mult_207_n2282), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1683) );
  XNOR2_X1 DP_mult_207_U2158 ( .A(DP_mult_207_n2308), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1545) );
  XNOR2_X1 DP_mult_207_U2157 ( .A(DP_mult_207_n2295), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1614) );
  XNOR2_X1 DP_mult_207_U2156 ( .A(DP_mult_207_n2290), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1637) );
  XNOR2_X1 DP_mult_207_U2155 ( .A(DP_mult_207_n2313), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1522) );
  XNOR2_X1 DP_mult_207_U2154 ( .A(DP_mult_207_n2281), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1687) );
  XNOR2_X1 DP_mult_207_U2153 ( .A(DP_mult_207_n2307), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1549) );
  XNOR2_X1 DP_mult_207_U2152 ( .A(DP_mult_207_n2287), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1664) );
  XNOR2_X1 DP_mult_207_U2151 ( .A(DP_mult_207_n2277), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1710) );
  XNOR2_X1 DP_mult_207_U2150 ( .A(DP_mult_207_n2299), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1593) );
  XNOR2_X1 DP_mult_207_U2149 ( .A(DP_mult_207_n2016), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1641) );
  XNOR2_X1 DP_mult_207_U2148 ( .A(DP_mult_207_n2299), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1595) );
  XNOR2_X1 DP_mult_207_U2147 ( .A(DP_mult_207_n2294), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1618) );
  XNOR2_X1 DP_mult_207_U2146 ( .A(DP_mult_207_n2303), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1572) );
  XNOR2_X1 DP_mult_207_U2145 ( .A(DP_mult_207_n2272), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1733) );
  XNOR2_X1 DP_mult_207_U2144 ( .A(DP_mult_207_n2303), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1568) );
  XNOR2_X1 DP_mult_207_U2143 ( .A(DP_mult_207_n2317), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1499) );
  XNOR2_X1 DP_mult_207_U2142 ( .A(DP_mult_207_n2287), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1660) );
  XNOR2_X1 DP_mult_207_U2141 ( .A(DP_mult_207_n2318), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1497) );
  XNOR2_X1 DP_mult_207_U2140 ( .A(DP_mult_207_n2271), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1749) );
  XNOR2_X1 DP_mult_207_U2139 ( .A(DP_mult_207_n2313), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1520) );
  XNOR2_X1 DP_mult_207_U2138 ( .A(DP_mult_207_n2294), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1612) );
  XNOR2_X1 DP_mult_207_U2137 ( .A(DP_mult_207_n2276), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1724) );
  XNOR2_X1 DP_mult_207_U2136 ( .A(DP_mult_207_n2276), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1722) );
  XNOR2_X1 DP_mult_207_U2135 ( .A(DP_mult_207_n2271), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1745) );
  XNOR2_X1 DP_mult_207_U2134 ( .A(DP_mult_207_n2287), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1658) );
  XNOR2_X1 DP_mult_207_U2133 ( .A(DP_mult_207_n2271), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1747) );
  XNOR2_X1 DP_mult_207_U2132 ( .A(DP_mult_207_n2276), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1720) );
  XNOR2_X1 DP_mult_207_U2131 ( .A(DP_mult_207_n2295), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1610) );
  XNOR2_X1 DP_mult_207_U2130 ( .A(DP_mult_207_n2303), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1566) );
  XNOR2_X1 DP_mult_207_U2129 ( .A(DP_mult_207_n2300), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1589) );
  XNOR2_X1 DP_mult_207_U2128 ( .A(DP_mult_207_n2290), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1635) );
  XNOR2_X1 DP_mult_207_U2127 ( .A(DP_mult_207_n2309), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1543) );
  XNOR2_X1 DP_mult_207_U2126 ( .A(DP_mult_207_n2282), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1697) );
  XNOR2_X1 DP_mult_207_U2125 ( .A(DP_mult_207_n2286), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1674) );
  XNOR2_X1 DP_mult_207_U2124 ( .A(DP_mult_207_n2271), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1743) );
  XNOR2_X1 DP_mult_207_U2123 ( .A(DP_mult_207_n2295), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1608) );
  XNOR2_X1 DP_mult_207_U2122 ( .A(DP_mult_207_n2272), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1735) );
  XNOR2_X1 DP_mult_207_U2121 ( .A(DP_mult_207_n2286), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1666) );
  XNOR2_X1 DP_mult_207_U2120 ( .A(DP_mult_207_n2299), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1597) );
  XNOR2_X1 DP_mult_207_U2119 ( .A(DP_mult_207_n2015), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1643) );
  XNOR2_X1 DP_mult_207_U2118 ( .A(DP_mult_207_n2303), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1574) );
  XNOR2_X1 DP_mult_207_U2117 ( .A(DP_mult_207_n2294), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1620) );
  XNOR2_X1 DP_mult_207_U2116 ( .A(DP_mult_207_n2290), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1633) );
  XNOR2_X1 DP_mult_207_U2115 ( .A(DP_mult_207_n2300), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1585) );
  XNOR2_X1 DP_mult_207_U2114 ( .A(DP_mult_207_n2276), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1712) );
  XNOR2_X1 DP_mult_207_U2113 ( .A(DP_mult_207_n2015), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1645) );
  XNOR2_X1 DP_mult_207_U2112 ( .A(DP_mult_207_n2317), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1493) );
  XNOR2_X1 DP_mult_207_U2111 ( .A(DP_mult_207_n2294), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1622) );
  XNOR2_X1 DP_mult_207_U2110 ( .A(DP_mult_207_n2286), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1668) );
  XNOR2_X1 DP_mult_207_U2109 ( .A(DP_mult_207_n2277), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1714) );
  XNOR2_X1 DP_mult_207_U2108 ( .A(DP_mult_207_n2299), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1599) );
  XNOR2_X1 DP_mult_207_U2107 ( .A(DP_mult_207_n2294), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1624) );
  XNOR2_X1 DP_mult_207_U2106 ( .A(DP_mult_207_n2281), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1689) );
  XNOR2_X1 DP_mult_207_U2105 ( .A(DP_mult_207_n2282), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1693) );
  XNOR2_X1 DP_mult_207_U2104 ( .A(DP_mult_207_n2015), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1647) );
  XNOR2_X1 DP_mult_207_U2103 ( .A(DP_mult_207_n2276), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1716) );
  XNOR2_X1 DP_mult_207_U2102 ( .A(DP_mult_207_n2272), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1739) );
  XNOR2_X1 DP_mult_207_U2101 ( .A(DP_mult_207_n2276), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1718) );
  XNOR2_X1 DP_mult_207_U2100 ( .A(DP_mult_207_n2286), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1670) );
  XNOR2_X1 DP_mult_207_U2099 ( .A(DP_mult_207_n2304), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1564) );
  XNOR2_X1 DP_mult_207_U2098 ( .A(DP_mult_207_n2299), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1587) );
  XNOR2_X1 DP_mult_207_U2097 ( .A(DP_mult_207_n2303), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1562) );
  XNOR2_X1 DP_mult_207_U2096 ( .A(DP_mult_207_n2286), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1672) );
  XNOR2_X1 DP_mult_207_U2095 ( .A(DP_mult_207_n2317), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1495) );
  XNOR2_X1 DP_mult_207_U2094 ( .A(DP_mult_207_n2290), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1649) );
  XNOR2_X1 DP_mult_207_U2093 ( .A(DP_mult_207_n2271), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1741) );
  XNOR2_X1 DP_mult_207_U2092 ( .A(DP_mult_207_n2271), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1737) );
  XNOR2_X1 DP_mult_207_U2091 ( .A(DP_mult_207_n2282), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1691) );
  XNOR2_X1 DP_mult_207_U2090 ( .A(DP_mult_207_n2313), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1518) );
  XNOR2_X1 DP_mult_207_U2089 ( .A(DP_mult_207_n2271), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1753) );
  XNOR2_X1 DP_mult_207_U2088 ( .A(DP_mult_207_n2318), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1501) );
  XNOR2_X1 DP_mult_207_U2087 ( .A(DP_mult_207_n2271), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1751) );
  XNOR2_X1 DP_mult_207_U2086 ( .A(DP_mult_207_n2276), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1728) );
  XNOR2_X1 DP_mult_207_U2085 ( .A(DP_mult_207_n2313), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1526) );
  XNOR2_X1 DP_mult_207_U2084 ( .A(DP_mult_207_n2318), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1503) );
  XNOR2_X1 DP_mult_207_U2083 ( .A(DP_mult_207_n2281), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1703) );
  XNOR2_X1 DP_mult_207_U2082 ( .A(DP_mult_207_n2286), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1676) );
  XNOR2_X1 DP_mult_207_U2081 ( .A(DP_mult_207_n2290), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1653) );
  XNOR2_X1 DP_mult_207_U2080 ( .A(DP_mult_207_n2286), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1678) );
  XNOR2_X1 DP_mult_207_U2079 ( .A(DP_mult_207_n2276), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1726) );
  XNOR2_X1 DP_mult_207_U2078 ( .A(DP_mult_207_n2281), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1701) );
  XNOR2_X1 DP_mult_207_U2077 ( .A(DP_mult_207_n2016), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1651) );
  XNOR2_X1 DP_mult_207_U2076 ( .A(DP_mult_207_n2313), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1528) );
  XNOR2_X1 DP_mult_207_U2075 ( .A(DP_mult_207_n2307), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1553) );
  XNOR2_X1 DP_mult_207_U2074 ( .A(DP_mult_207_n2308), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1551) );
  XNOR2_X1 DP_mult_207_U2073 ( .A(DP_mult_207_n2303), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1576) );
  XNOR2_X1 DP_mult_207_U2072 ( .A(DP_mult_207_n2299), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1603) );
  XNOR2_X1 DP_mult_207_U2071 ( .A(DP_mult_207_n2303), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1578) );
  XNOR2_X1 DP_mult_207_U2070 ( .A(DP_mult_207_n2299), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1601) );
  XNOR2_X1 DP_mult_207_U2069 ( .A(DP_mult_207_n2294), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1626) );
  XNOR2_X1 DP_mult_207_U2068 ( .A(DP_mult_207_n2294), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1628) );
  XNOR2_X1 DP_mult_207_U2067 ( .A(DP_mult_207_n2309), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1535) );
  XNOR2_X1 DP_mult_207_U2066 ( .A(DP_mult_207_n2314), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1510) );
  XNOR2_X1 DP_mult_207_U2065 ( .A(DP_mult_207_n2314), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1508) );
  XNOR2_X1 DP_mult_207_U2064 ( .A(DP_mult_207_n2308), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1533) );
  XNOR2_X1 DP_mult_207_U2063 ( .A(DP_mult_207_n2314), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1514) );
  XNOR2_X1 DP_mult_207_U2062 ( .A(DP_mult_207_n2313), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1512) );
  XNOR2_X1 DP_mult_207_U2061 ( .A(DP_mult_207_n2308), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1537) );
  XNOR2_X1 DP_mult_207_U2060 ( .A(DP_mult_207_n2308), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1541) );
  XNOR2_X1 DP_mult_207_U2059 ( .A(DP_mult_207_n2308), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1539) );
  XNOR2_X1 DP_mult_207_U2058 ( .A(DP_mult_207_n2313), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1516) );
  XNOR2_X1 DP_mult_207_U2057 ( .A(DP_mult_207_n2281), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1695) );
  XNOR2_X1 DP_mult_207_U2056 ( .A(DP_mult_207_n2317), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1491) );
  XNOR2_X1 DP_mult_207_U2055 ( .A(DP_mult_207_n2281), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1699) );
  XNOR2_X1 DP_mult_207_U2054 ( .A(DP_mult_207_n2265), .B(DP_pipe01[6]), .ZN(
        DP_mult_207_n1774) );
  XNOR2_X1 DP_mult_207_U2053 ( .A(DP_mult_207_n2265), .B(DP_pipe01[10]), .ZN(
        DP_mult_207_n1770) );
  XNOR2_X1 DP_mult_207_U2052 ( .A(DP_mult_207_n2265), .B(DP_pipe01[12]), .ZN(
        DP_mult_207_n1768) );
  XNOR2_X1 DP_mult_207_U2051 ( .A(DP_mult_207_n2265), .B(DP_pipe01[8]), .ZN(
        DP_mult_207_n1772) );
  XNOR2_X1 DP_mult_207_U2050 ( .A(DP_mult_207_n2265), .B(DP_pipe01[14]), .ZN(
        DP_mult_207_n1766) );
  XNOR2_X1 DP_mult_207_U2049 ( .A(DP_mult_207_n2266), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1758) );
  XNOR2_X1 DP_mult_207_U2048 ( .A(DP_mult_207_n2266), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1760) );
  XNOR2_X1 DP_mult_207_U2047 ( .A(DP_mult_207_n2265), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1762) );
  XNOR2_X1 DP_mult_207_U2046 ( .A(DP_mult_207_n2266), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1764) );
  XNOR2_X1 DP_mult_207_U2045 ( .A(DP_mult_207_n2317), .B(DP_pipe01[22]), .ZN(
        DP_mult_207_n1483) );
  XNOR2_X1 DP_mult_207_U2044 ( .A(DP_mult_207_n2317), .B(DP_pipe01[20]), .ZN(
        DP_mult_207_n1485) );
  XNOR2_X1 DP_mult_207_U2043 ( .A(DP_mult_207_n2317), .B(DP_pipe01[18]), .ZN(
        DP_mult_207_n1487) );
  XNOR2_X1 DP_mult_207_U2042 ( .A(DP_mult_207_n2317), .B(DP_pipe01[16]), .ZN(
        DP_mult_207_n1489) );
  XNOR2_X1 DP_mult_207_U2041 ( .A(DP_mult_207_n2265), .B(DP_pipe01[4]), .ZN(
        DP_mult_207_n1776) );
  XNOR2_X1 DP_mult_207_U2040 ( .A(DP_mult_207_n2265), .B(DP_pipe01[2]), .ZN(
        DP_mult_207_n1778) );
  XNOR2_X1 DP_mult_207_U2039 ( .A(DP_mult_207_n2287), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1680) );
  XNOR2_X1 DP_mult_207_U2038 ( .A(DP_mult_207_n2304), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1580) );
  XNOR2_X1 DP_mult_207_U2037 ( .A(DP_mult_207_n2309), .B(DP_pipe01[0]), .ZN(
        DP_mult_207_n1555) );
  INV_X1 DP_mult_207_U2036 ( .A(DP_mult_207_n1482), .ZN(DP_mult_207_n2331) );
  INV_X1 DP_mult_207_U2035 ( .A(DP_mult_207_n1732), .ZN(DP_mult_207_n2321) );
  INV_X1 DP_mult_207_U2034 ( .A(DP_mult_207_n1657), .ZN(DP_mult_207_n2324) );
  INV_X1 DP_mult_207_U2033 ( .A(DP_mult_207_n1582), .ZN(DP_mult_207_n2327) );
  OAI22_X1 DP_mult_207_U2032 ( .A1(DP_mult_207_n2095), .A2(DP_mult_207_n1489), 
        .B1(DP_mult_207_n1488), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n1200)
         );
  OAI22_X1 DP_mult_207_U2031 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1538), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1537), .ZN(DP_mult_207_n1247)
         );
  OAI22_X1 DP_mult_207_U2030 ( .A1(DP_mult_207_n2096), .A2(DP_mult_207_n1491), 
        .B1(DP_mult_207_n1490), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n1202)
         );
  INV_X1 DP_mult_207_U2029 ( .A(DP_mult_207_n1607), .ZN(DP_mult_207_n2326) );
  INV_X1 DP_mult_207_U2028 ( .A(DP_mult_207_n1557), .ZN(DP_mult_207_n2328) );
  OAI22_X1 DP_mult_207_U2027 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1534), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1533), .ZN(DP_mult_207_n1243)
         );
  OAI21_X1 DP_mult_207_U2026 ( .B1(DP_mult_207_n2187), .B2(DP_mult_207_n2130), 
        .A(DP_mult_207_n2328), .ZN(DP_mult_207_n1266) );
  INV_X1 DP_mult_207_U2025 ( .A(DP_mult_207_n874), .ZN(DP_mult_207_n875) );
  OAI22_X1 DP_mult_207_U2024 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1773), 
        .B1(DP_mult_207_n1772), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1474)
         );
  OAI22_X1 DP_mult_207_U2023 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1762), 
        .B1(DP_mult_207_n1761), .B2(DP_mult_207_n2262), .ZN(DP_mult_207_n1463)
         );
  OAI22_X1 DP_mult_207_U2022 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1758), 
        .B1(DP_mult_207_n1757), .B2(DP_mult_207_n2262), .ZN(DP_mult_207_n1459)
         );
  OAI22_X1 DP_mult_207_U2021 ( .A1(DP_mult_207_n2114), .A2(DP_mult_207_n1699), 
        .B1(DP_mult_207_n1698), .B2(DP_mult_207_n2255), .ZN(DP_mult_207_n1402)
         );
  NOR2_X1 DP_mult_207_U2020 ( .A1(DP_mult_207_n2246), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1337) );
  NOR2_X1 DP_mult_207_U2019 ( .A1(DP_mult_207_n2241), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1289) );
  INV_X1 DP_mult_207_U2018 ( .A(DP_mult_207_n1707), .ZN(DP_mult_207_n2322) );
  OAI21_X1 DP_mult_207_U2017 ( .B1(DP_mult_207_n2190), .B2(DP_mult_207_n2066), 
        .A(DP_mult_207_n2322), .ZN(DP_mult_207_n1410) );
  INV_X1 DP_mult_207_U2016 ( .A(DP_mult_207_n802), .ZN(DP_mult_207_n803) );
  NOR2_X1 DP_mult_207_U2015 ( .A1(DP_mult_207_n2239), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1241) );
  OAI22_X1 DP_mult_207_U2014 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1509), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1508), .ZN(DP_mult_207_n1219)
         );
  OAI22_X1 DP_mult_207_U2013 ( .A1(DP_mult_207_n2096), .A2(DP_mult_207_n1486), 
        .B1(DP_mult_207_n2238), .B2(DP_mult_207_n1485), .ZN(DP_mult_207_n1197)
         );
  OAI22_X1 DP_mult_207_U2012 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1766), 
        .B1(DP_mult_207_n1765), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1467)
         );
  NOR2_X1 DP_mult_207_U2011 ( .A1(DP_mult_207_n2077), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1265) );
  OAI22_X1 DP_mult_207_U2010 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1759), 
        .B1(DP_mult_207_n1758), .B2(DP_mult_207_n2262), .ZN(DP_mult_207_n1460)
         );
  OAI22_X1 DP_mult_207_U2009 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1775), 
        .B1(DP_mult_207_n1774), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1476)
         );
  OAI22_X1 DP_mult_207_U2008 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1771), 
        .B1(DP_mult_207_n1770), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1472)
         );
  OAI22_X1 DP_mult_207_U2007 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1772), 
        .B1(DP_mult_207_n1771), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1473)
         );
  INV_X1 DP_mult_207_U2006 ( .A(DP_mult_207_n1682), .ZN(DP_mult_207_n2323) );
  OAI21_X1 DP_mult_207_U2005 ( .B1(DP_mult_207_n2191), .B2(DP_mult_207_n1930), 
        .A(DP_mult_207_n2323), .ZN(DP_mult_207_n1386) );
  OAI22_X1 DP_mult_207_U2004 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1517), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1516), .ZN(DP_mult_207_n1227)
         );
  OAI22_X1 DP_mult_207_U2003 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1774), 
        .B1(DP_mult_207_n1773), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1475)
         );
  OAI22_X1 DP_mult_207_U2002 ( .A1(DP_mult_207_n2229), .A2(DP_mult_207_n1696), 
        .B1(DP_mult_207_n2255), .B2(DP_mult_207_n1695), .ZN(DP_mult_207_n1399)
         );
  OAI22_X1 DP_mult_207_U2001 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1770), 
        .B1(DP_mult_207_n1769), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1471)
         );
  OAI22_X1 DP_mult_207_U2000 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1769), 
        .B1(DP_mult_207_n1768), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1470)
         );
  NOR2_X1 DP_mult_207_U1999 ( .A1(DP_mult_207_n2250), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1361) );
  NOR2_X1 DP_mult_207_U1998 ( .A1(DP_mult_207_n1991), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1313) );
  OAI22_X1 DP_mult_207_U1997 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1763), 
        .B1(DP_mult_207_n1762), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1464)
         );
  NOR2_X1 DP_mult_207_U1996 ( .A1(DP_mult_207_n2238), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1217) );
  OAI22_X1 DP_mult_207_U1995 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1768), 
        .B1(DP_mult_207_n1767), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1469)
         );
  OAI22_X1 DP_mult_207_U1994 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1515), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1514), .ZN(DP_mult_207_n1225)
         );
  OAI22_X1 DP_mult_207_U1993 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1761), 
        .B1(DP_mult_207_n1760), .B2(DP_mult_207_n2262), .ZN(DP_mult_207_n1462)
         );
  OAI22_X1 DP_mult_207_U1992 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1767), 
        .B1(DP_mult_207_n1766), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1468)
         );
  OAI22_X1 DP_mult_207_U1991 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1542), 
        .B1(DP_mult_207_n2077), .B2(DP_mult_207_n1541), .ZN(DP_mult_207_n1251)
         );
  OAI22_X1 DP_mult_207_U1990 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1513), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1512), .ZN(DP_mult_207_n1223)
         );
  OAI22_X1 DP_mult_207_U1989 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1536), 
        .B1(DP_mult_207_n2140), .B2(DP_mult_207_n1535), .ZN(DP_mult_207_n1245)
         );
  OAI21_X1 DP_mult_207_U1988 ( .B1(DP_mult_207_n2189), .B2(DP_mult_207_n2244), 
        .A(DP_mult_207_n2327), .ZN(DP_mult_207_n1290) );
  INV_X1 DP_mult_207_U1987 ( .A(DP_mult_207_n1532), .ZN(DP_mult_207_n2329) );
  OAI21_X1 DP_mult_207_U1986 ( .B1(DP_mult_207_n1984), .B2(DP_mult_207_n2186), 
        .A(DP_mult_207_n2329), .ZN(DP_mult_207_n1242) );
  OAI22_X1 DP_mult_207_U1985 ( .A1(DP_mult_207_n2096), .A2(DP_mult_207_n1490), 
        .B1(DP_mult_207_n2238), .B2(DP_mult_207_n1489), .ZN(DP_mult_207_n1201)
         );
  OAI22_X1 DP_mult_207_U1984 ( .A1(DP_mult_207_n2218), .A2(DP_mult_207_n1540), 
        .B1(DP_mult_207_n2077), .B2(DP_mult_207_n1539), .ZN(DP_mult_207_n1249)
         );
  OAI22_X1 DP_mult_207_U1983 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1760), 
        .B1(DP_mult_207_n1759), .B2(DP_mult_207_n2262), .ZN(DP_mult_207_n1461)
         );
  INV_X1 DP_mult_207_U1982 ( .A(DP_mult_207_n1632), .ZN(DP_mult_207_n2325) );
  OAI22_X1 DP_mult_207_U1981 ( .A1(DP_mult_207_n2095), .A2(DP_mult_207_n1487), 
        .B1(DP_mult_207_n1486), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n1198)
         );
  INV_X1 DP_mult_207_U1980 ( .A(DP_mult_207_n692), .ZN(DP_mult_207_n693) );
  INV_X1 DP_mult_207_U1979 ( .A(DP_mult_207_n724), .ZN(DP_mult_207_n725) );
  CLKBUF_X1 DP_mult_207_U1978 ( .A(DP_mult_207_n251), .Z(DP_mult_207_n2262) );
  NOR2_X1 DP_mult_207_U1977 ( .A1(DP_mult_207_n1181), .A2(DP_mult_207_n1192), 
        .ZN(DP_mult_207_n644) );
  NAND2_X1 DP_mult_207_U1976 ( .A1(DP_mult_207_n1181), .A2(DP_mult_207_n1192), 
        .ZN(DP_mult_207_n645) );
  NAND2_X1 DP_mult_207_U1975 ( .A1(DP_mult_207_n2265), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1781) );
  NAND2_X1 DP_mult_207_U1974 ( .A1(DP_mult_207_n2281), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1706) );
  NAND2_X1 DP_mult_207_U1973 ( .A1(DP_mult_207_n2294), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1631) );
  NAND2_X1 DP_mult_207_U1972 ( .A1(DP_mult_207_n2015), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1656) );
  NAND2_X1 DP_mult_207_U1971 ( .A1(DP_mult_207_n2286), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1681) );
  NAND2_X1 DP_mult_207_U1970 ( .A1(DP_mult_207_n2317), .A2(DP_mult_207_n2012), 
        .ZN(DP_mult_207_n1506) );
  NAND2_X1 DP_mult_207_U1969 ( .A1(DP_mult_207_n2299), .A2(DP_mult_207_n2012), 
        .ZN(DP_mult_207_n1606) );
  NAND2_X1 DP_mult_207_U1968 ( .A1(DP_mult_207_n2313), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1531) );
  NAND2_X1 DP_mult_207_U1967 ( .A1(DP_mult_207_n2309), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1556) );
  NAND2_X1 DP_mult_207_U1966 ( .A1(DP_mult_207_n2303), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1581) );
  AOI21_X1 DP_mult_207_U1965 ( .B1(DP_mult_207_n1965), .B2(DP_mult_207_n1964), 
        .A(DP_mult_207_n1972), .ZN(DP_mult_207_n646) );
  INV_X2 DP_mult_207_U1964 ( .A(DP_mult_207_n2267), .ZN(DP_mult_207_n2264) );
  OAI22_X1 DP_mult_207_U1963 ( .A1(DP_mult_207_n2095), .A2(DP_mult_207_n1488), 
        .B1(DP_mult_207_n2238), .B2(DP_mult_207_n1487), .ZN(DP_mult_207_n1199)
         );
  OAI22_X1 DP_mult_207_U1962 ( .A1(DP_mult_207_n2216), .A2(DP_mult_207_n1511), 
        .B1(DP_mult_207_n2239), .B2(DP_mult_207_n1510), .ZN(DP_mult_207_n1221)
         );
  NOR2_X1 DP_mult_207_U1961 ( .A1(DP_mult_207_n2255), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1409) );
  NOR2_X1 DP_mult_207_U1960 ( .A1(DP_mult_207_n2253), .A2(DP_mult_207_n2014), 
        .ZN(DP_mult_207_n1385) );
  INV_X1 DP_mult_207_U1959 ( .A(DP_mult_207_n682), .ZN(DP_mult_207_n683) );
  OAI22_X1 DP_mult_207_U1958 ( .A1(DP_mult_207_n2095), .A2(DP_mult_207_n1485), 
        .B1(DP_mult_207_n1484), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n1196)
         );
  OAI22_X1 DP_mult_207_U1957 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1777), 
        .B1(DP_mult_207_n1776), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1478)
         );
  NAND2_X1 DP_mult_207_U1956 ( .A1(DP_mult_207_n2276), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1731) );
  INV_X1 DP_mult_207_U1955 ( .A(DP_mult_207_n1507), .ZN(DP_mult_207_n2330) );
  OAI22_X1 DP_mult_207_U1954 ( .A1(DP_mult_207_n2096), .A2(DP_mult_207_n1484), 
        .B1(DP_mult_207_n2238), .B2(DP_mult_207_n1483), .ZN(DP_mult_207_n1195)
         );
  OAI22_X1 DP_mult_207_U1953 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1764), 
        .B1(DP_mult_207_n1763), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1465)
         );
  OAI22_X1 DP_mult_207_U1952 ( .A1(DP_mult_207_n2236), .A2(DP_mult_207_n1765), 
        .B1(DP_mult_207_n1764), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1466)
         );
  INV_X1 DP_mult_207_U1951 ( .A(DP_mult_207_n1984), .ZN(DP_mult_207_n2218) );
  INV_X1 DP_mult_207_U1950 ( .A(DP_mult_207_n2194), .ZN(DP_mult_207_n2216) );
  NOR2_X1 DP_mult_207_U1949 ( .A1(DP_mult_207_n2259), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1457) );
  NOR2_X1 DP_mult_207_U1948 ( .A1(DP_mult_207_n2257), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1433) );
  OAI22_X1 DP_mult_207_U1947 ( .A1(DP_mult_207_n2235), .A2(DP_mult_207_n1779), 
        .B1(DP_mult_207_n1778), .B2(DP_mult_207_n2261), .ZN(DP_mult_207_n1480)
         );
  OAI22_X1 DP_mult_207_U1946 ( .A1(DP_mult_207_n2095), .A2(DP_mult_207_n1483), 
        .B1(DP_mult_207_n1482), .B2(DP_mult_207_n1937), .ZN(DP_mult_207_n676)
         );
  NAND2_X1 DP_mult_207_U1945 ( .A1(DP_mult_207_n2271), .A2(DP_mult_207_n2013), 
        .ZN(DP_mult_207_n1756) );
  OR2_X1 DP_mult_207_U1944 ( .A1(DP_mult_207_n1194), .A2(DP_mult_207_n676), 
        .ZN(DP_mult_207_n2183) );
  NAND2_X1 DP_mult_207_U1943 ( .A1(DP_mult_207_n678), .A2(DP_mult_207_n677), 
        .ZN(DP_mult_207_n335) );
  NAND2_X1 DP_mult_207_U1942 ( .A1(DP_mult_207_n1171), .A2(DP_mult_207_n1174), 
        .ZN(DP_mult_207_n634) );
  NAND2_X1 DP_mult_207_U1941 ( .A1(DP_mult_207_n1175), .A2(DP_mult_207_n1178), 
        .ZN(DP_mult_207_n637) );
  NAND2_X1 DP_mult_207_U1940 ( .A1(DP_mult_207_n1165), .A2(DP_mult_207_n1170), 
        .ZN(DP_mult_207_n632) );
  NAND2_X1 DP_mult_207_U1939 ( .A1(DP_mult_207_n1159), .A2(DP_mult_207_n1161), 
        .ZN(DP_mult_207_n627) );
  NOR2_X1 DP_mult_207_U1938 ( .A1(DP_mult_207_n1175), .A2(DP_mult_207_n1178), 
        .ZN(DP_mult_207_n636) );
  NOR2_X1 DP_mult_207_U1937 ( .A1(DP_mult_207_n1171), .A2(DP_mult_207_n1174), 
        .ZN(DP_mult_207_n633) );
  NAND2_X1 DP_mult_207_U1936 ( .A1(DP_mult_207_n679), .A2(DP_mult_207_n680), 
        .ZN(DP_mult_207_n341) );
  NAND2_X1 DP_mult_207_U1935 ( .A1(DP_mult_207_n681), .A2(DP_mult_207_n684), 
        .ZN(DP_mult_207_n352) );
  OR2_X1 DP_mult_207_U1934 ( .A1(DP_mult_207_n679), .A2(DP_mult_207_n680), 
        .ZN(DP_mult_207_n2182) );
  NOR2_X1 DP_mult_207_U1933 ( .A1(DP_mult_207_n1159), .A2(DP_mult_207_n1161), 
        .ZN(DP_mult_207_n626) );
  OR2_X1 DP_mult_207_U1932 ( .A1(DP_mult_207_n681), .A2(DP_mult_207_n684), 
        .ZN(DP_mult_207_n2181) );
  NOR2_X1 DP_mult_207_U1931 ( .A1(DP_mult_207_n1165), .A2(DP_mult_207_n1170), 
        .ZN(DP_mult_207_n631) );
  NOR2_X1 DP_mult_207_U1930 ( .A1(DP_mult_207_n678), .A2(DP_mult_207_n677), 
        .ZN(DP_mult_207_n334) );
  OAI21_X1 DP_mult_207_U1929 ( .B1(DP_mult_207_n646), .B2(DP_mult_207_n644), 
        .A(DP_mult_207_n645), .ZN(DP_mult_207_n643) );
  AOI21_X1 DP_mult_207_U1928 ( .B1(DP_mult_207_n643), .B2(DP_mult_207_n1967), 
        .A(DP_mult_207_n1974), .ZN(DP_mult_207_n638) );
  OR2_X1 DP_mult_207_U1927 ( .A1(DP_mult_207_n685), .A2(DP_mult_207_n688), 
        .ZN(DP_mult_207_n2180) );
  INV_X1 DP_mult_207_U1926 ( .A(DP_mult_207_n676), .ZN(DP_mult_207_n677) );
  AND2_X1 DP_mult_207_U1925 ( .A1(DP_mult_207_n1194), .A2(DP_mult_207_n676), 
        .ZN(DP_mult_207_n2179) );
  NOR2_X1 DP_mult_207_U1924 ( .A1(DP_mult_207_n590), .A2(DP_mult_207_n592), 
        .ZN(DP_mult_207_n588) );
  NAND2_X1 DP_mult_207_U1923 ( .A1(DP_mult_207_n588), .A2(DP_mult_207_n2166), 
        .ZN(DP_mult_207_n582) );
  AOI21_X1 DP_mult_207_U1922 ( .B1(DP_mult_207_n2176), .B2(DP_mult_207_n1969), 
        .A(DP_mult_207_n1977), .ZN(DP_mult_207_n600) );
  NAND2_X1 DP_mult_207_U1921 ( .A1(DP_mult_207_n1979), .A2(DP_mult_207_n2175), 
        .ZN(DP_mult_207_n610) );
  OR2_X1 DP_mult_207_U1920 ( .A1(DP_mult_207_n694), .A2(DP_mult_207_n689), 
        .ZN(DP_mult_207_n2178) );
  NAND2_X1 DP_mult_207_U1919 ( .A1(DP_mult_207_n709), .A2(DP_mult_207_n716), 
        .ZN(DP_mult_207_n409) );
  INV_X1 DP_mult_207_U1918 ( .A(DP_mult_207_n369), .ZN(DP_mult_207_n367) );
  OR2_X1 DP_mult_207_U1917 ( .A1(DP_mult_207_n709), .A2(DP_mult_207_n716), 
        .ZN(DP_mult_207_n2177) );
  NAND2_X1 DP_mult_207_U1916 ( .A1(DP_mult_207_n727), .A2(DP_mult_207_n736), 
        .ZN(DP_mult_207_n429) );
  NAND2_X1 DP_mult_207_U1915 ( .A1(DP_mult_207_n695), .A2(DP_mult_207_n700), 
        .ZN(DP_mult_207_n387) );
  OR2_X1 DP_mult_207_U1914 ( .A1(DP_mult_207_n1111), .A2(DP_mult_207_n1122), 
        .ZN(DP_mult_207_n2176) );
  OAI21_X1 DP_mult_207_U1913 ( .B1(DP_mult_207_n628), .B2(DP_mult_207_n626), 
        .A(DP_mult_207_n627), .ZN(DP_mult_207_n625) );
  AOI21_X1 DP_mult_207_U1912 ( .B1(DP_mult_207_n625), .B2(DP_mult_207_n1978), 
        .A(DP_mult_207_n1970), .ZN(DP_mult_207_n620) );
  AOI21_X1 DP_mult_207_U1911 ( .B1(DP_mult_207_n2175), .B2(DP_mult_207_n1968), 
        .A(DP_mult_207_n1976), .ZN(DP_mult_207_n611) );
  OR2_X1 DP_mult_207_U1910 ( .A1(DP_mult_207_n1133), .A2(DP_mult_207_n1142), 
        .ZN(DP_mult_207_n2175) );
  NAND2_X1 DP_mult_207_U1909 ( .A1(DP_mult_207_n2182), .A2(DP_mult_207_n341), 
        .ZN(DP_mult_207_n302) );
  NAND2_X1 DP_mult_207_U1908 ( .A1(DP_mult_207_n2181), .A2(DP_mult_207_n352), 
        .ZN(DP_mult_207_n303) );
  OR2_X1 DP_mult_207_U1907 ( .A1(DP_mult_207_n1123), .A2(DP_mult_207_n1132), 
        .ZN(DP_mult_207_n2174) );
  NAND2_X1 DP_mult_207_U1906 ( .A1(DP_mult_207_n2180), .A2(DP_mult_207_n369), 
        .ZN(DP_mult_207_n304) );
  INV_X1 DP_mult_207_U1905 ( .A(DP_mult_207_n341), .ZN(DP_mult_207_n339) );
  NOR2_X1 DP_mult_207_U1904 ( .A1(DP_mult_207_n727), .A2(DP_mult_207_n736), 
        .ZN(DP_mult_207_n428) );
  XNOR2_X1 DP_mult_207_U1903 ( .A(DP_mult_207_n920), .B(DP_mult_207_n901), 
        .ZN(DP_mult_207_n2173) );
  XNOR2_X1 DP_mult_207_U1902 ( .A(DP_mult_207_n2173), .B(DP_mult_207_n899), 
        .ZN(DP_mult_207_n897) );
  OR2_X1 DP_mult_207_U1901 ( .A1(DP_mult_207_n701), .A2(DP_mult_207_n708), 
        .ZN(DP_mult_207_n2172) );
  AOI21_X1 DP_mult_207_U1900 ( .B1(DP_mult_207_n376), .B2(DP_mult_207_n2180), 
        .A(DP_mult_207_n367), .ZN(DP_mult_207_n365) );
  OAI21_X1 DP_mult_207_U1899 ( .B1(DP_mult_207_n364), .B2(DP_mult_207_n387), 
        .A(DP_mult_207_n365), .ZN(DP_mult_207_n363) );
  AOI21_X1 DP_mult_207_U1898 ( .B1(DP_mult_207_n362), .B2(DP_mult_207_n394), 
        .A(DP_mult_207_n363), .ZN(DP_mult_207_n361) );
  INV_X1 DP_mult_207_U1897 ( .A(DP_mult_207_n352), .ZN(DP_mult_207_n350) );
  OR2_X1 DP_mult_207_U1896 ( .A1(DP_mult_207_n717), .A2(DP_mult_207_n726), 
        .ZN(DP_mult_207_n2171) );
  NOR2_X1 DP_mult_207_U1895 ( .A1(DP_mult_207_n695), .A2(DP_mult_207_n700), 
        .ZN(DP_mult_207_n384) );
  OR2_X1 DP_mult_207_U1894 ( .A1(DP_mult_207_n1039), .A2(DP_mult_207_n1054), 
        .ZN(DP_mult_207_n2170) );
  NAND2_X1 DP_mult_207_U1893 ( .A1(DP_mult_207_n400), .A2(DP_mult_207_n2172), 
        .ZN(DP_mult_207_n389) );
  NAND2_X1 DP_mult_207_U1892 ( .A1(DP_mult_207_n983), .A2(DP_mult_207_n1002), 
        .ZN(DP_mult_207_n564) );
  NOR2_X1 DP_mult_207_U1891 ( .A1(DP_mult_207_n389), .A2(DP_mult_207_n384), 
        .ZN(DP_mult_207_n382) );
  INV_X1 DP_mult_207_U1890 ( .A(DP_mult_207_n378), .ZN(DP_mult_207_n376) );
  NAND2_X1 DP_mult_207_U1889 ( .A1(DP_mult_207_n941), .A2(DP_mult_207_n962), 
        .ZN(DP_mult_207_n550) );
  NAND2_X1 DP_mult_207_U1888 ( .A1(DP_mult_207_n857), .A2(DP_mult_207_n876), 
        .ZN(DP_mult_207_n521) );
  OR2_X1 DP_mult_207_U1887 ( .A1(DP_mult_207_n761), .A2(DP_mult_207_n774), 
        .ZN(DP_mult_207_n2168) );
  INV_X1 DP_mult_207_U1886 ( .A(DP_mult_207_n418), .ZN(DP_mult_207_n416) );
  OAI21_X1 DP_mult_207_U1885 ( .B1(DP_mult_207_n590), .B2(DP_mult_207_n593), 
        .A(DP_mult_207_n591), .ZN(DP_mult_207_n589) );
  AOI21_X1 DP_mult_207_U1884 ( .B1(DP_mult_207_n589), .B2(DP_mult_207_n2166), 
        .A(DP_mult_207_n1975), .ZN(DP_mult_207_n583) );
  AOI21_X1 DP_mult_207_U1883 ( .B1(DP_mult_207_n423), .B2(DP_mult_207_n2171), 
        .A(DP_mult_207_n416), .ZN(DP_mult_207_n412) );
  OR2_X1 DP_mult_207_U1882 ( .A1(DP_mult_207_n788), .A2(DP_mult_207_n775), 
        .ZN(DP_mult_207_n2167) );
  NOR2_X1 DP_mult_207_U1881 ( .A1(DP_mult_207_n1003), .A2(DP_mult_207_n1020), 
        .ZN(DP_mult_207_n569) );
  OAI21_X1 DP_mult_207_U1880 ( .B1(DP_mult_207_n600), .B2(DP_mult_207_n597), 
        .A(DP_mult_207_n598), .ZN(DP_mult_207_n596) );
  OAI21_X1 DP_mult_207_U1879 ( .B1(DP_mult_207_n620), .B2(DP_mult_207_n610), 
        .A(DP_mult_207_n611), .ZN(DP_mult_207_n609) );
  NOR2_X1 DP_mult_207_U1878 ( .A1(DP_mult_207_n597), .A2(DP_mult_207_n599), 
        .ZN(DP_mult_207_n595) );
  AOI21_X1 DP_mult_207_U1877 ( .B1(DP_mult_207_n595), .B2(DP_mult_207_n609), 
        .A(DP_mult_207_n596), .ZN(DP_mult_207_n594) );
  NAND2_X1 DP_mult_207_U1876 ( .A1(DP_mult_207_n2171), .A2(DP_mult_207_n2177), 
        .ZN(DP_mult_207_n402) );
  NOR2_X1 DP_mult_207_U1875 ( .A1(DP_mult_207_n983), .A2(DP_mult_207_n1002), 
        .ZN(DP_mult_207_n563) );
  AOI21_X1 DP_mult_207_U1874 ( .B1(DP_mult_207_n401), .B2(DP_mult_207_n2172), 
        .A(DP_mult_207_n394), .ZN(DP_mult_207_n390) );
  NOR2_X1 DP_mult_207_U1873 ( .A1(DP_mult_207_n384), .A2(DP_mult_207_n364), 
        .ZN(DP_mult_207_n362) );
  INV_X1 DP_mult_207_U1872 ( .A(DP_mult_207_n396), .ZN(DP_mult_207_n394) );
  INV_X1 DP_mult_207_U1871 ( .A(DP_mult_207_n384), .ZN(DP_mult_207_n657) );
  NAND2_X1 DP_mult_207_U1870 ( .A1(DP_mult_207_n657), .A2(DP_mult_207_n387), 
        .ZN(DP_mult_207_n306) );
  INV_X1 DP_mult_207_U1869 ( .A(DP_mult_207_n400), .ZN(DP_mult_207_n398) );
  NAND2_X1 DP_mult_207_U1868 ( .A1(DP_mult_207_n2172), .A2(DP_mult_207_n396), 
        .ZN(DP_mult_207_n307) );
  NAND2_X1 DP_mult_207_U1867 ( .A1(DP_mult_207_n422), .A2(DP_mult_207_n2171), 
        .ZN(DP_mult_207_n411) );
  NAND2_X1 DP_mult_207_U1866 ( .A1(DP_mult_207_n821), .A2(DP_mult_207_n838), 
        .ZN(DP_mult_207_n503) );
  NOR2_X1 DP_mult_207_U1865 ( .A1(DP_mult_207_n435), .A2(DP_mult_207_n428), 
        .ZN(DP_mult_207_n426) );
  NAND2_X1 DP_mult_207_U1864 ( .A1(DP_mult_207_n661), .A2(DP_mult_207_n429), 
        .ZN(DP_mult_207_n310) );
  NAND2_X1 DP_mult_207_U1863 ( .A1(DP_mult_207_n789), .A2(DP_mult_207_n804), 
        .ZN(DP_mult_207_n481) );
  NOR2_X1 DP_mult_207_U1862 ( .A1(DP_mult_207_n896), .A2(DP_mult_207_n877), 
        .ZN(DP_mult_207_n531) );
  NAND2_X1 DP_mult_207_U1861 ( .A1(DP_mult_207_n2171), .A2(DP_mult_207_n418), 
        .ZN(DP_mult_207_n309) );
  OR2_X1 DP_mult_207_U1860 ( .A1(DP_mult_207_n1055), .A2(DP_mult_207_n1070), 
        .ZN(DP_mult_207_n2166) );
  NOR2_X1 DP_mult_207_U1859 ( .A1(DP_mult_207_n1071), .A2(DP_mult_207_n1084), 
        .ZN(DP_mult_207_n590) );
  INV_X1 DP_mult_207_U1858 ( .A(DP_mult_207_n409), .ZN(DP_mult_207_n407) );
  AOI21_X1 DP_mult_207_U1857 ( .B1(DP_mult_207_n2177), .B2(DP_mult_207_n416), 
        .A(DP_mult_207_n407), .ZN(DP_mult_207_n405) );
  NOR2_X1 DP_mult_207_U1856 ( .A1(DP_mult_207_n789), .A2(DP_mult_207_n804), 
        .ZN(DP_mult_207_n480) );
  INV_X1 DP_mult_207_U1855 ( .A(DP_mult_207_n461), .ZN(DP_mult_207_n459) );
  INV_X1 DP_mult_207_U1854 ( .A(DP_mult_207_n438), .ZN(DP_mult_207_n663) );
  INV_X1 DP_mult_207_U1853 ( .A(DP_mult_207_n436), .ZN(DP_mult_207_n434) );
  AOI21_X1 DP_mult_207_U1852 ( .B1(DP_mult_207_n662), .B2(DP_mult_207_n445), 
        .A(DP_mult_207_n434), .ZN(DP_mult_207_n432) );
  INV_X1 DP_mult_207_U1851 ( .A(DP_mult_207_n563), .ZN(DP_mult_207_n561) );
  INV_X1 DP_mult_207_U1850 ( .A(DP_mult_207_n564), .ZN(DP_mult_207_n562) );
  AOI21_X1 DP_mult_207_U1849 ( .B1(DP_mult_207_n565), .B2(DP_mult_207_n561), 
        .A(DP_mult_207_n562), .ZN(DP_mult_207_n560) );
  AOI21_X1 DP_mult_207_U1848 ( .B1(DP_mult_207_n565), .B2(DP_mult_207_n545), 
        .A(DP_mult_207_n546), .ZN(DP_mult_207_n544) );
  NOR2_X1 DP_mult_207_U1847 ( .A1(DP_mult_207_n402), .A2(DP_mult_207_n360), 
        .ZN(DP_mult_207_n356) );
  NAND2_X1 DP_mult_207_U1846 ( .A1(DP_mult_207_n662), .A2(DP_mult_207_n436), 
        .ZN(DP_mult_207_n311) );
  INV_X1 DP_mult_207_U1845 ( .A(DP_mult_207_n481), .ZN(DP_mult_207_n483) );
  NAND2_X1 DP_mult_207_U1844 ( .A1(DP_mult_207_n478), .A2(DP_mult_207_n2207), 
        .ZN(DP_mult_207_n476) );
  INV_X1 DP_mult_207_U1843 ( .A(DP_mult_207_n503), .ZN(DP_mult_207_n501) );
  NAND2_X1 DP_mult_207_U1842 ( .A1(DP_mult_207_n2207), .A2(DP_mult_207_n668), 
        .ZN(DP_mult_207_n498) );
  INV_X1 DP_mult_207_U1841 ( .A(DP_mult_207_n435), .ZN(DP_mult_207_n662) );
  NOR2_X1 DP_mult_207_U1840 ( .A1(DP_mult_207_n420), .A2(DP_mult_207_n402), 
        .ZN(DP_mult_207_n400) );
  OAI21_X1 DP_mult_207_U1839 ( .B1(DP_mult_207_n421), .B2(DP_mult_207_n402), 
        .A(DP_mult_207_n405), .ZN(DP_mult_207_n401) );
  INV_X1 DP_mult_207_U1838 ( .A(DP_mult_207_n401), .ZN(DP_mult_207_n399) );
  NAND2_X1 DP_mult_207_U1837 ( .A1(DP_mult_207_n663), .A2(DP_mult_207_n662), 
        .ZN(DP_mult_207_n431) );
  NAND2_X1 DP_mult_207_U1836 ( .A1(DP_mult_207_n465), .A2(DP_mult_207_n2207), 
        .ZN(DP_mult_207_n463) );
  AND2_X1 DP_mult_207_U1835 ( .A1(DP_mult_207_n511), .A2(DP_mult_207_n2088), 
        .ZN(DP_mult_207_n2207) );
  INV_X2 DP_mult_207_U1834 ( .A(DP_mult_207_n2268), .ZN(DP_mult_207_n2265) );
  INV_X2 DP_mult_207_U1833 ( .A(DP_mult_207_n2279), .ZN(DP_mult_207_n2276) );
  INV_X2 DP_mult_207_U1832 ( .A(DP_mult_207_n2289), .ZN(DP_mult_207_n2286) );
  INV_X2 DP_mult_207_U1831 ( .A(DP_mult_207_n2306), .ZN(DP_mult_207_n2303) );
  INV_X2 DP_mult_207_U1830 ( .A(DP_mult_207_n2302), .ZN(DP_mult_207_n2299) );
  INV_X2 DP_mult_207_U1829 ( .A(DP_mult_207_n2297), .ZN(DP_mult_207_n2294) );
  AOI21_X1 DP_mult_207_U1828 ( .B1(DP_mult_207_n526), .B2(DP_mult_207_n511), 
        .A(DP_mult_207_n512), .ZN(DP_mult_207_n2165) );
  OR2_X1 DP_mult_207_U1827 ( .A1(DP_mult_207_n805), .A2(DP_mult_207_n820), 
        .ZN(DP_mult_207_n2164) );
  INV_X1 DP_mult_207_U1826 ( .A(DP_mult_207_n492), .ZN(DP_mult_207_n2163) );
  NOR2_X1 DP_mult_207_U1825 ( .A1(DP_mult_207_n839), .A2(DP_mult_207_n856), 
        .ZN(DP_mult_207_n2162) );
  AND2_X2 DP_mult_207_U1824 ( .A1(DP_mult_207_n1812), .A2(DP_mult_207_n2248), 
        .ZN(DP_mult_207_n2188) );
  INV_X2 DP_mult_207_U1823 ( .A(DP_mult_207_n2278), .ZN(DP_mult_207_n2275) );
  OR2_X1 DP_mult_207_U1822 ( .A1(DP_mult_207_n896), .A2(DP_mult_207_n877), 
        .ZN(DP_mult_207_n2161) );
  CLKBUF_X1 DP_mult_207_U1821 ( .A(DP_mult_207_n526), .Z(DP_mult_207_n2160) );
  NAND3_X1 DP_mult_207_U1820 ( .A1(DP_mult_207_n2157), .A2(DP_mult_207_n2158), 
        .A3(DP_mult_207_n2159), .ZN(DP_mult_207_n972) );
  NAND2_X1 DP_mult_207_U1819 ( .A1(DP_mult_207_n996), .A2(DP_mult_207_n1217), 
        .ZN(DP_mult_207_n2159) );
  NAND2_X1 DP_mult_207_U1818 ( .A1(DP_mult_207_n994), .A2(DP_mult_207_n1217), 
        .ZN(DP_mult_207_n2158) );
  NAND2_X1 DP_mult_207_U1817 ( .A1(DP_mult_207_n994), .A2(DP_mult_207_n996), 
        .ZN(DP_mult_207_n2157) );
  XOR2_X1 DP_mult_207_U1816 ( .A(DP_mult_207_n2032), .B(DP_mult_207_n2156), 
        .Z(DP_mult_207_n973) );
  XOR2_X1 DP_mult_207_U1815 ( .A(DP_mult_207_n996), .B(DP_mult_207_n1217), .Z(
        DP_mult_207_n2156) );
  INV_X2 DP_mult_207_U1814 ( .A(DP_mult_207_n2296), .ZN(DP_mult_207_n2293) );
  INV_X2 DP_mult_207_U1813 ( .A(DP_mult_207_n2302), .ZN(DP_mult_207_n2298) );
  NOR2_X1 DP_mult_207_U1812 ( .A1(DP_mult_207_n1941), .A2(DP_mult_207_n940), 
        .ZN(DP_mult_207_n542) );
  NOR2_X1 DP_mult_207_U1811 ( .A1(DP_mult_207_n1941), .A2(DP_mult_207_n940), 
        .ZN(DP_mult_207_n2155) );
  NAND3_X1 DP_mult_207_U1810 ( .A1(DP_mult_207_n2152), .A2(DP_mult_207_n2153), 
        .A3(DP_mult_207_n2154), .ZN(DP_mult_207_n822) );
  NAND2_X1 DP_mult_207_U1809 ( .A1(DP_mult_207_n844), .A2(DP_mult_207_n827), 
        .ZN(DP_mult_207_n2154) );
  NAND2_X1 DP_mult_207_U1808 ( .A1(DP_mult_207_n842), .A2(DP_mult_207_n827), 
        .ZN(DP_mult_207_n2153) );
  NAND2_X1 DP_mult_207_U1807 ( .A1(DP_mult_207_n842), .A2(DP_mult_207_n844), 
        .ZN(DP_mult_207_n2152) );
  INV_X2 DP_mult_207_U1806 ( .A(DP_mult_207_n2102), .ZN(DP_mult_207_n2239) );
  INV_X2 DP_mult_207_U1805 ( .A(DP_mult_207_n2310), .ZN(DP_mult_207_n2307) );
  AND2_X2 DP_mult_207_U1804 ( .A1(DP_mult_207_n1815), .A2(DP_mult_207_n1990), 
        .ZN(DP_mult_207_n2190) );
  INV_X1 DP_mult_207_U1803 ( .A(DP_mult_207_n2190), .ZN(DP_mult_207_n2232) );
  INV_X1 DP_mult_207_U1802 ( .A(DP_mult_207_n2190), .ZN(DP_mult_207_n2150) );
  INV_X1 DP_mult_207_U1801 ( .A(DP_mult_207_n2190), .ZN(DP_mult_207_n2151) );
  CLKBUF_X1 DP_mult_207_U1800 ( .A(DP_mult_207_n520), .Z(DP_mult_207_n2149) );
  INV_X1 DP_mult_207_U1799 ( .A(DP_mult_207_n2043), .ZN(DP_mult_207_n2248) );
  AOI21_X1 DP_mult_207_U1798 ( .B1(DP_mult_207_n2000), .B2(DP_mult_207_n567), 
        .A(DP_mult_207_n2024), .ZN(DP_mult_207_n2148) );
  NAND3_X1 DP_mult_207_U1797 ( .A1(DP_mult_207_n2145), .A2(DP_mult_207_n2146), 
        .A3(DP_mult_207_n2147), .ZN(DP_mult_207_n1020) );
  NAND2_X1 DP_mult_207_U1796 ( .A1(DP_mult_207_n1025), .A2(DP_mult_207_n1040), 
        .ZN(DP_mult_207_n2147) );
  NAND2_X1 DP_mult_207_U1795 ( .A1(DP_mult_207_n1023), .A2(DP_mult_207_n1040), 
        .ZN(DP_mult_207_n2146) );
  NAND2_X1 DP_mult_207_U1794 ( .A1(DP_mult_207_n1023), .A2(DP_mult_207_n1025), 
        .ZN(DP_mult_207_n2145) );
  INV_X1 DP_mult_207_U1793 ( .A(DP_mult_207_n2187), .ZN(DP_mult_207_n2144) );
  INV_X2 DP_mult_207_U1792 ( .A(DP_mult_207_n2273), .ZN(DP_mult_207_n2270) );
  INV_X1 DP_mult_207_U1791 ( .A(DP_mult_207_n2273), .ZN(DP_mult_207_n2269) );
  NAND3_X1 DP_mult_207_U1790 ( .A1(DP_mult_207_n2141), .A2(DP_mult_207_n2142), 
        .A3(DP_mult_207_n2143), .ZN(DP_mult_207_n954) );
  NAND2_X1 DP_mult_207_U1789 ( .A1(DP_mult_207_n1304), .A2(DP_mult_207_n1414), 
        .ZN(DP_mult_207_n2143) );
  NAND2_X1 DP_mult_207_U1788 ( .A1(DP_mult_207_n1282), .A2(DP_mult_207_n1414), 
        .ZN(DP_mult_207_n2142) );
  NAND2_X1 DP_mult_207_U1787 ( .A1(DP_mult_207_n1282), .A2(DP_mult_207_n1304), 
        .ZN(DP_mult_207_n2141) );
  OR2_X1 DP_mult_207_U1786 ( .A1(DP_mult_207_n1941), .A2(DP_mult_207_n940), 
        .ZN(DP_mult_207_n2139) );
  NAND3_X1 DP_mult_207_U1785 ( .A1(DP_mult_207_n2136), .A2(DP_mult_207_n2137), 
        .A3(DP_mult_207_n2138), .ZN(DP_mult_207_n928) );
  NAND2_X1 DP_mult_207_U1784 ( .A1(DP_mult_207_n956), .A2(DP_mult_207_n958), 
        .ZN(DP_mult_207_n2138) );
  NAND2_X1 DP_mult_207_U1783 ( .A1(DP_mult_207_n954), .A2(DP_mult_207_n958), 
        .ZN(DP_mult_207_n2137) );
  NAND2_X1 DP_mult_207_U1782 ( .A1(DP_mult_207_n2019), .A2(DP_mult_207_n2001), 
        .ZN(DP_mult_207_n2136) );
  XOR2_X1 DP_mult_207_U1781 ( .A(DP_mult_207_n2135), .B(DP_mult_207_n958), .Z(
        DP_mult_207_n929) );
  XOR2_X1 DP_mult_207_U1780 ( .A(DP_mult_207_n2002), .B(DP_mult_207_n2020), 
        .Z(DP_mult_207_n2135) );
  NAND2_X1 DP_mult_207_U1779 ( .A1(DP_mult_207_n1348), .A2(DP_mult_207_n1182), 
        .ZN(DP_mult_207_n2134) );
  NAND2_X1 DP_mult_207_U1778 ( .A1(DP_mult_207_n1260), .A2(DP_mult_207_n1182), 
        .ZN(DP_mult_207_n2133) );
  NAND2_X1 DP_mult_207_U1777 ( .A1(DP_mult_207_n1260), .A2(DP_mult_207_n1348), 
        .ZN(DP_mult_207_n2132) );
  XOR2_X1 DP_mult_207_U1776 ( .A(DP_mult_207_n2131), .B(DP_mult_207_n1182), 
        .Z(DP_mult_207_n959) );
  XOR2_X1 DP_mult_207_U1775 ( .A(DP_mult_207_n1260), .B(DP_mult_207_n1348), 
        .Z(DP_mult_207_n2131) );
  AND2_X2 DP_mult_207_U1774 ( .A1(DP_mult_207_n1814), .A2(DP_mult_207_n2047), 
        .ZN(DP_mult_207_n2191) );
  XNOR2_X1 DP_mult_207_U1773 ( .A(DP_mult_207_n1040), .B(DP_mult_207_n1025), 
        .ZN(DP_mult_207_n2129) );
  XNOR2_X1 DP_mult_207_U1772 ( .A(DP_mult_207_n2129), .B(DP_mult_207_n1023), 
        .ZN(DP_mult_207_n1021) );
  INV_X2 DP_mult_207_U1771 ( .A(DP_mult_207_n2186), .ZN(DP_mult_207_n2140) );
  INV_X1 DP_mult_207_U1770 ( .A(DP_mult_207_n2128), .ZN(DP_mult_207_n2186) );
  OR2_X1 DP_mult_207_U1769 ( .A1(DP_mult_207_n941), .A2(DP_mult_207_n962), 
        .ZN(DP_mult_207_n2127) );
  NOR2_X1 DP_mult_207_U1768 ( .A1(DP_mult_207_n547), .A2(DP_mult_207_n542), 
        .ZN(DP_mult_207_n2126) );
  NAND3_X1 DP_mult_207_U1767 ( .A1(DP_mult_207_n2123), .A2(DP_mult_207_n2124), 
        .A3(DP_mult_207_n2125), .ZN(DP_mult_207_n940) );
  NAND2_X1 DP_mult_207_U1766 ( .A1(DP_mult_207_n945), .A2(DP_mult_207_n943), 
        .ZN(DP_mult_207_n2125) );
  NAND2_X1 DP_mult_207_U1765 ( .A1(DP_mult_207_n964), .A2(DP_mult_207_n943), 
        .ZN(DP_mult_207_n2124) );
  NAND2_X1 DP_mult_207_U1764 ( .A1(DP_mult_207_n964), .A2(DP_mult_207_n945), 
        .ZN(DP_mult_207_n2123) );
  NAND3_X1 DP_mult_207_U1763 ( .A1(DP_mult_207_n2120), .A2(DP_mult_207_n2121), 
        .A3(DP_mult_207_n2122), .ZN(DP_mult_207_n942) );
  NAND2_X1 DP_mult_207_U1762 ( .A1(DP_mult_207_n949), .A2(DP_mult_207_n966), 
        .ZN(DP_mult_207_n2122) );
  NAND2_X1 DP_mult_207_U1761 ( .A1(DP_mult_207_n947), .A2(DP_mult_207_n966), 
        .ZN(DP_mult_207_n2121) );
  NAND2_X1 DP_mult_207_U1760 ( .A1(DP_mult_207_n947), .A2(DP_mult_207_n949), 
        .ZN(DP_mult_207_n2120) );
  XOR2_X1 DP_mult_207_U1759 ( .A(DP_mult_207_n2119), .B(DP_mult_207_n966), .Z(
        DP_mult_207_n943) );
  XOR2_X1 DP_mult_207_U1758 ( .A(DP_mult_207_n947), .B(DP_mult_207_n949), .Z(
        DP_mult_207_n2119) );
  NAND3_X1 DP_mult_207_U1757 ( .A1(DP_mult_207_n2116), .A2(DP_mult_207_n2117), 
        .A3(DP_mult_207_n2118), .ZN(DP_mult_207_n918) );
  NAND2_X1 DP_mult_207_U1756 ( .A1(DP_mult_207_n2033), .A2(DP_mult_207_n923), 
        .ZN(DP_mult_207_n2118) );
  NAND2_X1 DP_mult_207_U1755 ( .A1(DP_mult_207_n921), .A2(DP_mult_207_n923), 
        .ZN(DP_mult_207_n2117) );
  NAND2_X1 DP_mult_207_U1754 ( .A1(DP_mult_207_n921), .A2(DP_mult_207_n2033), 
        .ZN(DP_mult_207_n2116) );
  INV_X1 DP_mult_207_U1753 ( .A(DP_mult_207_n491), .ZN(DP_mult_207_n2115) );
  INV_X1 DP_mult_207_U1752 ( .A(DP_mult_207_n2191), .ZN(DP_mult_207_n2114) );
  AND2_X2 DP_mult_207_U1751 ( .A1(DP_mult_207_n1813), .A2(DP_mult_207_n2251), 
        .ZN(DP_mult_207_n2193) );
  NAND3_X1 DP_mult_207_U1750 ( .A1(DP_mult_207_n2111), .A2(DP_mult_207_n2112), 
        .A3(DP_mult_207_n2113), .ZN(DP_mult_207_n882) );
  NAND2_X1 DP_mult_207_U1749 ( .A1(DP_mult_207_n889), .A2(DP_mult_207_n893), 
        .ZN(DP_mult_207_n2113) );
  NAND2_X1 DP_mult_207_U1748 ( .A1(DP_mult_207_n906), .A2(DP_mult_207_n893), 
        .ZN(DP_mult_207_n2112) );
  NAND2_X1 DP_mult_207_U1747 ( .A1(DP_mult_207_n906), .A2(DP_mult_207_n1929), 
        .ZN(DP_mult_207_n2111) );
  XOR2_X1 DP_mult_207_U1746 ( .A(DP_mult_207_n2110), .B(DP_mult_207_n906), .Z(
        DP_mult_207_n883) );
  XOR2_X1 DP_mult_207_U1745 ( .A(DP_mult_207_n889), .B(DP_mult_207_n893), .Z(
        DP_mult_207_n2110) );
  INV_X1 DP_mult_207_U1744 ( .A(DP_coeffs_ff_int[24]), .ZN(DP_mult_207_n2319)
         );
  NAND3_X1 DP_mult_207_U1743 ( .A1(DP_mult_207_n2107), .A2(DP_mult_207_n2108), 
        .A3(DP_mult_207_n2109), .ZN(DP_mult_207_n830) );
  NAND2_X1 DP_mult_207_U1742 ( .A1(DP_mult_207_n1320), .A2(DP_mult_207_n1254), 
        .ZN(DP_mult_207_n2109) );
  NAND2_X1 DP_mult_207_U1741 ( .A1(DP_mult_207_n1298), .A2(DP_mult_207_n1254), 
        .ZN(DP_mult_207_n2108) );
  NAND2_X1 DP_mult_207_U1740 ( .A1(DP_mult_207_n1298), .A2(DP_mult_207_n1320), 
        .ZN(DP_mult_207_n2107) );
  XOR2_X1 DP_mult_207_U1739 ( .A(DP_mult_207_n1994), .B(DP_mult_207_n2106), 
        .Z(DP_mult_207_n831) );
  XOR2_X1 DP_mult_207_U1738 ( .A(DP_mult_207_n1320), .B(DP_mult_207_n1254), 
        .Z(DP_mult_207_n2106) );
  INV_X2 DP_mult_207_U1737 ( .A(DP_mult_207_n2283), .ZN(DP_mult_207_n2280) );
  AND2_X1 DP_mult_207_U1736 ( .A1(DP_mult_207_n2214), .A2(DP_mult_207_n2213), 
        .ZN(DP_mult_207_n301) );
  INV_X2 DP_mult_207_U1735 ( .A(DP_mult_207_n2195), .ZN(DP_mult_207_n2105) );
  AND2_X1 DP_mult_207_U1734 ( .A1(DP_mult_207_n2214), .A2(DP_mult_207_n2213), 
        .ZN(DP_mult_207_n2103) );
  AND2_X1 DP_mult_207_U1733 ( .A1(DP_mult_207_n2214), .A2(DP_mult_207_n2213), 
        .ZN(DP_mult_207_n2104) );
  AND2_X1 DP_mult_207_U1732 ( .A1(DP_mult_207_n2213), .A2(DP_mult_207_n2214), 
        .ZN(DP_mult_207_n2212) );
  XNOR2_X1 DP_mult_207_U1731 ( .A(DP_mult_207_n942), .B(DP_mult_207_n923), 
        .ZN(DP_mult_207_n2101) );
  NAND3_X1 DP_mult_207_U1730 ( .A1(DP_mult_207_n2098), .A2(DP_mult_207_n2099), 
        .A3(DP_mult_207_n2100), .ZN(DP_mult_207_n1038) );
  NAND2_X1 DP_mult_207_U1729 ( .A1(DP_mult_207_n1056), .A2(DP_mult_207_n1043), 
        .ZN(DP_mult_207_n2100) );
  NAND2_X1 DP_mult_207_U1728 ( .A1(DP_mult_207_n1041), .A2(DP_mult_207_n1043), 
        .ZN(DP_mult_207_n2099) );
  NAND2_X1 DP_mult_207_U1727 ( .A1(DP_mult_207_n1041), .A2(DP_mult_207_n1056), 
        .ZN(DP_mult_207_n2098) );
  AND2_X2 DP_mult_207_U1726 ( .A1(DP_mult_207_n1811), .A2(DP_mult_207_n2245), 
        .ZN(DP_mult_207_n2192) );
  NOR2_X1 DP_mult_207_U1725 ( .A1(DP_mult_207_n963), .A2(DP_mult_207_n982), 
        .ZN(DP_mult_207_n558) );
  NOR2_X1 DP_mult_207_U1724 ( .A1(DP_mult_207_n963), .A2(DP_mult_207_n982), 
        .ZN(DP_mult_207_n2097) );
  NAND2_X1 DP_mult_207_U1723 ( .A1(DP_mult_207_n1806), .A2(DP_mult_207_n2185), 
        .ZN(DP_mult_207_n2184) );
  BUF_X2 DP_mult_207_U1722 ( .A(DP_mult_207_n2184), .Z(DP_mult_207_n2095) );
  CLKBUF_X3 DP_mult_207_U1721 ( .A(DP_mult_207_n2184), .Z(DP_mult_207_n2096)
         );
  BUF_X1 DP_mult_207_U1720 ( .A(DP_mult_207_n2184), .Z(DP_mult_207_n2094) );
  OAI22_X1 DP_mult_207_U1719 ( .A1(DP_mult_207_n2094), .A2(DP_mult_207_n1504), 
        .B1(DP_mult_207_n2237), .B2(DP_mult_207_n1503), .ZN(DP_mult_207_n2093)
         );
  INV_X1 DP_mult_207_U1718 ( .A(DP_mult_207_n2043), .ZN(DP_mult_207_n2250) );
  INV_X2 DP_mult_207_U1717 ( .A(DP_mult_207_n2289), .ZN(DP_mult_207_n2092) );
  OR2_X1 DP_mult_207_U1716 ( .A1(DP_mult_207_n856), .A2(DP_mult_207_n1932), 
        .ZN(DP_mult_207_n2091) );
  NOR2_X1 DP_mult_207_U1715 ( .A1(DP_mult_207_n877), .A2(DP_mult_207_n896), 
        .ZN(DP_mult_207_n2090) );
  OAI22_X1 DP_mult_207_U1714 ( .A1(DP_mult_207_n2234), .A2(DP_mult_207_n1733), 
        .B1(DP_mult_207_n1732), .B2(DP_mult_207_n2259), .ZN(DP_mult_207_n2089)
         );
  BUF_X2 DP_mult_207_U1713 ( .A(DP_mult_207_n2223), .Z(DP_mult_207_n2200) );
  NOR2_X1 DP_mult_207_U1712 ( .A1(DP_mult_207_n531), .A2(DP_mult_207_n534), 
        .ZN(DP_mult_207_n2088) );
  INV_X1 DP_mult_207_U1711 ( .A(DP_mult_207_n1987), .ZN(DP_mult_207_n2245) );
  INV_X2 DP_mult_207_U1710 ( .A(DP_mult_207_n2195), .ZN(DP_mult_207_n2233) );
  INV_X1 DP_mult_207_U1709 ( .A(DP_mult_207_n2082), .ZN(DP_mult_207_n2255) );
  INV_X1 DP_mult_207_U1708 ( .A(DP_mult_207_n2249), .ZN(DP_mult_207_n2087) );
  XNOR2_X1 DP_mult_207_U1707 ( .A(DP_mult_207_n964), .B(DP_mult_207_n945), 
        .ZN(DP_mult_207_n2086) );
  XNOR2_X1 DP_mult_207_U1706 ( .A(DP_mult_207_n2086), .B(DP_mult_207_n943), 
        .ZN(DP_mult_207_n941) );
  NOR2_X1 DP_mult_207_U1705 ( .A1(DP_mult_207_n805), .A2(DP_mult_207_n820), 
        .ZN(DP_mult_207_n2085) );
  INV_X1 DP_mult_207_U1704 ( .A(DP_mult_207_n1951), .ZN(DP_mult_207_n2249) );
  INV_X1 DP_mult_207_U1703 ( .A(DP_mult_207_n2066), .ZN(DP_mult_207_n2258) );
  BUF_X2 DP_mult_207_U1702 ( .A(DP_mult_207_n2114), .Z(DP_mult_207_n2196) );
  INV_X1 DP_mult_207_U1701 ( .A(DP_mult_207_n2188), .ZN(DP_mult_207_n2226) );
  INV_X1 DP_mult_207_U1700 ( .A(DP_mult_207_n2188), .ZN(DP_mult_207_n2080) );
  INV_X2 DP_mult_207_U1699 ( .A(DP_mult_207_n2130), .ZN(DP_mult_207_n2241) );
  CLKBUF_X1 DP_mult_207_U1698 ( .A(DP_mult_207_n2256), .Z(DP_mult_207_n2078)
         );
  XNOR2_X1 DP_mult_207_U1697 ( .A(DP_coeffs_ff_int[29]), .B(
        DP_coeffs_ff_int[30]), .ZN(DP_mult_207_n2128) );
  INV_X2 DP_mult_207_U1696 ( .A(DP_mult_207_n2076), .ZN(DP_mult_207_n2077) );
  INV_X1 DP_mult_207_U1695 ( .A(DP_mult_207_n2128), .ZN(DP_mult_207_n2076) );
  INV_X1 DP_mult_207_U1694 ( .A(DP_mult_207_n555), .ZN(DP_mult_207_n2075) );
  NAND2_X1 DP_mult_207_U1693 ( .A1(DP_mult_207_n2073), .A2(DP_mult_207_n2074), 
        .ZN(DP_mult_207_n1370) );
  OR2_X1 DP_mult_207_U1692 ( .A1(DP_mult_207_n1665), .A2(DP_mult_207_n2252), 
        .ZN(DP_mult_207_n2074) );
  OR2_X1 DP_mult_207_U1691 ( .A1(DP_mult_207_n2227), .A2(DP_mult_207_n1666), 
        .ZN(DP_mult_207_n2073) );
  NAND3_X1 DP_mult_207_U1690 ( .A1(DP_mult_207_n2070), .A2(DP_mult_207_n2071), 
        .A3(DP_mult_207_n2072), .ZN(DP_mult_207_n956) );
  NAND2_X1 DP_mult_207_U1689 ( .A1(DP_mult_207_n1459), .A2(DP_mult_207_n1436), 
        .ZN(DP_mult_207_n2072) );
  NAND2_X1 DP_mult_207_U1688 ( .A1(DP_mult_207_n1370), .A2(DP_mult_207_n1436), 
        .ZN(DP_mult_207_n2071) );
  NAND2_X1 DP_mult_207_U1687 ( .A1(DP_mult_207_n1370), .A2(DP_mult_207_n1459), 
        .ZN(DP_mult_207_n2070) );
  XOR2_X1 DP_mult_207_U1686 ( .A(DP_mult_207_n1370), .B(DP_mult_207_n2069), 
        .Z(DP_mult_207_n957) );
  XOR2_X1 DP_mult_207_U1685 ( .A(DP_mult_207_n1436), .B(DP_mult_207_n1459), 
        .Z(DP_mult_207_n2069) );
  INV_X1 DP_mult_207_U1684 ( .A(DP_mult_207_n2209), .ZN(DP_mult_207_n2215) );
  INV_X1 DP_mult_207_U1683 ( .A(DP_mult_207_n2079), .ZN(DP_mult_207_n2130) );
  XNOR2_X1 DP_mult_207_U1682 ( .A(DP_mult_207_n1414), .B(DP_mult_207_n1304), 
        .ZN(DP_mult_207_n2068) );
  XNOR2_X1 DP_mult_207_U1681 ( .A(DP_mult_207_n2068), .B(DP_mult_207_n1282), 
        .ZN(DP_mult_207_n955) );
  INV_X1 DP_mult_207_U1680 ( .A(DP_mult_207_n2216), .ZN(DP_mult_207_n2067) );
  INV_X1 DP_mult_207_U1679 ( .A(DP_mult_207_n2193), .ZN(DP_mult_207_n2227) );
  INV_X1 DP_mult_207_U1678 ( .A(DP_mult_207_n2188), .ZN(DP_mult_207_n2081) );
  NAND3_X1 DP_mult_207_U1677 ( .A1(DP_mult_207_n2063), .A2(DP_mult_207_n2064), 
        .A3(DP_mult_207_n2065), .ZN(DP_mult_207_n1126) );
  NAND2_X1 DP_mult_207_U1676 ( .A1(DP_mult_207_n1337), .A2(DP_mult_207_n1138), 
        .ZN(DP_mult_207_n2065) );
  NAND2_X1 DP_mult_207_U1675 ( .A1(DP_mult_207_n1140), .A2(DP_mult_207_n1138), 
        .ZN(DP_mult_207_n2064) );
  NAND2_X1 DP_mult_207_U1674 ( .A1(DP_mult_207_n1140), .A2(DP_mult_207_n1337), 
        .ZN(DP_mult_207_n2063) );
  XOR2_X1 DP_mult_207_U1673 ( .A(DP_mult_207_n2062), .B(DP_mult_207_n1138), 
        .Z(DP_mult_207_n1127) );
  XOR2_X1 DP_mult_207_U1672 ( .A(DP_mult_207_n1140), .B(DP_mult_207_n1337), 
        .Z(DP_mult_207_n2062) );
  NAND3_X1 DP_mult_207_U1671 ( .A1(DP_mult_207_n2059), .A2(DP_mult_207_n2060), 
        .A3(DP_mult_207_n2061), .ZN(DP_mult_207_n1138) );
  NAND2_X1 DP_mult_207_U1670 ( .A1(DP_mult_207_n1188), .A2(DP_mult_207_n1426), 
        .ZN(DP_mult_207_n2061) );
  NAND2_X1 DP_mult_207_U1669 ( .A1(DP_mult_207_n1471), .A2(DP_mult_207_n1426), 
        .ZN(DP_mult_207_n2060) );
  NAND2_X1 DP_mult_207_U1668 ( .A1(DP_mult_207_n1471), .A2(DP_mult_207_n1188), 
        .ZN(DP_mult_207_n2059) );
  XOR2_X1 DP_mult_207_U1667 ( .A(DP_mult_207_n2058), .B(DP_mult_207_n1426), 
        .Z(DP_mult_207_n1139) );
  XOR2_X1 DP_mult_207_U1666 ( .A(DP_mult_207_n1471), .B(DP_mult_207_n1188), 
        .Z(DP_mult_207_n2058) );
  NAND3_X1 DP_mult_207_U1665 ( .A1(DP_mult_207_n2054), .A2(DP_mult_207_n2055), 
        .A3(DP_mult_207_n2056), .ZN(DP_mult_207_n920) );
  NAND2_X1 DP_mult_207_U1664 ( .A1(DP_mult_207_n925), .A2(DP_mult_207_n927), 
        .ZN(DP_mult_207_n2056) );
  NAND2_X1 DP_mult_207_U1663 ( .A1(DP_mult_207_n944), .A2(DP_mult_207_n927), 
        .ZN(DP_mult_207_n2055) );
  NAND2_X1 DP_mult_207_U1662 ( .A1(DP_mult_207_n944), .A2(DP_mult_207_n925), 
        .ZN(DP_mult_207_n2054) );
  INV_X1 DP_mult_207_U1661 ( .A(DP_mult_207_n2209), .ZN(DP_mult_207_n2053) );
  NOR2_X1 DP_mult_207_U1660 ( .A1(DP_mult_207_n2102), .A2(DP_mult_207_n2052), 
        .ZN(DP_mult_207_n2194) );
  BUF_X2 DP_mult_207_U1659 ( .A(DP_mult_207_n2217), .Z(DP_mult_207_n2202) );
  XNOR2_X1 DP_mult_207_U1658 ( .A(DP_coeffs_ff_int[41]), .B(DP_mult_207_n2283), 
        .ZN(DP_mult_207_n1814) );
  NAND3_X1 DP_mult_207_U1657 ( .A1(DP_mult_207_n2049), .A2(DP_mult_207_n2050), 
        .A3(DP_mult_207_n2051), .ZN(DP_mult_207_n790) );
  NAND2_X1 DP_mult_207_U1656 ( .A1(DP_mult_207_n795), .A2(DP_mult_207_n810), 
        .ZN(DP_mult_207_n2051) );
  NAND2_X1 DP_mult_207_U1655 ( .A1(DP_mult_207_n808), .A2(DP_mult_207_n810), 
        .ZN(DP_mult_207_n2050) );
  NAND2_X1 DP_mult_207_U1654 ( .A1(DP_mult_207_n808), .A2(DP_mult_207_n795), 
        .ZN(DP_mult_207_n2049) );
  XOR2_X1 DP_mult_207_U1653 ( .A(DP_mult_207_n808), .B(DP_mult_207_n2048), .Z(
        DP_mult_207_n791) );
  XOR2_X1 DP_mult_207_U1652 ( .A(DP_mult_207_n795), .B(DP_mult_207_n810), .Z(
        DP_mult_207_n2048) );
  INV_X1 DP_mult_207_U1651 ( .A(DP_mult_207_n2316), .ZN(DP_mult_207_n2311) );
  XNOR2_X1 DP_mult_207_U1650 ( .A(DP_coeffs_ff_int[25]), .B(DP_mult_207_n2316), 
        .ZN(DP_mult_207_n2210) );
  INV_X1 DP_mult_207_U1649 ( .A(DP_mult_207_n2193), .ZN(DP_mult_207_n2228) );
  INV_X1 DP_mult_207_U1648 ( .A(DP_mult_207_n2193), .ZN(DP_mult_207_n2044) );
  INV_X1 DP_mult_207_U1647 ( .A(DP_mult_207_n2193), .ZN(DP_mult_207_n2045) );
  INV_X1 DP_mult_207_U1646 ( .A(DP_mult_207_n2188), .ZN(DP_mult_207_n2225) );
  NOR2_X1 DP_mult_207_U1645 ( .A1(DP_mult_207_n495), .A2(DP_mult_207_n502), 
        .ZN(DP_mult_207_n2042) );
  NAND3_X1 DP_mult_207_U1644 ( .A1(DP_mult_207_n2039), .A2(DP_mult_207_n2040), 
        .A3(DP_mult_207_n2041), .ZN(DP_mult_207_n842) );
  NAND2_X1 DP_mult_207_U1643 ( .A1(DP_mult_207_n849), .A2(DP_mult_207_n864), 
        .ZN(DP_mult_207_n2041) );
  NAND2_X1 DP_mult_207_U1642 ( .A1(DP_mult_207_n862), .A2(DP_mult_207_n864), 
        .ZN(DP_mult_207_n2040) );
  NAND2_X1 DP_mult_207_U1641 ( .A1(DP_mult_207_n862), .A2(DP_mult_207_n849), 
        .ZN(DP_mult_207_n2039) );
  XOR2_X1 DP_mult_207_U1640 ( .A(DP_mult_207_n862), .B(DP_mult_207_n2038), .Z(
        DP_mult_207_n843) );
  XOR2_X1 DP_mult_207_U1639 ( .A(DP_mult_207_n849), .B(DP_mult_207_n864), .Z(
        DP_mult_207_n2038) );
  BUF_X1 DP_mult_207_U1638 ( .A(DP_mult_207_n1372), .Z(DP_mult_207_n2037) );
  NAND3_X1 DP_mult_207_U1637 ( .A1(DP_mult_207_n2034), .A2(DP_mult_207_n2035), 
        .A3(DP_mult_207_n2036), .ZN(DP_mult_207_n996) );
  NAND2_X1 DP_mult_207_U1636 ( .A1(DP_mult_207_n1284), .A2(DP_mult_207_n1438), 
        .ZN(DP_mult_207_n2036) );
  NAND2_X1 DP_mult_207_U1635 ( .A1(DP_mult_207_n1372), .A2(DP_mult_207_n1438), 
        .ZN(DP_mult_207_n2035) );
  NAND2_X1 DP_mult_207_U1634 ( .A1(DP_mult_207_n1372), .A2(DP_mult_207_n1284), 
        .ZN(DP_mult_207_n2034) );
  INV_X1 DP_mult_207_U1633 ( .A(DP_mult_207_n2288), .ZN(DP_mult_207_n2285) );
  XNOR2_X1 DP_mult_207_U1632 ( .A(DP_coeffs_ff_int[39]), .B(DP_mult_207_n2289), 
        .ZN(DP_mult_207_n1813) );
  NAND3_X1 DP_mult_207_U1631 ( .A1(DP_mult_207_n2120), .A2(DP_mult_207_n2121), 
        .A3(DP_mult_207_n2122), .ZN(DP_mult_207_n2033) );
  CLKBUF_X1 DP_mult_207_U1630 ( .A(DP_mult_207_n994), .Z(DP_mult_207_n2032) );
  NAND3_X1 DP_mult_207_U1629 ( .A1(DP_mult_207_n2029), .A2(DP_mult_207_n2030), 
        .A3(DP_mult_207_n2031), .ZN(DP_mult_207_n846) );
  NAND2_X1 DP_mult_207_U1628 ( .A1(DP_mult_207_n870), .A2(DP_mult_207_n868), 
        .ZN(DP_mult_207_n2031) );
  NAND2_X1 DP_mult_207_U1627 ( .A1(DP_mult_207_n851), .A2(DP_mult_207_n868), 
        .ZN(DP_mult_207_n2030) );
  NAND2_X1 DP_mult_207_U1626 ( .A1(DP_mult_207_n851), .A2(DP_mult_207_n870), 
        .ZN(DP_mult_207_n2029) );
  XOR2_X1 DP_mult_207_U1625 ( .A(DP_mult_207_n851), .B(DP_mult_207_n2028), .Z(
        DP_mult_207_n847) );
  XOR2_X1 DP_mult_207_U1624 ( .A(DP_mult_207_n870), .B(DP_mult_207_n868), .Z(
        DP_mult_207_n2028) );
  NAND3_X1 DP_mult_207_U1623 ( .A1(DP_mult_207_n2025), .A2(DP_mult_207_n2026), 
        .A3(DP_mult_207_n2027), .ZN(DP_mult_207_n908) );
  NAND2_X1 DP_mult_207_U1622 ( .A1(DP_mult_207_n1390), .A2(DP_mult_207_n1368), 
        .ZN(DP_mult_207_n2027) );
  NAND2_X1 DP_mult_207_U1621 ( .A1(DP_mult_207_n938), .A2(DP_mult_207_n1390), 
        .ZN(DP_mult_207_n2026) );
  NAND2_X1 DP_mult_207_U1620 ( .A1(DP_mult_207_n938), .A2(DP_mult_207_n1368), 
        .ZN(DP_mult_207_n2025) );
  INV_X2 DP_mult_207_U1619 ( .A(DP_mult_207_n2244), .ZN(DP_mult_207_n2242) );
  INV_X1 DP_mult_207_U1618 ( .A(DP_mult_207_n2189), .ZN(DP_mult_207_n2222) );
  INV_X1 DP_mult_207_U1617 ( .A(DP_mult_207_n2189), .ZN(DP_mult_207_n2022) );
  INV_X1 DP_mult_207_U1616 ( .A(DP_mult_207_n2189), .ZN(DP_mult_207_n2023) );
  INV_X1 DP_mult_207_U1615 ( .A(DP_mult_207_n2319), .ZN(DP_mult_207_n2318) );
  XNOR2_X1 DP_mult_207_U1614 ( .A(DP_coeffs_ff_int[25]), .B(DP_mult_207_n2319), 
        .ZN(DP_mult_207_n1806) );
  CLKBUF_X1 DP_mult_207_U1613 ( .A(DP_mult_207_n2256), .Z(DP_mult_207_n2021)
         );
  AOI21_X2 DP_mult_207_U1612 ( .B1(DP_mult_207_n426), .B2(DP_mult_207_n445), 
        .A(DP_mult_207_n427), .ZN(DP_mult_207_n421) );
  NAND3_X1 DP_mult_207_U1611 ( .A1(DP_mult_207_n2141), .A2(DP_mult_207_n2142), 
        .A3(DP_mult_207_n2143), .ZN(DP_mult_207_n2019) );
  NAND3_X1 DP_mult_207_U1610 ( .A1(DP_mult_207_n2141), .A2(DP_mult_207_n2142), 
        .A3(DP_mult_207_n2143), .ZN(DP_mult_207_n2020) );
  XNOR2_X1 DP_mult_207_U1609 ( .A(DP_mult_207_n925), .B(DP_mult_207_n927), 
        .ZN(DP_mult_207_n2018) );
  XNOR2_X1 DP_mult_207_U1608 ( .A(DP_mult_207_n944), .B(DP_mult_207_n2018), 
        .ZN(DP_mult_207_n921) );
  INV_X1 DP_mult_207_U1607 ( .A(DP_mult_207_n2188), .ZN(DP_mult_207_n2017) );
  INV_X1 DP_mult_207_U1606 ( .A(DP_mult_207_n2291), .ZN(DP_mult_207_n2015) );
  INV_X1 DP_mult_207_U1605 ( .A(DP_mult_207_n2291), .ZN(DP_mult_207_n2016) );
  INV_X1 DP_mult_207_U1604 ( .A(DP_pipe01[0]), .ZN(DP_mult_207_n2013) );
  INV_X1 DP_mult_207_U1603 ( .A(DP_pipe01[0]), .ZN(DP_mult_207_n2014) );
  INV_X1 DP_mult_207_U1602 ( .A(DP_pipe01[0]), .ZN(DP_mult_207_n2012) );
  INV_X1 DP_mult_207_U1601 ( .A(DP_mult_207_n1811), .ZN(DP_mult_207_n2011) );
  OR2_X1 DP_mult_207_U1600 ( .A1(DP_mult_207_n2011), .A2(DP_mult_207_n1988), 
        .ZN(DP_mult_207_n2199) );
  BUF_X4 DP_mult_207_U1599 ( .A(DP_mult_207_n251), .Z(DP_mult_207_n2261) );
  INV_X2 DP_mult_207_U1598 ( .A(DP_mult_207_n2010), .ZN(DP_mult_207_n2236) );
  AND2_X1 DP_mult_207_U1597 ( .A1(DP_mult_207_n2261), .A2(DP_coeffs_ff_int[46]), .ZN(DP_mult_207_n2010) );
  INV_X1 DP_mult_207_U1596 ( .A(DP_mult_207_n2189), .ZN(DP_mult_207_n2221) );
  XNOR2_X1 DP_mult_207_U1595 ( .A(DP_mult_207_n844), .B(DP_mult_207_n827), 
        .ZN(DP_mult_207_n2009) );
  XNOR2_X1 DP_mult_207_U1594 ( .A(DP_mult_207_n842), .B(DP_mult_207_n2009), 
        .ZN(DP_mult_207_n823) );
  XNOR2_X1 DP_mult_207_U1593 ( .A(DP_coeffs_ff_int[31]), .B(
        DP_coeffs_ff_int[32]), .ZN(DP_mult_207_n2079) );
  INV_X2 DP_mult_207_U1592 ( .A(DP_mult_207_n2007), .ZN(DP_mult_207_n2008) );
  INV_X1 DP_mult_207_U1591 ( .A(DP_mult_207_n2079), .ZN(DP_mult_207_n2007) );
  INV_X1 DP_mult_207_U1590 ( .A(DP_mult_207_n2244), .ZN(DP_mult_207_n2243) );
  XNOR2_X1 DP_mult_207_U1589 ( .A(DP_mult_207_n1056), .B(DP_mult_207_n1043), 
        .ZN(DP_mult_207_n2006) );
  XNOR2_X1 DP_mult_207_U1588 ( .A(DP_mult_207_n1041), .B(DP_mult_207_n2006), 
        .ZN(DP_mult_207_n1039) );
  BUF_X2 DP_mult_207_U1587 ( .A(DP_mult_207_n2217), .Z(DP_mult_207_n2201) );
  INV_X2 DP_mult_207_U1586 ( .A(DP_mult_207_n2066), .ZN(DP_mult_207_n2257) );
  INV_X1 DP_mult_207_U1585 ( .A(DP_mult_207_n2247), .ZN(DP_mult_207_n2005) );
  XNOR2_X1 DP_mult_207_U1584 ( .A(DP_mult_207_n1368), .B(DP_mult_207_n1390), 
        .ZN(DP_mult_207_n2004) );
  XNOR2_X1 DP_mult_207_U1583 ( .A(DP_mult_207_n2004), .B(DP_mult_207_n938), 
        .ZN(DP_mult_207_n909) );
  INV_X1 DP_mult_207_U1582 ( .A(DP_mult_207_n1988), .ZN(DP_mult_207_n2247) );
  INV_X2 DP_mult_207_U1581 ( .A(DP_mult_207_n1971), .ZN(DP_mult_207_n2235) );
  XOR2_X1 DP_mult_207_U1580 ( .A(DP_coeffs_ff_int[38]), .B(
        DP_coeffs_ff_int[37]), .Z(DP_mult_207_n2043) );
  INV_X1 DP_mult_207_U1579 ( .A(DP_mult_207_n2189), .ZN(DP_mult_207_n2003) );
  AND2_X2 DP_mult_207_U1578 ( .A1(DP_mult_207_n1809), .A2(DP_mult_207_n2079), 
        .ZN(DP_mult_207_n2187) );
  INV_X2 DP_mult_207_U1577 ( .A(DP_mult_207_n2187), .ZN(DP_mult_207_n2219) );
  XOR2_X1 DP_mult_207_U1576 ( .A(DP_coeffs_ff_int[45]), .B(
        DP_coeffs_ff_int[46]), .Z(DP_mult_207_n2083) );
  NAND3_X1 DP_mult_207_U1575 ( .A1(DP_mult_207_n2070), .A2(DP_mult_207_n2071), 
        .A3(DP_mult_207_n2072), .ZN(DP_mult_207_n2001) );
  NAND3_X1 DP_mult_207_U1574 ( .A1(DP_mult_207_n2070), .A2(DP_mult_207_n2071), 
        .A3(DP_mult_207_n2072), .ZN(DP_mult_207_n2002) );
  CLKBUF_X1 DP_mult_207_U1573 ( .A(DP_mult_207_n581), .Z(DP_mult_207_n2000) );
  XNOR2_X1 DP_mult_207_U1572 ( .A(DP_coeffs_ff_int[43]), .B(DP_mult_207_n2274), 
        .ZN(DP_mult_207_n2066) );
  INV_X1 DP_mult_207_U1571 ( .A(DP_mult_207_n2254), .ZN(DP_mult_207_n2251) );
  INV_X4 DP_mult_207_U1570 ( .A(DP_mult_207_n1931), .ZN(DP_mult_207_n2317) );
  NAND3_X1 DP_mult_207_U1569 ( .A1(DP_mult_207_n1997), .A2(DP_mult_207_n1998), 
        .A3(DP_mult_207_n1999), .ZN(DP_mult_207_n994) );
  NAND2_X1 DP_mult_207_U1568 ( .A1(DP_mult_207_n1306), .A2(DP_mult_207_n1416), 
        .ZN(DP_mult_207_n1999) );
  NAND2_X1 DP_mult_207_U1567 ( .A1(DP_mult_207_n1328), .A2(DP_mult_207_n1416), 
        .ZN(DP_mult_207_n1998) );
  NAND2_X1 DP_mult_207_U1566 ( .A1(DP_mult_207_n1328), .A2(DP_mult_207_n1306), 
        .ZN(DP_mult_207_n1997) );
  XOR2_X1 DP_mult_207_U1565 ( .A(DP_mult_207_n1996), .B(DP_mult_207_n1328), 
        .Z(DP_mult_207_n995) );
  XOR2_X1 DP_mult_207_U1564 ( .A(DP_mult_207_n1306), .B(DP_mult_207_n1416), 
        .Z(DP_mult_207_n1996) );
  NAND3_X1 DP_mult_207_U1563 ( .A1(DP_mult_207_n2054), .A2(DP_mult_207_n2055), 
        .A3(DP_mult_207_n2056), .ZN(DP_mult_207_n1995) );
  BUF_X1 DP_mult_207_U1562 ( .A(DP_mult_207_n1298), .Z(DP_mult_207_n1994) );
  INV_X1 DP_mult_207_U1561 ( .A(DP_mult_207_n2192), .ZN(DP_mult_207_n2224) );
  INV_X1 DP_mult_207_U1560 ( .A(DP_mult_207_n2192), .ZN(DP_mult_207_n1993) );
  XNOR2_X1 DP_mult_207_U1559 ( .A(DP_coeffs_ff_int[37]), .B(DP_mult_207_n2291), 
        .ZN(DP_mult_207_n1812) );
  XNOR2_X1 DP_mult_207_U1558 ( .A(DP_coeffs_ff_int[45]), .B(DP_mult_207_n2268), 
        .ZN(DP_mult_207_n2084) );
  BUF_X1 DP_mult_207_U1557 ( .A(DP_mult_207_n2167), .Z(DP_mult_207_n1992) );
  BUF_X1 DP_mult_207_U1556 ( .A(DP_mult_207_n2223), .Z(DP_mult_207_n2198) );
  XOR2_X1 DP_mult_207_U1555 ( .A(DP_coeffs_ff_int[41]), .B(
        DP_coeffs_ff_int[42]), .Z(DP_mult_207_n2082) );
  XNOR2_X1 DP_mult_207_U1554 ( .A(DP_coeffs_ff_int[41]), .B(
        DP_coeffs_ff_int[42]), .ZN(DP_mult_207_n2047) );
  INV_X2 DP_mult_207_U1553 ( .A(DP_mult_207_n2316), .ZN(DP_mult_207_n2313) );
  INV_X1 DP_mult_207_U1552 ( .A(DP_mult_207_n2244), .ZN(DP_mult_207_n1991) );
  XNOR2_X1 DP_mult_207_U1551 ( .A(DP_coeffs_ff_int[43]), .B(DP_mult_207_n2269), 
        .ZN(DP_mult_207_n1990) );
  XNOR2_X1 DP_mult_207_U1550 ( .A(DP_mult_207_n1284), .B(DP_mult_207_n1438), 
        .ZN(DP_mult_207_n1989) );
  XNOR2_X1 DP_mult_207_U1549 ( .A(DP_mult_207_n2037), .B(DP_mult_207_n1989), 
        .ZN(DP_mult_207_n997) );
  INV_X2 DP_mult_207_U1548 ( .A(DP_mult_207_n2305), .ZN(DP_mult_207_n2057) );
  INV_X1 DP_mult_207_U1547 ( .A(DP_mult_207_n2102), .ZN(DP_mult_207_n2240) );
  XOR2_X1 DP_mult_207_U1546 ( .A(DP_coeffs_ff_int[35]), .B(
        DP_coeffs_ff_int[36]), .Z(DP_mult_207_n1988) );
  XOR2_X1 DP_mult_207_U1545 ( .A(DP_coeffs_ff_int[35]), .B(
        DP_coeffs_ff_int[36]), .Z(DP_mult_207_n1987) );
  AND2_X1 DP_mult_207_U1544 ( .A1(DP_mult_207_n663), .A2(DP_mult_207_n439), 
        .ZN(DP_mult_207_n1986) );
  XNOR2_X1 DP_mult_207_U1543 ( .A(DP_mult_207_n2212), .B(DP_mult_207_n1986), 
        .ZN(DP_pipe0_coeff_pipe01[12]) );
  NOR2_X1 DP_mult_207_U1542 ( .A1(DP_mult_207_n558), .A2(DP_mult_207_n563), 
        .ZN(DP_mult_207_n552) );
  INV_X1 DP_mult_207_U1541 ( .A(DP_mult_207_n1942), .ZN(DP_mult_207_n1985) );
  AND2_X1 DP_mult_207_U1540 ( .A1(DP_mult_207_n672), .A2(DP_mult_207_n535), 
        .ZN(DP_mult_207_n1983) );
  XNOR2_X1 DP_mult_207_U1539 ( .A(DP_mult_207_n536), .B(DP_mult_207_n1983), 
        .ZN(DP_pipe0_coeff_pipe01[3]) );
  AND2_X1 DP_mult_207_U1538 ( .A1(DP_mult_207_n1957), .A2(DP_mult_207_n559), 
        .ZN(DP_mult_207_n1982) );
  XNOR2_X1 DP_mult_207_U1537 ( .A(DP_mult_207_n560), .B(DP_mult_207_n1982), 
        .ZN(DP_pipe0_coeff_pipe01[0]) );
  AND2_X1 DP_mult_207_U1536 ( .A1(DP_mult_207_n2139), .A2(DP_mult_207_n543), 
        .ZN(DP_mult_207_n1981) );
  XNOR2_X1 DP_mult_207_U1535 ( .A(DP_mult_207_n544), .B(DP_mult_207_n1981), 
        .ZN(DP_pipe0_coeff_pipe01[2]) );
  AND2_X1 DP_mult_207_U1534 ( .A1(DP_mult_207_n2127), .A2(DP_mult_207_n550), 
        .ZN(DP_mult_207_n1980) );
  XNOR2_X1 DP_mult_207_U1533 ( .A(DP_mult_207_n551), .B(DP_mult_207_n1980), 
        .ZN(DP_pipe0_coeff_pipe01[1]) );
  OR2_X1 DP_mult_207_U1532 ( .A1(DP_mult_207_n1143), .A2(DP_mult_207_n1150), 
        .ZN(DP_mult_207_n1979) );
  OR2_X1 DP_mult_207_U1531 ( .A1(DP_mult_207_n1151), .A2(DP_mult_207_n1158), 
        .ZN(DP_mult_207_n1978) );
  AND2_X1 DP_mult_207_U1530 ( .A1(DP_mult_207_n1111), .A2(DP_mult_207_n1122), 
        .ZN(DP_mult_207_n1977) );
  AND2_X1 DP_mult_207_U1529 ( .A1(DP_mult_207_n1133), .A2(DP_mult_207_n1142), 
        .ZN(DP_mult_207_n1976) );
  AND2_X1 DP_mult_207_U1528 ( .A1(DP_mult_207_n1055), .A2(DP_mult_207_n1070), 
        .ZN(DP_mult_207_n1975) );
  AND2_X1 DP_mult_207_U1527 ( .A1(DP_mult_207_n1179), .A2(DP_mult_207_n1433), 
        .ZN(DP_mult_207_n1974) );
  AND2_X1 DP_mult_207_U1526 ( .A1(DP_mult_207_n1021), .A2(DP_mult_207_n1038), 
        .ZN(DP_mult_207_n1973) );
  AND2_X1 DP_mult_207_U1525 ( .A1(DP_mult_207_n1457), .A2(DP_mult_207_n1480), 
        .ZN(DP_mult_207_n1972) );
  AND2_X1 DP_mult_207_U1524 ( .A1(DP_mult_207_n1817), .A2(DP_mult_207_n2261), 
        .ZN(DP_mult_207_n1971) );
  AND2_X1 DP_mult_207_U1523 ( .A1(DP_mult_207_n1151), .A2(DP_mult_207_n1158), 
        .ZN(DP_mult_207_n1970) );
  AND2_X1 DP_mult_207_U1522 ( .A1(DP_mult_207_n1123), .A2(DP_mult_207_n1132), 
        .ZN(DP_mult_207_n1969) );
  AND2_X1 DP_mult_207_U1521 ( .A1(DP_mult_207_n1143), .A2(DP_mult_207_n1150), 
        .ZN(DP_mult_207_n1968) );
  OR2_X1 DP_mult_207_U1520 ( .A1(DP_mult_207_n1179), .A2(DP_mult_207_n1433), 
        .ZN(DP_mult_207_n1967) );
  AND2_X1 DP_mult_207_U1519 ( .A1(DP_mult_207_n1039), .A2(DP_mult_207_n1054), 
        .ZN(DP_mult_207_n1966) );
  OR2_X1 DP_mult_207_U1518 ( .A1(DP_mult_207_n1457), .A2(DP_mult_207_n1480), 
        .ZN(DP_mult_207_n1965) );
  AND2_X1 DP_mult_207_U1517 ( .A1(DP_mult_207_n1193), .A2(DP_mult_207_n1481), 
        .ZN(DP_mult_207_n1964) );
  NOR2_X1 DP_mult_207_U1516 ( .A1(DP_mult_207_n941), .A2(DP_mult_207_n962), 
        .ZN(DP_mult_207_n547) );
  NOR2_X1 DP_mult_207_U1515 ( .A1(DP_mult_207_n1099), .A2(DP_mult_207_n1110), 
        .ZN(DP_mult_207_n597) );
  NAND3_X1 DP_mult_207_U1514 ( .A1(DP_mult_207_n2132), .A2(DP_mult_207_n2133), 
        .A3(DP_mult_207_n2134), .ZN(DP_mult_207_n958) );
  BUF_X2 DP_mult_207_U1513 ( .A(DP_mult_207_n2232), .Z(DP_mult_207_n2203) );
  XNOR2_X1 DP_mult_207_U1512 ( .A(DP_coeffs_ff_int[45]), .B(DP_mult_207_n2273), 
        .ZN(DP_mult_207_n1816) );
  INV_X2 DP_mult_207_U1511 ( .A(DP_mult_207_n2210), .ZN(DP_mult_207_n2238) );
  INV_X1 DP_mult_207_U1510 ( .A(DP_mult_207_n2210), .ZN(DP_mult_207_n2237) );
  OR2_X2 DP_mult_207_U1509 ( .A1(DP_mult_207_n2102), .A2(DP_mult_207_n2052), 
        .ZN(DP_mult_207_n2046) );
  BUF_X1 DP_mult_207_U1508 ( .A(DP_mult_207_n874), .Z(DP_mult_207_n1963) );
  NAND3_X1 DP_mult_207_U1507 ( .A1(DP_mult_207_n1960), .A2(DP_mult_207_n1961), 
        .A3(DP_mult_207_n1962), .ZN(DP_mult_207_n806) );
  NAND2_X1 DP_mult_207_U1506 ( .A1(DP_mult_207_n811), .A2(DP_mult_207_n826), 
        .ZN(DP_mult_207_n1962) );
  NAND2_X1 DP_mult_207_U1505 ( .A1(DP_mult_207_n824), .A2(DP_mult_207_n826), 
        .ZN(DP_mult_207_n1961) );
  NAND2_X1 DP_mult_207_U1504 ( .A1(DP_mult_207_n824), .A2(DP_mult_207_n811), 
        .ZN(DP_mult_207_n1960) );
  XOR2_X1 DP_mult_207_U1503 ( .A(DP_mult_207_n824), .B(DP_mult_207_n1959), .Z(
        DP_mult_207_n807) );
  XOR2_X1 DP_mult_207_U1502 ( .A(DP_mult_207_n811), .B(DP_mult_207_n826), .Z(
        DP_mult_207_n1959) );
  CLKBUF_X1 DP_mult_207_U1501 ( .A(DP_mult_207_n2256), .Z(DP_mult_207_n1958)
         );
  XNOR2_X1 DP_mult_207_U1500 ( .A(DP_coeffs_ff_int[34]), .B(
        DP_coeffs_ff_int[33]), .ZN(DP_mult_207_n265) );
  XNOR2_X1 DP_mult_207_U1499 ( .A(DP_coeffs_ff_int[43]), .B(DP_mult_207_n2278), 
        .ZN(DP_mult_207_n1815) );
  OR2_X1 DP_mult_207_U1498 ( .A1(DP_mult_207_n963), .A2(DP_mult_207_n982), 
        .ZN(DP_mult_207_n1957) );
  INV_X1 DP_mult_207_U1497 ( .A(DP_mult_207_n2315), .ZN(DP_mult_207_n2312) );
  CLKBUF_X1 DP_mult_207_U1496 ( .A(DP_mult_207_n568), .Z(DP_mult_207_n2024) );
  NAND2_X1 DP_mult_207_U1495 ( .A1(DP_mult_207_n1955), .A2(DP_mult_207_n1956), 
        .ZN(DP_mult_207_n1436) );
  OR2_X1 DP_mult_207_U1494 ( .A1(DP_mult_207_n1734), .A2(DP_mult_207_n2259), 
        .ZN(DP_mult_207_n1956) );
  OR2_X1 DP_mult_207_U1493 ( .A1(DP_mult_207_n2105), .A2(DP_mult_207_n1735), 
        .ZN(DP_mult_207_n1955) );
  XNOR2_X1 DP_mult_207_U1492 ( .A(DP_coeffs_ff_int[45]), .B(
        DP_coeffs_ff_int[46]), .ZN(DP_mult_207_n1954) );
  INV_X1 DP_mult_207_U1491 ( .A(DP_mult_207_n519), .ZN(DP_mult_207_n1953) );
  CLKBUF_X1 DP_mult_207_U1490 ( .A(DP_mult_207_n532), .Z(DP_mult_207_n1952) );
  XOR2_X1 DP_mult_207_U1489 ( .A(DP_mult_207_n1938), .B(DP_coeffs_ff_int[37]), 
        .Z(DP_mult_207_n1951) );
  AND2_X2 DP_mult_207_U1488 ( .A1(DP_mult_207_n1806), .A2(DP_mult_207_n2185), 
        .ZN(DP_mult_207_n2209) );
  NOR2_X1 DP_mult_207_U1487 ( .A1(DP_mult_207_n1003), .A2(DP_mult_207_n1020), 
        .ZN(DP_mult_207_n1950) );
  NAND3_X1 DP_mult_207_U1486 ( .A1(DP_mult_207_n1947), .A2(DP_mult_207_n1948), 
        .A3(DP_mult_207_n1949), .ZN(DP_mult_207_n966) );
  NAND2_X1 DP_mult_207_U1485 ( .A1(DP_mult_207_n973), .A2(DP_mult_207_n990), 
        .ZN(DP_mult_207_n1949) );
  NAND2_X1 DP_mult_207_U1484 ( .A1(DP_mult_207_n988), .A2(DP_mult_207_n990), 
        .ZN(DP_mult_207_n1948) );
  NAND2_X1 DP_mult_207_U1483 ( .A1(DP_mult_207_n988), .A2(DP_mult_207_n973), 
        .ZN(DP_mult_207_n1947) );
  XOR2_X1 DP_mult_207_U1482 ( .A(DP_mult_207_n988), .B(DP_mult_207_n1946), .Z(
        DP_mult_207_n967) );
  XOR2_X1 DP_mult_207_U1481 ( .A(DP_mult_207_n973), .B(DP_mult_207_n990), .Z(
        DP_mult_207_n1946) );
  INV_X2 DP_mult_207_U1480 ( .A(DP_mult_207_n2254), .ZN(DP_mult_207_n2252) );
  INV_X1 DP_mult_207_U1479 ( .A(DP_mult_207_n2252), .ZN(DP_mult_207_n1945) );
  INV_X1 DP_mult_207_U1478 ( .A(DP_mult_207_n2240), .ZN(DP_mult_207_n1944) );
  INV_X1 DP_mult_207_U1477 ( .A(DP_mult_207_n2084), .ZN(DP_mult_207_n1943) );
  OR2_X1 DP_mult_207_U1476 ( .A1(DP_mult_207_n558), .A2(DP_mult_207_n563), 
        .ZN(DP_mult_207_n1942) );
  INV_X2 DP_mult_207_U1475 ( .A(DP_mult_207_n2284), .ZN(DP_mult_207_n2281) );
  XOR2_X1 DP_mult_207_U1474 ( .A(DP_coeffs_ff_int[35]), .B(
        DP_coeffs_ff_int[34]), .Z(DP_mult_207_n1811) );
  XNOR2_X1 DP_mult_207_U1473 ( .A(DP_mult_207_n921), .B(DP_mult_207_n2101), 
        .ZN(DP_mult_207_n1941) );
  CLKBUF_X1 DP_mult_207_U1472 ( .A(DP_mult_207_n547), .Z(DP_mult_207_n1940) );
  XNOR2_X1 DP_mult_207_U1471 ( .A(DP_coeffs_ff_int[31]), .B(DP_mult_207_n2305), 
        .ZN(DP_mult_207_n1809) );
  CLKBUF_X1 DP_mult_207_U1470 ( .A(DP_coeffs_ff_int[30]), .Z(DP_mult_207_n1939) );
  OR2_X2 DP_mult_207_U1469 ( .A1(DP_mult_207_n1021), .A2(DP_mult_207_n1038), 
        .ZN(DP_mult_207_n2169) );
  XNOR2_X1 DP_mult_207_U1468 ( .A(DP_coeffs_ff_int[33]), .B(DP_mult_207_n2301), 
        .ZN(DP_mult_207_n1810) );
  CLKBUF_X1 DP_mult_207_U1467 ( .A(DP_coeffs_ff_int[38]), .Z(DP_mult_207_n1938) );
  BUF_X2 DP_mult_207_U1466 ( .A(DP_mult_207_n2230), .Z(DP_mult_207_n2197) );
  XNOR2_X1 DP_mult_207_U1465 ( .A(DP_coeffs_ff_int[25]), .B(
        DP_coeffs_ff_int[26]), .ZN(DP_mult_207_n2185) );
  BUF_X2 DP_mult_207_U1464 ( .A(DP_mult_207_n2185), .Z(DP_mult_207_n1937) );
  NAND3_X1 DP_mult_207_U1463 ( .A1(DP_mult_207_n1934), .A2(DP_mult_207_n1935), 
        .A3(DP_mult_207_n1936), .ZN(DP_mult_207_n796) );
  NAND2_X1 DP_mult_207_U1462 ( .A1(DP_mult_207_n1274), .A2(DP_mult_207_n1296), 
        .ZN(DP_mult_207_n1936) );
  NAND2_X1 DP_mult_207_U1461 ( .A1(DP_mult_207_n818), .A2(DP_mult_207_n1296), 
        .ZN(DP_mult_207_n1935) );
  NAND2_X1 DP_mult_207_U1460 ( .A1(DP_mult_207_n818), .A2(DP_mult_207_n1274), 
        .ZN(DP_mult_207_n1934) );
  XOR2_X1 DP_mult_207_U1459 ( .A(DP_mult_207_n818), .B(DP_mult_207_n1933), .Z(
        DP_mult_207_n797) );
  XOR2_X1 DP_mult_207_U1458 ( .A(DP_mult_207_n1274), .B(DP_mult_207_n1296), 
        .Z(DP_mult_207_n1933) );
  CLKBUF_X1 DP_mult_207_U1457 ( .A(DP_mult_207_n839), .Z(DP_mult_207_n1932) );
  XOR2_X1 DP_mult_207_U1456 ( .A(DP_coeffs_ff_int[29]), .B(
        DP_coeffs_ff_int[28]), .Z(DP_mult_207_n1808) );
  INV_X1 DP_mult_207_U1455 ( .A(DP_coeffs_ff_int[24]), .ZN(DP_mult_207_n1931)
         );
  INV_X1 DP_mult_207_U1454 ( .A(DP_mult_207_n2047), .ZN(DP_mult_207_n1930) );
  INV_X2 DP_mult_207_U1453 ( .A(DP_mult_207_n2310), .ZN(DP_mult_207_n2308) );
  XOR2_X2 DP_mult_207_U1452 ( .A(DP_coeffs_ff_int[27]), .B(
        DP_coeffs_ff_int[28]), .Z(DP_mult_207_n2102) );
  CLKBUF_X1 DP_mult_207_U1451 ( .A(DP_mult_207_n889), .Z(DP_mult_207_n1929) );
  AND2_X2 DP_mult_207_U1450 ( .A1(DP_mult_207_n1808), .A2(DP_mult_207_n2128), 
        .ZN(DP_mult_207_n1984) );
  INV_X1 DP_mult_207_U1449 ( .A(DP_mult_207_n537), .ZN(DP_mult_207_n536) );
  XNOR2_X1 DP_mult_207_U1448 ( .A(DP_coeffs_ff_int[27]), .B(
        DP_coeffs_ff_int[26]), .ZN(DP_mult_207_n2052) );
  HA_X1 DP_mult_207_U798 ( .A(DP_mult_207_n1456), .B(DP_mult_207_n1479), .CO(
        DP_mult_207_n1180), .S(DP_mult_207_n1181) );
  FA_X1 DP_mult_207_U797 ( .A(DP_mult_207_n1455), .B(DP_mult_207_n1478), .CI(
        DP_mult_207_n1180), .CO(DP_mult_207_n1178), .S(DP_mult_207_n1179) );
  HA_X1 DP_mult_207_U796 ( .A(DP_mult_207_n1432), .B(DP_mult_207_n1477), .CO(
        DP_mult_207_n1176), .S(DP_mult_207_n1177) );
  FA_X1 DP_mult_207_U795 ( .A(DP_mult_207_n1191), .B(DP_mult_207_n1454), .CI(
        DP_mult_207_n1177), .CO(DP_mult_207_n1174), .S(DP_mult_207_n1175) );
  FA_X1 DP_mult_207_U794 ( .A(DP_mult_207_n1476), .B(DP_mult_207_n1453), .CI(
        DP_mult_207_n1431), .CO(DP_mult_207_n1172), .S(DP_mult_207_n1173) );
  FA_X1 DP_mult_207_U793 ( .A(DP_mult_207_n1409), .B(DP_mult_207_n1176), .CI(
        DP_mult_207_n1173), .CO(DP_mult_207_n1170), .S(DP_mult_207_n1171) );
  HA_X1 DP_mult_207_U792 ( .A(DP_mult_207_n1408), .B(DP_mult_207_n1430), .CO(
        DP_mult_207_n1168), .S(DP_mult_207_n1169) );
  FA_X1 DP_mult_207_U791 ( .A(DP_mult_207_n1452), .B(DP_mult_207_n1475), .CI(
        DP_mult_207_n1190), .CO(DP_mult_207_n1166), .S(DP_mult_207_n1167) );
  FA_X1 DP_mult_207_U790 ( .A(DP_mult_207_n1172), .B(DP_mult_207_n1169), .CI(
        DP_mult_207_n1167), .CO(DP_mult_207_n1164), .S(DP_mult_207_n1165) );
  FA_X1 DP_mult_207_U789 ( .A(DP_mult_207_n1451), .B(DP_mult_207_n1474), .CI(
        DP_mult_207_n1407), .CO(DP_mult_207_n1162), .S(DP_mult_207_n1163) );
  FA_X1 DP_mult_207_U788 ( .A(DP_mult_207_n1168), .B(DP_mult_207_n1429), .CI(
        DP_mult_207_n1166), .CO(DP_mult_207_n1160), .S(DP_mult_207_n1161) );
  FA_X1 DP_mult_207_U787 ( .A(DP_mult_207_n1163), .B(DP_mult_207_n1385), .CI(
        DP_mult_207_n1164), .CO(DP_mult_207_n1158), .S(DP_mult_207_n1159) );
  HA_X1 DP_mult_207_U786 ( .A(DP_mult_207_n1384), .B(DP_mult_207_n1406), .CO(
        DP_mult_207_n1156), .S(DP_mult_207_n1157) );
  FA_X1 DP_mult_207_U785 ( .A(DP_mult_207_n1450), .B(DP_mult_207_n1428), .CI(
        DP_mult_207_n1189), .CO(DP_mult_207_n1154), .S(DP_mult_207_n1155) );
  FA_X1 DP_mult_207_U784 ( .A(DP_mult_207_n1157), .B(DP_mult_207_n1473), .CI(
        DP_mult_207_n1162), .CO(DP_mult_207_n1152), .S(DP_mult_207_n1153) );
  FA_X1 DP_mult_207_U783 ( .A(DP_mult_207_n1160), .B(DP_mult_207_n1155), .CI(
        DP_mult_207_n1153), .CO(DP_mult_207_n1150), .S(DP_mult_207_n1151) );
  FA_X1 DP_mult_207_U782 ( .A(DP_mult_207_n1383), .B(DP_mult_207_n1472), .CI(
        DP_mult_207_n1405), .CO(DP_mult_207_n1148), .S(DP_mult_207_n1149) );
  FA_X1 DP_mult_207_U781 ( .A(DP_mult_207_n1427), .B(DP_mult_207_n1449), .CI(
        DP_mult_207_n1156), .CO(DP_mult_207_n1146), .S(DP_mult_207_n1147) );
  FA_X1 DP_mult_207_U780 ( .A(DP_mult_207_n1361), .B(DP_mult_207_n1154), .CI(
        DP_mult_207_n1149), .CO(DP_mult_207_n1144), .S(DP_mult_207_n1145) );
  FA_X1 DP_mult_207_U779 ( .A(DP_mult_207_n1152), .B(DP_mult_207_n1147), .CI(
        DP_mult_207_n1145), .CO(DP_mult_207_n1142), .S(DP_mult_207_n1143) );
  HA_X1 DP_mult_207_U778 ( .A(DP_mult_207_n1360), .B(DP_mult_207_n1382), .CO(
        DP_mult_207_n1140), .S(DP_mult_207_n1141) );
  FA_X1 DP_mult_207_U776 ( .A(DP_mult_207_n1404), .B(DP_mult_207_n1448), .CI(
        DP_mult_207_n1141), .CO(DP_mult_207_n1136), .S(DP_mult_207_n1137) );
  FA_X1 DP_mult_207_U775 ( .A(DP_mult_207_n1146), .B(DP_mult_207_n1148), .CI(
        DP_mult_207_n1139), .CO(DP_mult_207_n1134), .S(DP_mult_207_n1135) );
  FA_X1 DP_mult_207_U774 ( .A(DP_mult_207_n1144), .B(DP_mult_207_n1137), .CI(
        DP_mult_207_n1135), .CO(DP_mult_207_n1132), .S(DP_mult_207_n1133) );
  FA_X1 DP_mult_207_U773 ( .A(DP_mult_207_n1359), .B(DP_mult_207_n1381), .CI(
        DP_mult_207_n1470), .CO(DP_mult_207_n1130), .S(DP_mult_207_n1131) );
  FA_X1 DP_mult_207_U772 ( .A(DP_mult_207_n1425), .B(DP_mult_207_n1447), .CI(
        DP_mult_207_n1403), .CO(DP_mult_207_n1128), .S(DP_mult_207_n1129) );
  FA_X1 DP_mult_207_U770 ( .A(DP_mult_207_n1131), .B(DP_mult_207_n1129), .CI(
        DP_mult_207_n1136), .CO(DP_mult_207_n1124), .S(DP_mult_207_n1125) );
  FA_X1 DP_mult_207_U769 ( .A(DP_mult_207_n1127), .B(DP_mult_207_n1134), .CI(
        DP_mult_207_n1125), .CO(DP_mult_207_n1122), .S(DP_mult_207_n1123) );
  HA_X1 DP_mult_207_U768 ( .A(DP_mult_207_n1336), .B(DP_mult_207_n1358), .CO(
        DP_mult_207_n1120), .S(DP_mult_207_n1121) );
  FA_X1 DP_mult_207_U767 ( .A(DP_mult_207_n1380), .B(DP_mult_207_n1402), .CI(
        DP_mult_207_n1187), .CO(DP_mult_207_n1118), .S(DP_mult_207_n1119) );
  FA_X1 DP_mult_207_U766 ( .A(DP_mult_207_n1424), .B(DP_mult_207_n1469), .CI(
        DP_mult_207_n1446), .CO(DP_mult_207_n1116), .S(DP_mult_207_n1117) );
  FA_X1 DP_mult_207_U765 ( .A(DP_mult_207_n1130), .B(DP_mult_207_n1121), .CI(
        DP_mult_207_n1128), .CO(DP_mult_207_n1114), .S(DP_mult_207_n1115) );
  FA_X1 DP_mult_207_U764 ( .A(DP_mult_207_n1119), .B(DP_mult_207_n1117), .CI(
        DP_mult_207_n1126), .CO(DP_mult_207_n1112), .S(DP_mult_207_n1113) );
  FA_X1 DP_mult_207_U763 ( .A(DP_mult_207_n1124), .B(DP_mult_207_n1115), .CI(
        DP_mult_207_n1113), .CO(DP_mult_207_n1110), .S(DP_mult_207_n1111) );
  FA_X1 DP_mult_207_U762 ( .A(DP_mult_207_n1335), .B(DP_mult_207_n1468), .CI(
        DP_mult_207_n1357), .CO(DP_mult_207_n1108), .S(DP_mult_207_n1109) );
  FA_X1 DP_mult_207_U761 ( .A(DP_mult_207_n1379), .B(DP_mult_207_n1445), .CI(
        DP_mult_207_n1401), .CO(DP_mult_207_n1106), .S(DP_mult_207_n1107) );
  FA_X1 DP_mult_207_U760 ( .A(DP_mult_207_n1120), .B(DP_mult_207_n1423), .CI(
        DP_mult_207_n1118), .CO(DP_mult_207_n1104), .S(DP_mult_207_n1105) );
  FA_X1 DP_mult_207_U759 ( .A(DP_mult_207_n1313), .B(DP_mult_207_n1116), .CI(
        DP_mult_207_n1107), .CO(DP_mult_207_n1102), .S(DP_mult_207_n1103) );
  FA_X1 DP_mult_207_U758 ( .A(DP_mult_207_n1114), .B(DP_mult_207_n1109), .CI(
        DP_mult_207_n1105), .CO(DP_mult_207_n1100), .S(DP_mult_207_n1101) );
  FA_X1 DP_mult_207_U757 ( .A(DP_mult_207_n1103), .B(DP_mult_207_n1112), .CI(
        DP_mult_207_n1101), .CO(DP_mult_207_n1098), .S(DP_mult_207_n1099) );
  HA_X1 DP_mult_207_U756 ( .A(DP_mult_207_n1334), .B(DP_mult_207_n1312), .CO(
        DP_mult_207_n1096), .S(DP_mult_207_n1097) );
  FA_X1 DP_mult_207_U755 ( .A(DP_mult_207_n1186), .B(DP_mult_207_n1400), .CI(
        DP_mult_207_n1467), .CO(DP_mult_207_n1094), .S(DP_mult_207_n1095) );
  FA_X1 DP_mult_207_U754 ( .A(DP_mult_207_n1444), .B(DP_mult_207_n1378), .CI(
        DP_mult_207_n1356), .CO(DP_mult_207_n1092), .S(DP_mult_207_n1093) );
  FA_X1 DP_mult_207_U753 ( .A(DP_mult_207_n1097), .B(DP_mult_207_n1422), .CI(
        DP_mult_207_n1108), .CO(DP_mult_207_n1090), .S(DP_mult_207_n1091) );
  FA_X1 DP_mult_207_U752 ( .A(DP_mult_207_n1093), .B(DP_mult_207_n1106), .CI(
        DP_mult_207_n1095), .CO(DP_mult_207_n1088), .S(DP_mult_207_n1089) );
  FA_X1 DP_mult_207_U751 ( .A(DP_mult_207_n1102), .B(DP_mult_207_n1104), .CI(
        DP_mult_207_n1091), .CO(DP_mult_207_n1086), .S(DP_mult_207_n1087) );
  FA_X1 DP_mult_207_U750 ( .A(DP_mult_207_n1100), .B(DP_mult_207_n1089), .CI(
        DP_mult_207_n1087), .CO(DP_mult_207_n1084), .S(DP_mult_207_n1085) );
  FA_X1 DP_mult_207_U749 ( .A(DP_mult_207_n1311), .B(DP_mult_207_n1466), .CI(
        DP_mult_207_n1333), .CO(DP_mult_207_n1082), .S(DP_mult_207_n1083) );
  FA_X1 DP_mult_207_U748 ( .A(DP_mult_207_n1355), .B(DP_mult_207_n1443), .CI(
        DP_mult_207_n1377), .CO(DP_mult_207_n1080), .S(DP_mult_207_n1081) );
  FA_X1 DP_mult_207_U747 ( .A(DP_mult_207_n1399), .B(DP_mult_207_n1096), .CI(
        DP_mult_207_n1421), .CO(DP_mult_207_n1078), .S(DP_mult_207_n1079) );
  FA_X1 DP_mult_207_U746 ( .A(DP_mult_207_n1092), .B(DP_mult_207_n1094), .CI(
        DP_mult_207_n1289), .CO(DP_mult_207_n1076), .S(DP_mult_207_n1077) );
  FA_X1 DP_mult_207_U745 ( .A(DP_mult_207_n1083), .B(DP_mult_207_n1081), .CI(
        DP_mult_207_n1079), .CO(DP_mult_207_n1074), .S(DP_mult_207_n1075) );
  FA_X1 DP_mult_207_U744 ( .A(DP_mult_207_n1088), .B(DP_mult_207_n1090), .CI(
        DP_mult_207_n1077), .CO(DP_mult_207_n1072), .S(DP_mult_207_n1073) );
  FA_X1 DP_mult_207_U743 ( .A(DP_mult_207_n1086), .B(DP_mult_207_n1075), .CI(
        DP_mult_207_n1073), .CO(DP_mult_207_n1070), .S(DP_mult_207_n1071) );
  HA_X1 DP_mult_207_U742 ( .A(DP_mult_207_n1288), .B(DP_mult_207_n1310), .CO(
        DP_mult_207_n1068), .S(DP_mult_207_n1069) );
  FA_X1 DP_mult_207_U741 ( .A(DP_mult_207_n1465), .B(DP_mult_207_n1376), .CI(
        DP_mult_207_n1185), .CO(DP_mult_207_n1066), .S(DP_mult_207_n1067) );
  FA_X1 DP_mult_207_U740 ( .A(DP_mult_207_n1442), .B(DP_mult_207_n1354), .CI(
        DP_mult_207_n1332), .CO(DP_mult_207_n1064), .S(DP_mult_207_n1065) );
  FA_X1 DP_mult_207_U739 ( .A(DP_mult_207_n1398), .B(DP_mult_207_n1420), .CI(
        DP_mult_207_n1069), .CO(DP_mult_207_n1062), .S(DP_mult_207_n1063) );
  FA_X1 DP_mult_207_U738 ( .A(DP_mult_207_n1080), .B(DP_mult_207_n1082), .CI(
        DP_mult_207_n1078), .CO(DP_mult_207_n1060), .S(DP_mult_207_n1061) );
  FA_X1 DP_mult_207_U737 ( .A(DP_mult_207_n1067), .B(DP_mult_207_n1065), .CI(
        DP_mult_207_n1076), .CO(DP_mult_207_n1058), .S(DP_mult_207_n1059) );
  FA_X1 DP_mult_207_U736 ( .A(DP_mult_207_n1061), .B(DP_mult_207_n1063), .CI(
        DP_mult_207_n1074), .CO(DP_mult_207_n1056), .S(DP_mult_207_n1057) );
  FA_X1 DP_mult_207_U735 ( .A(DP_mult_207_n1072), .B(DP_mult_207_n1059), .CI(
        DP_mult_207_n1057), .CO(DP_mult_207_n1054), .S(DP_mult_207_n1055) );
  FA_X1 DP_mult_207_U734 ( .A(DP_mult_207_n1309), .B(DP_mult_207_n1464), .CI(
        DP_mult_207_n1287), .CO(DP_mult_207_n1052), .S(DP_mult_207_n1053) );
  FA_X1 DP_mult_207_U733 ( .A(DP_mult_207_n1331), .B(DP_mult_207_n1353), .CI(
        DP_mult_207_n1375), .CO(DP_mult_207_n1050), .S(DP_mult_207_n1051) );
  FA_X1 DP_mult_207_U732 ( .A(DP_mult_207_n1397), .B(DP_mult_207_n1441), .CI(
        DP_mult_207_n1419), .CO(DP_mult_207_n1048), .S(DP_mult_207_n1049) );
  FA_X1 DP_mult_207_U731 ( .A(DP_mult_207_n1064), .B(DP_mult_207_n1068), .CI(
        DP_mult_207_n1066), .CO(DP_mult_207_n1046), .S(DP_mult_207_n1047) );
  FA_X1 DP_mult_207_U730 ( .A(DP_mult_207_n1049), .B(DP_mult_207_n1265), .CI(
        DP_mult_207_n1051), .CO(DP_mult_207_n1044), .S(DP_mult_207_n1045) );
  FA_X1 DP_mult_207_U729 ( .A(DP_mult_207_n1062), .B(DP_mult_207_n1053), .CI(
        DP_mult_207_n1060), .CO(DP_mult_207_n1042), .S(DP_mult_207_n1043) );
  FA_X1 DP_mult_207_U728 ( .A(DP_mult_207_n1058), .B(DP_mult_207_n1047), .CI(
        DP_mult_207_n1045), .CO(DP_mult_207_n1040), .S(DP_mult_207_n1041) );
  HA_X1 DP_mult_207_U726 ( .A(DP_mult_207_n1264), .B(DP_mult_207_n1286), .CO(
        DP_mult_207_n1036), .S(DP_mult_207_n1037) );
  FA_X1 DP_mult_207_U725 ( .A(DP_mult_207_n1308), .B(DP_mult_207_n1184), .CI(
        DP_mult_207_n1374), .CO(DP_mult_207_n1034), .S(DP_mult_207_n1035) );
  FA_X1 DP_mult_207_U724 ( .A(DP_mult_207_n1330), .B(DP_mult_207_n1396), .CI(
        DP_mult_207_n1463), .CO(DP_mult_207_n1032), .S(DP_mult_207_n1033) );
  FA_X1 DP_mult_207_U723 ( .A(DP_mult_207_n1418), .B(DP_mult_207_n1440), .CI(
        DP_mult_207_n1352), .CO(DP_mult_207_n1030), .S(DP_mult_207_n1031) );
  FA_X1 DP_mult_207_U722 ( .A(DP_mult_207_n1052), .B(DP_mult_207_n1037), .CI(
        DP_mult_207_n1050), .CO(DP_mult_207_n1028), .S(DP_mult_207_n1029) );
  FA_X1 DP_mult_207_U721 ( .A(DP_mult_207_n1031), .B(DP_mult_207_n1048), .CI(
        DP_mult_207_n1033), .CO(DP_mult_207_n1026), .S(DP_mult_207_n1027) );
  FA_X1 DP_mult_207_U720 ( .A(DP_mult_207_n1046), .B(DP_mult_207_n1035), .CI(
        DP_mult_207_n1029), .CO(DP_mult_207_n1024), .S(DP_mult_207_n1025) );
  FA_X1 DP_mult_207_U719 ( .A(DP_mult_207_n1027), .B(DP_mult_207_n1044), .CI(
        DP_mult_207_n1042), .CO(DP_mult_207_n1022), .S(DP_mult_207_n1023) );
  FA_X1 DP_mult_207_U717 ( .A(DP_mult_207_n1351), .B(DP_mult_207_n1263), .CI(
        DP_mult_207_n1285), .CO(DP_mult_207_n1018), .S(DP_mult_207_n1019) );
  FA_X1 DP_mult_207_U716 ( .A(DP_mult_207_n1307), .B(DP_mult_207_n1373), .CI(
        DP_mult_207_n1329), .CO(DP_mult_207_n1016), .S(DP_mult_207_n1017) );
  FA_X1 DP_mult_207_U715 ( .A(DP_mult_207_n1395), .B(DP_mult_207_n1462), .CI(
        DP_mult_207_n1417), .CO(DP_mult_207_n1014), .S(DP_mult_207_n1015) );
  FA_X1 DP_mult_207_U714 ( .A(DP_mult_207_n1036), .B(DP_mult_207_n1439), .CI(
        DP_mult_207_n1032), .CO(DP_mult_207_n1012), .S(DP_mult_207_n1013) );
  FA_X1 DP_mult_207_U713 ( .A(DP_mult_207_n1030), .B(DP_mult_207_n1034), .CI(
        DP_mult_207_n1241), .CO(DP_mult_207_n1010), .S(DP_mult_207_n1011) );
  FA_X1 DP_mult_207_U712 ( .A(DP_mult_207_n1019), .B(DP_mult_207_n1015), .CI(
        DP_mult_207_n1017), .CO(DP_mult_207_n1008), .S(DP_mult_207_n1009) );
  FA_X1 DP_mult_207_U711 ( .A(DP_mult_207_n1013), .B(DP_mult_207_n1028), .CI(
        DP_mult_207_n1026), .CO(DP_mult_207_n1006), .S(DP_mult_207_n1007) );
  FA_X1 DP_mult_207_U710 ( .A(DP_mult_207_n1009), .B(DP_mult_207_n1011), .CI(
        DP_mult_207_n1024), .CO(DP_mult_207_n1004), .S(DP_mult_207_n1005) );
  FA_X1 DP_mult_207_U709 ( .A(DP_mult_207_n1022), .B(DP_mult_207_n1007), .CI(
        DP_mult_207_n1005), .CO(DP_mult_207_n1002), .S(DP_mult_207_n1003) );
  HA_X1 DP_mult_207_U708 ( .A(DP_mult_207_n1240), .B(DP_mult_207_n1262), .CO(
        DP_mult_207_n1000), .S(DP_mult_207_n1001) );
  FA_X1 DP_mult_207_U707 ( .A(DP_mult_207_n1461), .B(DP_mult_207_n1350), .CI(
        DP_mult_207_n1183), .CO(DP_mult_207_n998), .S(DP_mult_207_n999) );
  FA_X1 DP_mult_207_U704 ( .A(DP_mult_207_n1001), .B(DP_mult_207_n1394), .CI(
        DP_mult_207_n1018), .CO(DP_mult_207_n992), .S(DP_mult_207_n993) );
  FA_X1 DP_mult_207_U703 ( .A(DP_mult_207_n1014), .B(DP_mult_207_n1016), .CI(
        DP_mult_207_n995), .CO(DP_mult_207_n990), .S(DP_mult_207_n991) );
  FA_X1 DP_mult_207_U702 ( .A(DP_mult_207_n999), .B(DP_mult_207_n997), .CI(
        DP_mult_207_n1012), .CO(DP_mult_207_n988), .S(DP_mult_207_n989) );
  FA_X1 DP_mult_207_U701 ( .A(DP_mult_207_n993), .B(DP_mult_207_n1010), .CI(
        DP_mult_207_n1008), .CO(DP_mult_207_n986), .S(DP_mult_207_n987) );
  FA_X1 DP_mult_207_U700 ( .A(DP_mult_207_n989), .B(DP_mult_207_n991), .CI(
        DP_mult_207_n1006), .CO(DP_mult_207_n984), .S(DP_mult_207_n985) );
  FA_X1 DP_mult_207_U699 ( .A(DP_mult_207_n1004), .B(DP_mult_207_n987), .CI(
        DP_mult_207_n985), .CO(DP_mult_207_n982), .S(DP_mult_207_n983) );
  FA_X1 DP_mult_207_U698 ( .A(DP_mult_207_n1239), .B(DP_mult_207_n1349), .CI(
        DP_mult_207_n1261), .CO(DP_mult_207_n980), .S(DP_mult_207_n981) );
  FA_X1 DP_mult_207_U697 ( .A(DP_mult_207_n1460), .B(DP_mult_207_n1371), .CI(
        DP_mult_207_n1283), .CO(DP_mult_207_n978), .S(DP_mult_207_n979) );
  FA_X1 DP_mult_207_U696 ( .A(DP_mult_207_n1305), .B(DP_mult_207_n1327), .CI(
        DP_mult_207_n1437), .CO(DP_mult_207_n976), .S(DP_mult_207_n977) );
  FA_X1 DP_mult_207_U695 ( .A(DP_mult_207_n1000), .B(DP_mult_207_n1415), .CI(
        DP_mult_207_n1393), .CO(DP_mult_207_n974), .S(DP_mult_207_n975) );
  FA_X1 DP_mult_207_U693 ( .A(DP_mult_207_n977), .B(DP_mult_207_n998), .CI(
        DP_mult_207_n979), .CO(DP_mult_207_n970), .S(DP_mult_207_n971) );
  FA_X1 DP_mult_207_U692 ( .A(DP_mult_207_n992), .B(DP_mult_207_n981), .CI(
        DP_mult_207_n975), .CO(DP_mult_207_n968), .S(DP_mult_207_n969) );
  FA_X1 DP_mult_207_U690 ( .A(DP_mult_207_n969), .B(DP_mult_207_n971), .CI(
        DP_mult_207_n986), .CO(DP_mult_207_n964), .S(DP_mult_207_n965) );
  FA_X1 DP_mult_207_U689 ( .A(DP_mult_207_n984), .B(DP_mult_207_n967), .CI(
        DP_mult_207_n965), .CO(DP_mult_207_n962), .S(DP_mult_207_n963) );
  HA_X1 DP_mult_207_U688 ( .A(DP_mult_207_n1238), .B(DP_mult_207_n1216), .CO(
        DP_mult_207_n960), .S(DP_mult_207_n961) );
  FA_X1 DP_mult_207_U684 ( .A(DP_mult_207_n1326), .B(DP_mult_207_n1392), .CI(
        DP_mult_207_n961), .CO(DP_mult_207_n952), .S(DP_mult_207_n953) );
  FA_X1 DP_mult_207_U683 ( .A(DP_mult_207_n976), .B(DP_mult_207_n980), .CI(
        DP_mult_207_n978), .CO(DP_mult_207_n950), .S(DP_mult_207_n951) );
  FA_X1 DP_mult_207_U682 ( .A(DP_mult_207_n955), .B(DP_mult_207_n974), .CI(
        DP_mult_207_n957), .CO(DP_mult_207_n948), .S(DP_mult_207_n949) );
  FA_X1 DP_mult_207_U681 ( .A(DP_mult_207_n972), .B(DP_mult_207_n959), .CI(
        DP_mult_207_n953), .CO(DP_mult_207_n946), .S(DP_mult_207_n947) );
  FA_X1 DP_mult_207_U680 ( .A(DP_mult_207_n951), .B(DP_mult_207_n970), .CI(
        DP_mult_207_n968), .CO(DP_mult_207_n944), .S(DP_mult_207_n945) );
  FA_X1 DP_mult_207_U675 ( .A(DP_mult_207_n1259), .B(DP_mult_207_n1303), .CI(
        DP_mult_207_n1347), .CO(DP_mult_207_n936), .S(DP_mult_207_n937) );
  FA_X1 DP_mult_207_U674 ( .A(DP_mult_207_n1281), .B(DP_mult_207_n1369), .CI(
        DP_mult_207_n1391), .CO(DP_mult_207_n934), .S(DP_mult_207_n935) );
  FA_X1 DP_mult_207_U673 ( .A(DP_mult_207_n1325), .B(DP_mult_207_n1435), .CI(
        DP_mult_207_n1413), .CO(DP_mult_207_n932), .S(DP_mult_207_n933) );
  FA_X1 DP_mult_207_U672 ( .A(DP_mult_207_n939), .B(DP_mult_207_n960), .CI(
        DP_mult_207_n1458), .CO(DP_mult_207_n930), .S(DP_mult_207_n931) );
  FA_X1 DP_mult_207_U670 ( .A(DP_mult_207_n933), .B(DP_mult_207_n937), .CI(
        DP_mult_207_n952), .CO(DP_mult_207_n926), .S(DP_mult_207_n927) );
  FA_X1 DP_mult_207_U669 ( .A(DP_mult_207_n931), .B(DP_mult_207_n935), .CI(
        DP_mult_207_n950), .CO(DP_mult_207_n924), .S(DP_mult_207_n925) );
  FA_X1 DP_mult_207_U668 ( .A(DP_mult_207_n929), .B(DP_mult_207_n948), .CI(
        DP_mult_207_n946), .CO(DP_mult_207_n922), .S(DP_mult_207_n923) );
  FA_X1 DP_mult_207_U664 ( .A(DP_mult_207_n1214), .B(DP_mult_207_n917), .CI(
        DP_mult_207_n1302), .CO(DP_mult_207_n914), .S(DP_mult_207_n915) );
  FA_X1 DP_mult_207_U663 ( .A(DP_mult_207_n1258), .B(DP_mult_207_n1236), .CI(
        DP_mult_207_n1412), .CO(DP_mult_207_n912), .S(DP_mult_207_n913) );
  FA_X1 DP_mult_207_U662 ( .A(DP_mult_207_n1324), .B(DP_mult_207_n1346), .CI(
        DP_mult_207_n1280), .CO(DP_mult_207_n910), .S(DP_mult_207_n911) );
  FA_X1 DP_mult_207_U660 ( .A(DP_mult_207_n932), .B(DP_mult_207_n936), .CI(
        DP_mult_207_n934), .CO(DP_mult_207_n906), .S(DP_mult_207_n907) );
  FA_X1 DP_mult_207_U659 ( .A(DP_mult_207_n915), .B(DP_mult_207_n913), .CI(
        DP_mult_207_n911), .CO(DP_mult_207_n904), .S(DP_mult_207_n905) );
  FA_X1 DP_mult_207_U658 ( .A(DP_mult_207_n909), .B(DP_mult_207_n930), .CI(
        DP_mult_207_n928), .CO(DP_mult_207_n902), .S(DP_mult_207_n903) );
  FA_X1 DP_mult_207_U657 ( .A(DP_mult_207_n907), .B(DP_mult_207_n926), .CI(
        DP_mult_207_n905), .CO(DP_mult_207_n900), .S(DP_mult_207_n901) );
  FA_X1 DP_mult_207_U656 ( .A(DP_mult_207_n903), .B(DP_mult_207_n924), .CI(
        DP_mult_207_n922), .CO(DP_mult_207_n898), .S(DP_mult_207_n899) );
  FA_X1 DP_mult_207_U654 ( .A(DP_mult_207_n1235), .B(DP_mult_207_n1213), .CI(
        DP_mult_207_n1411), .CO(DP_mult_207_n894), .S(DP_mult_207_n895) );
  FA_X1 DP_mult_207_U653 ( .A(DP_mult_207_n916), .B(DP_mult_207_n1323), .CI(
        DP_mult_207_n1279), .CO(DP_mult_207_n892), .S(DP_mult_207_n893) );
  FA_X1 DP_mult_207_U652 ( .A(DP_mult_207_n1257), .B(DP_mult_207_n1345), .CI(
        DP_mult_207_n1301), .CO(DP_mult_207_n890), .S(DP_mult_207_n891) );
  FA_X1 DP_mult_207_U651 ( .A(DP_mult_207_n1367), .B(DP_mult_207_n1389), .CI(
        DP_mult_207_n1434), .CO(DP_mult_207_n888), .S(DP_mult_207_n889) );
  FA_X1 DP_mult_207_U650 ( .A(DP_mult_207_n910), .B(DP_mult_207_n914), .CI(
        DP_mult_207_n912), .CO(DP_mult_207_n886), .S(DP_mult_207_n887) );
  FA_X1 DP_mult_207_U649 ( .A(DP_mult_207_n891), .B(DP_mult_207_n908), .CI(
        DP_mult_207_n895), .CO(DP_mult_207_n884), .S(DP_mult_207_n885) );
  FA_X1 DP_mult_207_U647 ( .A(DP_mult_207_n887), .B(DP_mult_207_n904), .CI(
        DP_mult_207_n902), .CO(DP_mult_207_n880), .S(DP_mult_207_n881) );
  FA_X1 DP_mult_207_U646 ( .A(DP_mult_207_n883), .B(DP_mult_207_n885), .CI(
        DP_mult_207_n900), .CO(DP_mult_207_n878), .S(DP_mult_207_n879) );
  FA_X1 DP_mult_207_U645 ( .A(DP_mult_207_n898), .B(DP_mult_207_n881), .CI(
        DP_mult_207_n879), .CO(DP_mult_207_n876), .S(DP_mult_207_n877) );
  FA_X1 DP_mult_207_U643 ( .A(DP_mult_207_n1388), .B(DP_mult_207_n1278), .CI(
        DP_mult_207_n875), .CO(DP_mult_207_n872), .S(DP_mult_207_n873) );
  FA_X1 DP_mult_207_U642 ( .A(DP_mult_207_n1212), .B(DP_mult_207_n1366), .CI(
        DP_mult_207_n1344), .CO(DP_mult_207_n870), .S(DP_mult_207_n871) );
  FA_X1 DP_mult_207_U641 ( .A(DP_mult_207_n1322), .B(DP_mult_207_n1234), .CI(
        DP_mult_207_n1256), .CO(DP_mult_207_n868), .S(DP_mult_207_n869) );
  FA_X1 DP_mult_207_U640 ( .A(DP_mult_207_n894), .B(DP_mult_207_n1300), .CI(
        DP_mult_207_n892), .CO(DP_mult_207_n866), .S(DP_mult_207_n867) );
  FA_X1 DP_mult_207_U639 ( .A(DP_mult_207_n869), .B(DP_mult_207_n890), .CI(
        DP_mult_207_n871), .CO(DP_mult_207_n864), .S(DP_mult_207_n865) );
  FA_X1 DP_mult_207_U638 ( .A(DP_mult_207_n888), .B(DP_mult_207_n873), .CI(
        DP_mult_207_n886), .CO(DP_mult_207_n862), .S(DP_mult_207_n863) );
  FA_X1 DP_mult_207_U637 ( .A(DP_mult_207_n884), .B(DP_mult_207_n867), .CI(
        DP_mult_207_n865), .CO(DP_mult_207_n860), .S(DP_mult_207_n861) );
  FA_X1 DP_mult_207_U636 ( .A(DP_mult_207_n863), .B(DP_mult_207_n882), .CI(
        DP_mult_207_n880), .CO(DP_mult_207_n858), .S(DP_mult_207_n859) );
  FA_X1 DP_mult_207_U635 ( .A(DP_mult_207_n878), .B(DP_mult_207_n861), .CI(
        DP_mult_207_n859), .CO(DP_mult_207_n856), .S(DP_mult_207_n857) );
  FA_X1 DP_mult_207_U634 ( .A(DP_mult_207_n1233), .B(DP_mult_207_n1211), .CI(
        DP_mult_207_n1387), .CO(DP_mult_207_n854), .S(DP_mult_207_n855) );
  FA_X1 DP_mult_207_U633 ( .A(DP_mult_207_n1255), .B(DP_mult_207_n1321), .CI(
        DP_mult_207_n1963), .CO(DP_mult_207_n852), .S(DP_mult_207_n853) );
  FA_X1 DP_mult_207_U632 ( .A(DP_mult_207_n1343), .B(DP_mult_207_n1299), .CI(
        DP_mult_207_n1277), .CO(DP_mult_207_n850), .S(DP_mult_207_n851) );
  FA_X1 DP_mult_207_U631 ( .A(DP_mult_207_n1410), .B(DP_mult_207_n1365), .CI(
        DP_mult_207_n872), .CO(DP_mult_207_n848), .S(DP_mult_207_n849) );
  FA_X1 DP_mult_207_U629 ( .A(DP_mult_207_n855), .B(DP_mult_207_n853), .CI(
        DP_mult_207_n866), .CO(DP_mult_207_n844), .S(DP_mult_207_n845) );
  FA_X1 DP_mult_207_U627 ( .A(DP_mult_207_n845), .B(DP_mult_207_n847), .CI(
        DP_mult_207_n860), .CO(DP_mult_207_n840), .S(DP_mult_207_n841) );
  FA_X1 DP_mult_207_U626 ( .A(DP_mult_207_n858), .B(DP_mult_207_n843), .CI(
        DP_mult_207_n841), .CO(DP_mult_207_n838), .S(DP_mult_207_n839) );
  FA_X1 DP_mult_207_U624 ( .A(DP_mult_207_n1210), .B(DP_mult_207_n837), .CI(
        DP_mult_207_n1276), .CO(DP_mult_207_n834), .S(DP_mult_207_n835) );
  FA_X1 DP_mult_207_U623 ( .A(DP_mult_207_n1232), .B(DP_mult_207_n1364), .CI(
        DP_mult_207_n1342), .CO(DP_mult_207_n832), .S(DP_mult_207_n833) );
  FA_X1 DP_mult_207_U621 ( .A(DP_mult_207_n850), .B(DP_mult_207_n854), .CI(
        DP_mult_207_n852), .CO(DP_mult_207_n828), .S(DP_mult_207_n829) );
  FA_X1 DP_mult_207_U620 ( .A(DP_mult_207_n835), .B(DP_mult_207_n831), .CI(
        DP_mult_207_n833), .CO(DP_mult_207_n826), .S(DP_mult_207_n827) );
  FA_X1 DP_mult_207_U619 ( .A(DP_mult_207_n846), .B(DP_mult_207_n848), .CI(
        DP_mult_207_n829), .CO(DP_mult_207_n824), .S(DP_mult_207_n825) );
  FA_X1 DP_mult_207_U617 ( .A(DP_mult_207_n840), .B(DP_mult_207_n825), .CI(
        DP_mult_207_n823), .CO(DP_mult_207_n820), .S(DP_mult_207_n821) );
  FA_X1 DP_mult_207_U616 ( .A(DP_mult_207_n1209), .B(DP_mult_207_n1363), .CI(
        DP_mult_207_n836), .CO(DP_mult_207_n818), .S(DP_mult_207_n819) );
  FA_X1 DP_mult_207_U615 ( .A(DP_mult_207_n1231), .B(DP_mult_207_n1297), .CI(
        DP_mult_207_n1275), .CO(DP_mult_207_n816), .S(DP_mult_207_n817) );
  FA_X1 DP_mult_207_U614 ( .A(DP_mult_207_n1319), .B(DP_mult_207_n1253), .CI(
        DP_mult_207_n1341), .CO(DP_mult_207_n814), .S(DP_mult_207_n815) );
  FA_X1 DP_mult_207_U613 ( .A(DP_mult_207_n830), .B(DP_mult_207_n1386), .CI(
        DP_mult_207_n834), .CO(DP_mult_207_n812), .S(DP_mult_207_n813) );
  FA_X1 DP_mult_207_U612 ( .A(DP_mult_207_n815), .B(DP_mult_207_n832), .CI(
        DP_mult_207_n817), .CO(DP_mult_207_n810), .S(DP_mult_207_n811) );
  FA_X1 DP_mult_207_U611 ( .A(DP_mult_207_n828), .B(DP_mult_207_n819), .CI(
        DP_mult_207_n813), .CO(DP_mult_207_n808), .S(DP_mult_207_n809) );
  FA_X1 DP_mult_207_U609 ( .A(DP_mult_207_n807), .B(DP_mult_207_n809), .CI(
        DP_mult_207_n822), .CO(DP_mult_207_n804), .S(DP_mult_207_n805) );
  FA_X1 DP_mult_207_U607 ( .A(DP_mult_207_n1340), .B(DP_mult_207_n1252), .CI(
        DP_mult_207_n803), .CO(DP_mult_207_n800), .S(DP_mult_207_n801) );
  FA_X1 DP_mult_207_U606 ( .A(DP_mult_207_n1208), .B(DP_mult_207_n1318), .CI(
        DP_mult_207_n1230), .CO(DP_mult_207_n798), .S(DP_mult_207_n799) );
  FA_X1 DP_mult_207_U604 ( .A(DP_mult_207_n814), .B(DP_mult_207_n816), .CI(
        DP_mult_207_n799), .CO(DP_mult_207_n794), .S(DP_mult_207_n795) );
  FA_X1 DP_mult_207_U603 ( .A(DP_mult_207_n797), .B(DP_mult_207_n801), .CI(
        DP_mult_207_n812), .CO(DP_mult_207_n792), .S(DP_mult_207_n793) );
  FA_X1 DP_mult_207_U601 ( .A(DP_mult_207_n806), .B(DP_mult_207_n793), .CI(
        DP_mult_207_n791), .CO(DP_mult_207_n788), .S(DP_mult_207_n789) );
  FA_X1 DP_mult_207_U600 ( .A(DP_mult_207_n1251), .B(DP_mult_207_n1207), .CI(
        DP_mult_207_n802), .CO(DP_mult_207_n786), .S(DP_mult_207_n787) );
  FA_X1 DP_mult_207_U599 ( .A(DP_mult_207_n1273), .B(DP_mult_207_n1317), .CI(
        DP_mult_207_n1295), .CO(DP_mult_207_n784), .S(DP_mult_207_n785) );
  FA_X1 DP_mult_207_U598 ( .A(DP_mult_207_n1339), .B(DP_mult_207_n1229), .CI(
        DP_mult_207_n1362), .CO(DP_mult_207_n782), .S(DP_mult_207_n783) );
  FA_X1 DP_mult_207_U597 ( .A(DP_mult_207_n798), .B(DP_mult_207_n800), .CI(
        DP_mult_207_n785), .CO(DP_mult_207_n780), .S(DP_mult_207_n781) );
  FA_X1 DP_mult_207_U596 ( .A(DP_mult_207_n796), .B(DP_mult_207_n787), .CI(
        DP_mult_207_n783), .CO(DP_mult_207_n778), .S(DP_mult_207_n779) );
  FA_X1 DP_mult_207_U595 ( .A(DP_mult_207_n781), .B(DP_mult_207_n794), .CI(
        DP_mult_207_n792), .CO(DP_mult_207_n776), .S(DP_mult_207_n777) );
  FA_X1 DP_mult_207_U594 ( .A(DP_mult_207_n790), .B(DP_mult_207_n779), .CI(
        DP_mult_207_n777), .CO(DP_mult_207_n774), .S(DP_mult_207_n775) );
  FA_X1 DP_mult_207_U592 ( .A(DP_mult_207_n1316), .B(DP_mult_207_n1250), .CI(
        DP_mult_207_n773), .CO(DP_mult_207_n770), .S(DP_mult_207_n771) );
  FA_X1 DP_mult_207_U591 ( .A(DP_mult_207_n1294), .B(DP_mult_207_n1206), .CI(
        DP_mult_207_n1272), .CO(DP_mult_207_n768), .S(DP_mult_207_n769) );
  FA_X1 DP_mult_207_U590 ( .A(DP_mult_207_n786), .B(DP_mult_207_n1228), .CI(
        DP_mult_207_n784), .CO(DP_mult_207_n766), .S(DP_mult_207_n767) );
  FA_X1 DP_mult_207_U589 ( .A(DP_mult_207_n771), .B(DP_mult_207_n769), .CI(
        DP_mult_207_n782), .CO(DP_mult_207_n764), .S(DP_mult_207_n765) );
  FA_X1 DP_mult_207_U588 ( .A(DP_mult_207_n767), .B(DP_mult_207_n780), .CI(
        DP_mult_207_n778), .CO(DP_mult_207_n762), .S(DP_mult_207_n763) );
  FA_X1 DP_mult_207_U587 ( .A(DP_mult_207_n776), .B(DP_mult_207_n765), .CI(
        DP_mult_207_n763), .CO(DP_mult_207_n760), .S(DP_mult_207_n761) );
  FA_X1 DP_mult_207_U586 ( .A(DP_mult_207_n772), .B(DP_mult_207_n1205), .CI(
        DP_mult_207_n1227), .CO(DP_mult_207_n758), .S(DP_mult_207_n759) );
  FA_X1 DP_mult_207_U585 ( .A(DP_mult_207_n1249), .B(DP_mult_207_n1293), .CI(
        DP_mult_207_n1315), .CO(DP_mult_207_n756), .S(DP_mult_207_n757) );
  FA_X1 DP_mult_207_U584 ( .A(DP_mult_207_n1338), .B(DP_mult_207_n1271), .CI(
        DP_mult_207_n770), .CO(DP_mult_207_n754), .S(DP_mult_207_n755) );
  FA_X1 DP_mult_207_U583 ( .A(DP_mult_207_n757), .B(DP_mult_207_n768), .CI(
        DP_mult_207_n759), .CO(DP_mult_207_n752), .S(DP_mult_207_n753) );
  FA_X1 DP_mult_207_U582 ( .A(DP_mult_207_n755), .B(DP_mult_207_n766), .CI(
        DP_mult_207_n764), .CO(DP_mult_207_n750), .S(DP_mult_207_n751) );
  FA_X1 DP_mult_207_U581 ( .A(DP_mult_207_n762), .B(DP_mult_207_n753), .CI(
        DP_mult_207_n751), .CO(DP_mult_207_n748), .S(DP_mult_207_n749) );
  FA_X1 DP_mult_207_U579 ( .A(DP_mult_207_n1292), .B(DP_mult_207_n1248), .CI(
        DP_mult_207_n747), .CO(DP_mult_207_n744), .S(DP_mult_207_n745) );
  FA_X1 DP_mult_207_U578 ( .A(DP_mult_207_n1226), .B(DP_mult_207_n1204), .CI(
        DP_mult_207_n1270), .CO(DP_mult_207_n742), .S(DP_mult_207_n743) );
  FA_X1 DP_mult_207_U577 ( .A(DP_mult_207_n756), .B(DP_mult_207_n758), .CI(
        DP_mult_207_n743), .CO(DP_mult_207_n740), .S(DP_mult_207_n741) );
  FA_X1 DP_mult_207_U576 ( .A(DP_mult_207_n754), .B(DP_mult_207_n745), .CI(
        DP_mult_207_n752), .CO(DP_mult_207_n738), .S(DP_mult_207_n739) );
  FA_X1 DP_mult_207_U575 ( .A(DP_mult_207_n750), .B(DP_mult_207_n741), .CI(
        DP_mult_207_n739), .CO(DP_mult_207_n736), .S(DP_mult_207_n737) );
  FA_X1 DP_mult_207_U574 ( .A(DP_mult_207_n746), .B(DP_mult_207_n1203), .CI(
        DP_mult_207_n1247), .CO(DP_mult_207_n734), .S(DP_mult_207_n735) );
  FA_X1 DP_mult_207_U573 ( .A(DP_mult_207_n1225), .B(DP_mult_207_n1291), .CI(
        DP_mult_207_n1269), .CO(DP_mult_207_n732), .S(DP_mult_207_n733) );
  FA_X1 DP_mult_207_U572 ( .A(DP_mult_207_n744), .B(DP_mult_207_n1314), .CI(
        DP_mult_207_n742), .CO(DP_mult_207_n730), .S(DP_mult_207_n731) );
  FA_X1 DP_mult_207_U571 ( .A(DP_mult_207_n735), .B(DP_mult_207_n733), .CI(
        DP_mult_207_n740), .CO(DP_mult_207_n728), .S(DP_mult_207_n729) );
  FA_X1 DP_mult_207_U570 ( .A(DP_mult_207_n738), .B(DP_mult_207_n731), .CI(
        DP_mult_207_n729), .CO(DP_mult_207_n726), .S(DP_mult_207_n727) );
  FA_X1 DP_mult_207_U568 ( .A(DP_mult_207_n1268), .B(DP_mult_207_n1224), .CI(
        DP_mult_207_n725), .CO(DP_mult_207_n722), .S(DP_mult_207_n723) );
  FA_X1 DP_mult_207_U567 ( .A(DP_mult_207_n1202), .B(DP_mult_207_n1246), .CI(
        DP_mult_207_n734), .CO(DP_mult_207_n720), .S(DP_mult_207_n721) );
  FA_X1 DP_mult_207_U566 ( .A(DP_mult_207_n723), .B(DP_mult_207_n732), .CI(
        DP_mult_207_n730), .CO(DP_mult_207_n718), .S(DP_mult_207_n719) );
  FA_X1 DP_mult_207_U565 ( .A(DP_mult_207_n728), .B(DP_mult_207_n721), .CI(
        DP_mult_207_n719), .CO(DP_mult_207_n716), .S(DP_mult_207_n717) );
  FA_X1 DP_mult_207_U564 ( .A(DP_mult_207_n1267), .B(DP_mult_207_n1201), .CI(
        DP_mult_207_n724), .CO(DP_mult_207_n714), .S(DP_mult_207_n715) );
  FA_X1 DP_mult_207_U563 ( .A(DP_mult_207_n1245), .B(DP_mult_207_n1223), .CI(
        DP_mult_207_n1290), .CO(DP_mult_207_n712), .S(DP_mult_207_n713) );
  FA_X1 DP_mult_207_U562 ( .A(DP_mult_207_n715), .B(DP_mult_207_n722), .CI(
        DP_mult_207_n720), .CO(DP_mult_207_n710), .S(DP_mult_207_n711) );
  FA_X1 DP_mult_207_U561 ( .A(DP_mult_207_n718), .B(DP_mult_207_n713), .CI(
        DP_mult_207_n711), .CO(DP_mult_207_n708), .S(DP_mult_207_n709) );
  FA_X1 DP_mult_207_U559 ( .A(DP_mult_207_n1222), .B(DP_mult_207_n1200), .CI(
        DP_mult_207_n707), .CO(DP_mult_207_n704), .S(DP_mult_207_n705) );
  FA_X1 DP_mult_207_U558 ( .A(DP_mult_207_n714), .B(DP_mult_207_n1244), .CI(
        DP_mult_207_n705), .CO(DP_mult_207_n702), .S(DP_mult_207_n703) );
  FA_X1 DP_mult_207_U557 ( .A(DP_mult_207_n710), .B(DP_mult_207_n712), .CI(
        DP_mult_207_n703), .CO(DP_mult_207_n700), .S(DP_mult_207_n701) );
  FA_X1 DP_mult_207_U556 ( .A(DP_mult_207_n1221), .B(DP_mult_207_n1199), .CI(
        DP_mult_207_n706), .CO(DP_mult_207_n698), .S(DP_mult_207_n699) );
  FA_X1 DP_mult_207_U555 ( .A(DP_mult_207_n1266), .B(DP_mult_207_n1243), .CI(
        DP_mult_207_n704), .CO(DP_mult_207_n696), .S(DP_mult_207_n697) );
  FA_X1 DP_mult_207_U554 ( .A(DP_mult_207_n702), .B(DP_mult_207_n699), .CI(
        DP_mult_207_n697), .CO(DP_mult_207_n694), .S(DP_mult_207_n695) );
  FA_X1 DP_mult_207_U552 ( .A(DP_mult_207_n1198), .B(DP_mult_207_n1220), .CI(
        DP_mult_207_n693), .CO(DP_mult_207_n690), .S(DP_mult_207_n691) );
  FA_X1 DP_mult_207_U551 ( .A(DP_mult_207_n691), .B(DP_mult_207_n698), .CI(
        DP_mult_207_n696), .CO(DP_mult_207_n688), .S(DP_mult_207_n689) );
  FA_X1 DP_mult_207_U550 ( .A(DP_mult_207_n1219), .B(DP_mult_207_n692), .CI(
        DP_mult_207_n1197), .CO(DP_mult_207_n686), .S(DP_mult_207_n687) );
  FA_X1 DP_mult_207_U549 ( .A(DP_mult_207_n690), .B(DP_mult_207_n1242), .CI(
        DP_mult_207_n687), .CO(DP_mult_207_n684), .S(DP_mult_207_n685) );
  FA_X1 DP_mult_207_U547 ( .A(DP_mult_207_n683), .B(DP_mult_207_n1196), .CI(
        DP_mult_207_n686), .CO(DP_mult_207_n680), .S(DP_mult_207_n681) );
  FA_X1 DP_mult_207_U546 ( .A(DP_mult_207_n1195), .B(DP_mult_207_n682), .CI(
        DP_mult_207_n1218), .CO(DP_mult_207_n678), .S(DP_mult_207_n679) );
  INV_X2 DP_mult_208_U2757 ( .A(DP_pipe02[0]), .ZN(DP_mult_208_n2270) );
  INV_X1 DP_mult_208_U2756 ( .A(DP_coeffs_ff_int[50]), .ZN(DP_mult_208_n2268)
         );
  INV_X1 DP_mult_208_U2755 ( .A(DP_coeffs_ff_int[50]), .ZN(DP_mult_208_n2267)
         );
  INV_X1 DP_mult_208_U2754 ( .A(DP_mult_208_n2268), .ZN(DP_mult_208_n2266) );
  INV_X1 DP_mult_208_U2753 ( .A(DP_coeffs_ff_int[52]), .ZN(DP_mult_208_n2264)
         );
  INV_X1 DP_mult_208_U2752 ( .A(DP_coeffs_ff_int[52]), .ZN(DP_mult_208_n2263)
         );
  INV_X1 DP_mult_208_U2751 ( .A(DP_coeffs_ff_int[54]), .ZN(DP_mult_208_n2259)
         );
  INV_X1 DP_mult_208_U2750 ( .A(DP_coeffs_ff_int[54]), .ZN(DP_mult_208_n2258)
         );
  INV_X1 DP_mult_208_U2749 ( .A(DP_coeffs_ff_int[56]), .ZN(DP_mult_208_n2254)
         );
  INV_X1 DP_mult_208_U2748 ( .A(DP_coeffs_ff_int[56]), .ZN(DP_mult_208_n2253)
         );
  INV_X1 DP_mult_208_U2747 ( .A(DP_mult_208_n2254), .ZN(DP_mult_208_n2252) );
  INV_X1 DP_mult_208_U2746 ( .A(DP_coeffs_ff_int[58]), .ZN(DP_mult_208_n2248)
         );
  INV_X1 DP_mult_208_U2745 ( .A(DP_mult_208_n2248), .ZN(DP_mult_208_n2247) );
  INV_X1 DP_mult_208_U2744 ( .A(DP_coeffs_ff_int[60]), .ZN(DP_mult_208_n2245)
         );
  INV_X1 DP_mult_208_U2743 ( .A(DP_coeffs_ff_int[60]), .ZN(DP_mult_208_n2244)
         );
  INV_X1 DP_mult_208_U2742 ( .A(DP_mult_208_n2245), .ZN(DP_mult_208_n2243) );
  INV_X1 DP_mult_208_U2741 ( .A(DP_coeffs_ff_int[62]), .ZN(DP_mult_208_n2239)
         );
  INV_X1 DP_mult_208_U2740 ( .A(DP_coeffs_ff_int[62]), .ZN(DP_mult_208_n2238)
         );
  INV_X1 DP_mult_208_U2739 ( .A(DP_mult_208_n2238), .ZN(DP_mult_208_n2237) );
  INV_X1 DP_mult_208_U2738 ( .A(DP_coeffs_ff_int[66]), .ZN(DP_mult_208_n2230)
         );
  INV_X1 DP_mult_208_U2737 ( .A(DP_coeffs_ff_int[66]), .ZN(DP_mult_208_n2229)
         );
  INV_X1 DP_mult_208_U2736 ( .A(DP_mult_208_n2230), .ZN(DP_mult_208_n2228) );
  INV_X1 DP_mult_208_U2735 ( .A(DP_coeffs_ff_int[68]), .ZN(DP_mult_208_n2225)
         );
  INV_X1 DP_mult_208_U2734 ( .A(DP_coeffs_ff_int[68]), .ZN(DP_mult_208_n2224)
         );
  INV_X1 DP_mult_208_U2733 ( .A(DP_mult_208_n2224), .ZN(DP_mult_208_n2223) );
  INV_X1 DP_mult_208_U2732 ( .A(DP_coeffs_ff_int[70]), .ZN(DP_mult_208_n2221)
         );
  INV_X1 DP_mult_208_U2731 ( .A(DP_coeffs_ff_int[70]), .ZN(DP_mult_208_n2220)
         );
  INV_X1 DP_mult_208_U2730 ( .A(DP_mult_208_n2220), .ZN(DP_mult_208_n2219) );
  INV_X1 DP_mult_208_U2729 ( .A(DP_mult_208_n2054), .ZN(DP_mult_208_n2204) );
  INV_X1 DP_mult_208_U2728 ( .A(DP_mult_208_n277), .ZN(DP_mult_208_n2197) );
  INV_X2 DP_mult_208_U2727 ( .A(DP_mult_208_n2268), .ZN(DP_mult_208_n2265) );
  INV_X2 DP_mult_208_U2726 ( .A(DP_mult_208_n2264), .ZN(DP_mult_208_n2261) );
  INV_X2 DP_mult_208_U2725 ( .A(DP_mult_208_n2208), .ZN(DP_mult_208_n2206) );
  INV_X2 DP_mult_208_U2724 ( .A(DP_mult_208_n2097), .ZN(DP_mult_208_n2186) );
  INV_X2 DP_mult_208_U2723 ( .A(DP_mult_208_n2145), .ZN(DP_mult_208_n2180) );
  XNOR2_X1 DP_mult_208_U2722 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1713) );
  XNOR2_X1 DP_mult_208_U2721 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1711) );
  XNOR2_X1 DP_mult_208_U2720 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1719) );
  XNOR2_X1 DP_mult_208_U2719 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1715) );
  XNOR2_X1 DP_mult_208_U2718 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2227), .ZN(
        DP_mult_208_n1709) );
  OAI22_X1 DP_mult_208_U2717 ( .A1(DP_mult_208_n2193), .A2(DP_mult_208_n1683), 
        .B1(DP_mult_208_n1682), .B2(DP_mult_208_n2049), .ZN(DP_mult_208_n836)
         );
  XNOR2_X1 DP_mult_208_U2716 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1717) );
  OAI22_X1 DP_mult_208_U2715 ( .A1(DP_mult_208_n1693), .A2(DP_mult_208_n2193), 
        .B1(DP_mult_208_n1692), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n1396)
         );
  OAI22_X1 DP_mult_208_U2714 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1962), 
        .B1(DP_mult_208_n1706), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n1190)
         );
  OAI22_X1 DP_mult_208_U2713 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1684), 
        .B1(DP_mult_208_n2049), .B2(DP_mult_208_n1683), .ZN(DP_mult_208_n1387)
         );
  INV_X1 DP_mult_208_U2712 ( .A(DP_mult_208_n836), .ZN(DP_mult_208_n837) );
  OAI22_X1 DP_mult_208_U2711 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1688), 
        .B1(DP_mult_208_n2048), .B2(DP_mult_208_n1687), .ZN(DP_mult_208_n1391)
         );
  OAI22_X1 DP_mult_208_U2710 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1685), 
        .B1(DP_mult_208_n1684), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n1388)
         );
  OAI22_X1 DP_mult_208_U2709 ( .A1(DP_mult_208_n2193), .A2(DP_mult_208_n1692), 
        .B1(DP_mult_208_n2048), .B2(DP_mult_208_n1691), .ZN(DP_mult_208_n1395)
         );
  OAI22_X1 DP_mult_208_U2708 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1687), 
        .B1(DP_mult_208_n1686), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n1390)
         );
  OAI22_X1 DP_mult_208_U2707 ( .A1(DP_mult_208_n2193), .A2(DP_mult_208_n1690), 
        .B1(DP_mult_208_n2050), .B2(DP_mult_208_n1689), .ZN(DP_mult_208_n1393)
         );
  OAI22_X1 DP_mult_208_U2706 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1689), 
        .B1(DP_mult_208_n1688), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n1392)
         );
  OAI22_X1 DP_mult_208_U2705 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1686), 
        .B1(DP_mult_208_n2048), .B2(DP_mult_208_n1685), .ZN(DP_mult_208_n1389)
         );
  OAI22_X1 DP_mult_208_U2704 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1691), 
        .B1(DP_mult_208_n1690), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n1394)
         );
  OAI21_X1 DP_mult_208_U2703 ( .B1(DP_mult_208_n2177), .B2(DP_mult_208_n398), 
        .A(DP_mult_208_n399), .ZN(DP_mult_208_n397) );
  OAI21_X1 DP_mult_208_U2702 ( .B1(DP_mult_208_n2177), .B2(DP_mult_208_n389), 
        .A(DP_mult_208_n390), .ZN(DP_mult_208_n388) );
  OAI21_X1 DP_mult_208_U2701 ( .B1(DP_mult_208_n301), .B2(DP_mult_208_n431), 
        .A(DP_mult_208_n432), .ZN(DP_mult_208_n430) );
  OAI21_X1 DP_mult_208_U2700 ( .B1(DP_mult_208_n2178), .B2(DP_mult_208_n411), 
        .A(DP_mult_208_n412), .ZN(DP_mult_208_n410) );
  OAI21_X1 DP_mult_208_U2699 ( .B1(DP_mult_208_n301), .B2(DP_mult_208_n420), 
        .A(DP_mult_208_n421), .ZN(DP_mult_208_n419) );
  OAI21_X1 DP_mult_208_U2698 ( .B1(DP_mult_208_n2177), .B2(DP_mult_208_n343), 
        .A(DP_mult_208_n344), .ZN(DP_mult_208_n342) );
  OAI21_X1 DP_mult_208_U2697 ( .B1(DP_mult_208_n301), .B2(DP_mult_208_n380), 
        .A(DP_mult_208_n381), .ZN(DP_mult_208_n379) );
  OAI21_X1 DP_mult_208_U2696 ( .B1(DP_mult_208_n2178), .B2(DP_mult_208_n371), 
        .A(DP_mult_208_n372), .ZN(DP_mult_208_n370) );
  OAI21_X1 DP_mult_208_U2695 ( .B1(DP_mult_208_n2178), .B2(DP_mult_208_n354), 
        .A(DP_mult_208_n355), .ZN(DP_mult_208_n353) );
  OAI21_X1 DP_mult_208_U2694 ( .B1(DP_mult_208_n301), .B2(DP_mult_208_n438), 
        .A(DP_mult_208_n439), .ZN(DP_mult_208_n437) );
  INV_X1 DP_mult_208_U2693 ( .A(DP_mult_208_n2178), .ZN(DP_mult_208_n448) );
  OAI21_X1 DP_mult_208_U2692 ( .B1(DP_mult_208_n2177), .B2(DP_mult_208_n326), 
        .A(DP_mult_208_n327), .ZN(DP_mult_208_n325) );
  XNOR2_X1 DP_mult_208_U2691 ( .A(DP_mult_208_n437), .B(DP_mult_208_n311), 
        .ZN(DP_pipe0_coeff_pipe02[13]) );
  AOI21_X1 DP_mult_208_U2690 ( .B1(DP_mult_208_n333), .B2(DP_mult_208_n2137), 
        .A(DP_mult_208_n2133), .ZN(DP_mult_208_n327) );
  NAND2_X1 DP_mult_208_U2689 ( .A1(DP_mult_208_n356), .A2(DP_mult_208_n2135), 
        .ZN(DP_mult_208_n347) );
  XNOR2_X1 DP_mult_208_U2688 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2222), .ZN(
        DP_mult_208_n1742) );
  XNOR2_X1 DP_mult_208_U2687 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2223), .ZN(
        DP_mult_208_n1738) );
  XNOR2_X1 DP_mult_208_U2686 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2223), .ZN(
        DP_mult_208_n1744) );
  XNOR2_X1 DP_mult_208_U2685 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2223), .ZN(
        DP_mult_208_n1736) );
  XNOR2_X1 DP_mult_208_U2684 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2223), .ZN(
        DP_mult_208_n1740) );
  OAI22_X1 DP_mult_208_U2683 ( .A1(DP_mult_208_n2017), .A2(DP_mult_208_n1724), 
        .B1(DP_mult_208_n1723), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n1426)
         );
  XNOR2_X1 DP_mult_208_U2682 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2222), .ZN(
        DP_mult_208_n1734) );
  OAI22_X1 DP_mult_208_U2681 ( .A1(DP_mult_208_n2018), .A2(DP_mult_208_n1719), 
        .B1(DP_mult_208_n2212), .B2(DP_mult_208_n1718), .ZN(DP_mult_208_n1421)
         );
  OAI22_X1 DP_mult_208_U2680 ( .A1(DP_mult_208_n2018), .A2(DP_mult_208_n1722), 
        .B1(DP_mult_208_n1721), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n1424)
         );
  OAI22_X1 DP_mult_208_U2679 ( .A1(DP_mult_208_n2017), .A2(DP_mult_208_n1729), 
        .B1(DP_mult_208_n2212), .B2(DP_mult_208_n1728), .ZN(DP_mult_208_n1431)
         );
  OAI22_X1 DP_mult_208_U2678 ( .A1(DP_mult_208_n2194), .A2(DP_mult_208_n1728), 
        .B1(DP_mult_208_n1727), .B2(DP_mult_208_n2213), .ZN(DP_mult_208_n1430)
         );
  OAI22_X1 DP_mult_208_U2677 ( .A1(DP_mult_208_n2017), .A2(DP_mult_208_n1723), 
        .B1(DP_mult_208_n2213), .B2(DP_mult_208_n1722), .ZN(DP_mult_208_n1425)
         );
  OAI22_X1 DP_mult_208_U2676 ( .A1(DP_mult_208_n2018), .A2(DP_mult_208_n1725), 
        .B1(DP_mult_208_n2213), .B2(DP_mult_208_n1724), .ZN(DP_mult_208_n1427)
         );
  OAI22_X1 DP_mult_208_U2675 ( .A1(DP_mult_208_n2017), .A2(DP_mult_208_n1730), 
        .B1(DP_mult_208_n1729), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n1432)
         );
  OAI22_X1 DP_mult_208_U2674 ( .A1(DP_mult_208_n2017), .A2(DP_mult_208_n1726), 
        .B1(DP_mult_208_n1725), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n1428)
         );
  OAI22_X1 DP_mult_208_U2673 ( .A1(DP_mult_208_n2018), .A2(DP_mult_208_n1721), 
        .B1(DP_mult_208_n2213), .B2(DP_mult_208_n1720), .ZN(DP_mult_208_n1423)
         );
  OAI22_X1 DP_mult_208_U2672 ( .A1(DP_mult_208_n2018), .A2(DP_mult_208_n1720), 
        .B1(DP_mult_208_n1719), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n1422)
         );
  OAI22_X1 DP_mult_208_U2671 ( .A1(DP_mult_208_n2194), .A2(DP_mult_208_n1727), 
        .B1(DP_mult_208_n2213), .B2(DP_mult_208_n1726), .ZN(DP_mult_208_n1429)
         );
  OAI21_X1 DP_mult_208_U2670 ( .B1(DP_mult_208_n536), .B2(DP_mult_208_n498), 
        .A(DP_mult_208_n499), .ZN(DP_mult_208_n497) );
  OAI21_X1 DP_mult_208_U2669 ( .B1(DP_mult_208_n536), .B2(DP_mult_208_n2113), 
        .A(DP_mult_208_n2163), .ZN(DP_mult_208_n504) );
  OAI21_X1 DP_mult_208_U2668 ( .B1(DP_mult_208_n536), .B2(DP_mult_208_n516), 
        .A(DP_mult_208_n517), .ZN(DP_mult_208_n515) );
  OAI21_X1 DP_mult_208_U2667 ( .B1(DP_mult_208_n536), .B2(DP_mult_208_n476), 
        .A(DP_mult_208_n477), .ZN(DP_mult_208_n475) );
  OAI21_X1 DP_mult_208_U2666 ( .B1(DP_mult_208_n536), .B2(DP_mult_208_n523), 
        .A(DP_mult_208_n524), .ZN(DP_mult_208_n522) );
  OAI21_X1 DP_mult_208_U2665 ( .B1(DP_mult_208_n536), .B2(DP_mult_208_n463), 
        .A(DP_mult_208_n464), .ZN(DP_mult_208_n462) );
  OAI21_X1 DP_mult_208_U2664 ( .B1(DP_mult_208_n536), .B2(DP_mult_208_n487), 
        .A(DP_mult_208_n488), .ZN(DP_mult_208_n486) );
  OAI21_X1 DP_mult_208_U2663 ( .B1(DP_mult_208_n536), .B2(DP_mult_208_n2058), 
        .A(DP_mult_208_n2111), .ZN(DP_mult_208_n533) );
  XNOR2_X1 DP_mult_208_U2662 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2216), .ZN(
        DP_mult_208_n1769) );
  XNOR2_X1 DP_mult_208_U2661 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2216), .ZN(
        DP_mult_208_n1765) );
  XNOR2_X1 DP_mult_208_U2660 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2216), .ZN(
        DP_mult_208_n1761) );
  XNOR2_X1 DP_mult_208_U2659 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2216), .ZN(
        DP_mult_208_n1767) );
  XNOR2_X1 DP_mult_208_U2658 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2216), .ZN(
        DP_mult_208_n1759) );
  OAI22_X1 DP_mult_208_U2657 ( .A1(DP_mult_208_n2196), .A2(DP_mult_208_n1733), 
        .B1(DP_mult_208_n1732), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n916)
         );
  XNOR2_X1 DP_mult_208_U2656 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2216), .ZN(
        DP_mult_208_n1763) );
  OAI22_X1 DP_mult_208_U2655 ( .A1(DP_mult_208_n2062), .A2(DP_mult_208_n1742), 
        .B1(DP_mult_208_n2011), .B2(DP_mult_208_n1741), .ZN(DP_mult_208_n1443)
         );
  OAI22_X1 DP_mult_208_U2654 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1737), 
        .B1(DP_mult_208_n1736), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n1438)
         );
  OAI22_X1 DP_mult_208_U2653 ( .A1(DP_mult_208_n2062), .A2(DP_mult_208_n1743), 
        .B1(DP_mult_208_n1742), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n1444)
         );
  OAI22_X1 DP_mult_208_U2652 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1734), 
        .B1(DP_mult_208_n2011), .B2(DP_mult_208_n1733), .ZN(DP_mult_208_n1435)
         );
  OAI22_X1 DP_mult_208_U2651 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1739), 
        .B1(DP_mult_208_n1738), .B2(DP_mult_208_n2011), .ZN(DP_mult_208_n1440)
         );
  OAI22_X1 DP_mult_208_U2650 ( .A1(DP_mult_208_n2062), .A2(DP_mult_208_n1735), 
        .B1(DP_mult_208_n1734), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n1436)
         );
  OAI22_X1 DP_mult_208_U2649 ( .A1(DP_mult_208_n2196), .A2(DP_mult_208_n1736), 
        .B1(DP_mult_208_n1937), .B2(DP_mult_208_n1735), .ZN(DP_mult_208_n1437)
         );
  OAI22_X1 DP_mult_208_U2648 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1740), 
        .B1(DP_mult_208_n1937), .B2(DP_mult_208_n1739), .ZN(DP_mult_208_n1441)
         );
  OAI22_X1 DP_mult_208_U2647 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1741), 
        .B1(DP_mult_208_n1740), .B2(DP_mult_208_n2011), .ZN(DP_mult_208_n1442)
         );
  OAI22_X1 DP_mult_208_U2646 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1738), 
        .B1(DP_mult_208_n2011), .B2(DP_mult_208_n1737), .ZN(DP_mult_208_n1439)
         );
  OAI22_X1 DP_mult_208_U2645 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n2225), 
        .B1(DP_mult_208_n1756), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n1192)
         );
  INV_X1 DP_mult_208_U2644 ( .A(DP_mult_208_n2096), .ZN(DP_mult_208_n492) );
  AOI21_X1 DP_mult_208_U2643 ( .B1(DP_mult_208_n508), .B2(DP_mult_208_n2116), 
        .A(DP_mult_208_n2174), .ZN(DP_mult_208_n488) );
  XNOR2_X1 DP_mult_208_U2642 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2240), .ZN(
        DP_mult_208_n1642) );
  XNOR2_X1 DP_mult_208_U2641 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2240), .ZN(
        DP_mult_208_n1640) );
  XNOR2_X1 DP_mult_208_U2640 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2240), .ZN(
        DP_mult_208_n1644) );
  XNOR2_X1 DP_mult_208_U2639 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2240), .ZN(
        DP_mult_208_n1638) );
  OAI22_X1 DP_mult_208_U2638 ( .A1(DP_mult_208_n2108), .A2(DP_mult_208_n1608), 
        .B1(DP_mult_208_n1607), .B2(DP_mult_208_n2003), .ZN(DP_mult_208_n746)
         );
  XNOR2_X1 DP_mult_208_U2637 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2240), .ZN(
        DP_mult_208_n1634) );
  XNOR2_X1 DP_mult_208_U2636 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2240), .ZN(
        DP_mult_208_n1636) );
  OAI22_X1 DP_mult_208_U2635 ( .A1(DP_mult_208_n2188), .A2(DP_mult_208_n1614), 
        .B1(DP_mult_208_n1613), .B2(DP_mult_208_n2003), .ZN(DP_mult_208_n1320)
         );
  OAI22_X1 DP_mult_208_U2634 ( .A1(DP_mult_208_n2189), .A2(DP_mult_208_n1616), 
        .B1(DP_mult_208_n1615), .B2(DP_mult_208_n2003), .ZN(DP_mult_208_n1322)
         );
  OAI22_X1 DP_mult_208_U2633 ( .A1(DP_mult_208_n2109), .A2(DP_mult_208_n1618), 
        .B1(DP_mult_208_n1617), .B2(DP_mult_208_n2209), .ZN(DP_mult_208_n1324)
         );
  OAI22_X1 DP_mult_208_U2632 ( .A1(DP_mult_208_n2109), .A2(DP_mult_208_n1953), 
        .B1(DP_mult_208_n1631), .B2(DP_mult_208_n2003), .ZN(DP_mult_208_n1187)
         );
  OAI22_X1 DP_mult_208_U2631 ( .A1(DP_mult_208_n2188), .A2(DP_mult_208_n1609), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1608), .ZN(DP_mult_208_n1315)
         );
  INV_X1 DP_mult_208_U2630 ( .A(DP_mult_208_n746), .ZN(DP_mult_208_n747) );
  OAI22_X1 DP_mult_208_U2629 ( .A1(DP_mult_208_n2188), .A2(DP_mult_208_n1611), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1610), .ZN(DP_mult_208_n1317)
         );
  OAI22_X1 DP_mult_208_U2628 ( .A1(DP_mult_208_n2109), .A2(DP_mult_208_n1615), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1614), .ZN(DP_mult_208_n1321)
         );
  OAI22_X1 DP_mult_208_U2627 ( .A1(DP_mult_208_n2109), .A2(DP_mult_208_n1617), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1616), .ZN(DP_mult_208_n1323)
         );
  OAI22_X1 DP_mult_208_U2626 ( .A1(DP_mult_208_n2109), .A2(DP_mult_208_n1610), 
        .B1(DP_mult_208_n1609), .B2(DP_mult_208_n2003), .ZN(DP_mult_208_n1316)
         );
  OAI22_X1 DP_mult_208_U2625 ( .A1(DP_mult_208_n2109), .A2(DP_mult_208_n1612), 
        .B1(DP_mult_208_n1611), .B2(DP_mult_208_n2003), .ZN(DP_mult_208_n1318)
         );
  OAI22_X1 DP_mult_208_U2624 ( .A1(DP_mult_208_n2108), .A2(DP_mult_208_n1613), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1612), .ZN(DP_mult_208_n1319)
         );
  NAND2_X1 DP_mult_208_U2623 ( .A1(DP_mult_208_n717), .A2(DP_mult_208_n726), 
        .ZN(DP_mult_208_n418) );
  NOR2_X1 DP_mult_208_U2622 ( .A1(DP_mult_208_n420), .A2(DP_mult_208_n347), 
        .ZN(DP_mult_208_n345) );
  NAND2_X1 DP_mult_208_U2621 ( .A1(DP_mult_208_n345), .A2(DP_mult_208_n2134), 
        .ZN(DP_mult_208_n336) );
  INV_X1 DP_mult_208_U2620 ( .A(DP_mult_208_n345), .ZN(DP_mult_208_n343) );
  XNOR2_X1 DP_mult_208_U2619 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1667) );
  XNOR2_X1 DP_mult_208_U2618 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1659) );
  XNOR2_X1 DP_mult_208_U2617 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1665) );
  XNOR2_X1 DP_mult_208_U2616 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1661) );
  XNOR2_X1 DP_mult_208_U2615 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1663) );
  XNOR2_X1 DP_mult_208_U2614 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1669) );
  OAI22_X1 DP_mult_208_U2613 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n2245), 
        .B1(DP_mult_208_n1656), .B2(DP_mult_208_n2210), .ZN(DP_mult_208_n1188)
         );
  OAI22_X1 DP_mult_208_U2612 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1643), 
        .B1(DP_mult_208_n1642), .B2(DP_mult_208_n2210), .ZN(DP_mult_208_n1348)
         );
  OAI22_X1 DP_mult_208_U2611 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1641), 
        .B1(DP_mult_208_n1640), .B2(DP_mult_208_n2210), .ZN(DP_mult_208_n1346)
         );
  OAI22_X1 DP_mult_208_U2610 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1642), 
        .B1(DP_mult_208_n2210), .B2(DP_mult_208_n1641), .ZN(DP_mult_208_n1347)
         );
  OAI22_X1 DP_mult_208_U2609 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1638), 
        .B1(DP_mult_208_n2210), .B2(DP_mult_208_n1637), .ZN(DP_mult_208_n1343)
         );
  OAI22_X1 DP_mult_208_U2608 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1633), 
        .B1(DP_mult_208_n1632), .B2(DP_mult_208_n2211), .ZN(DP_mult_208_n772)
         );
  OAI22_X1 DP_mult_208_U2607 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1640), 
        .B1(DP_mult_208_n2211), .B2(DP_mult_208_n1639), .ZN(DP_mult_208_n1345)
         );
  OAI22_X1 DP_mult_208_U2606 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1639), 
        .B1(DP_mult_208_n1638), .B2(DP_mult_208_n2211), .ZN(DP_mult_208_n1344)
         );
  OAI22_X1 DP_mult_208_U2605 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1635), 
        .B1(DP_mult_208_n1634), .B2(DP_mult_208_n2210), .ZN(DP_mult_208_n1340)
         );
  OAI22_X1 DP_mult_208_U2604 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1634), 
        .B1(DP_mult_208_n2211), .B2(DP_mult_208_n1633), .ZN(DP_mult_208_n1339)
         );
  OAI22_X1 DP_mult_208_U2603 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1636), 
        .B1(DP_mult_208_n2211), .B2(DP_mult_208_n1635), .ZN(DP_mult_208_n1341)
         );
  OAI22_X1 DP_mult_208_U2602 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1637), 
        .B1(DP_mult_208_n1636), .B2(DP_mult_208_n2210), .ZN(DP_mult_208_n1342)
         );
  OAI21_X1 DP_mult_208_U2601 ( .B1(DP_mult_208_n594), .B2(DP_mult_208_n582), 
        .A(DP_mult_208_n583), .ZN(DP_mult_208_n581) );
  XNOR2_X1 DP_mult_208_U2600 ( .A(DP_mult_208_n430), .B(DP_mult_208_n310), 
        .ZN(DP_pipe0_coeff_pipe02[14]) );
  OAI22_X1 DP_mult_208_U2599 ( .A1(DP_mult_208_n2187), .A2(DP_mult_208_n1605), 
        .B1(DP_mult_208_n1604), .B2(DP_mult_208_n2207), .ZN(DP_mult_208_n1312)
         );
  AOI21_X1 DP_mult_208_U2598 ( .B1(DP_mult_208_n553), .B2(DP_mult_208_n540), 
        .A(DP_mult_208_n541), .ZN(DP_mult_208_n539) );
  NAND2_X1 DP_mult_208_U2597 ( .A1(DP_mult_208_n540), .A2(DP_mult_208_n552), 
        .ZN(DP_mult_208_n538) );
  OAI22_X1 DP_mult_208_U2596 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1499), 
        .B1(DP_mult_208_n1498), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1210)
         );
  OAI22_X1 DP_mult_208_U2595 ( .A1(DP_mult_208_n2179), .A2(DP_mult_208_n1498), 
        .B1(DP_mult_208_n2051), .B2(DP_mult_208_n1497), .ZN(DP_mult_208_n1209)
         );
  OAI22_X1 DP_mult_208_U2594 ( .A1(DP_mult_208_n2179), .A2(DP_mult_208_n1504), 
        .B1(DP_mult_208_n2051), .B2(DP_mult_208_n1503), .ZN(DP_mult_208_n1215)
         );
  OAI22_X1 DP_mult_208_U2593 ( .A1(DP_mult_208_n2179), .A2(DP_mult_208_n1503), 
        .B1(DP_mult_208_n1502), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1214)
         );
  OAI22_X1 DP_mult_208_U2592 ( .A1(DP_mult_208_n2179), .A2(DP_mult_208_n1505), 
        .B1(DP_mult_208_n1504), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1216)
         );
  OAI22_X1 DP_mult_208_U2591 ( .A1(DP_mult_208_n2179), .A2(DP_mult_208_n1500), 
        .B1(DP_mult_208_n2051), .B2(DP_mult_208_n1499), .ZN(DP_mult_208_n1211)
         );
  OAI22_X1 DP_mult_208_U2590 ( .A1(DP_mult_208_n2179), .A2(DP_mult_208_n1501), 
        .B1(DP_mult_208_n1500), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1212)
         );
  OAI22_X1 DP_mult_208_U2589 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1494), 
        .B1(DP_mult_208_n2200), .B2(DP_mult_208_n1493), .ZN(DP_mult_208_n1205)
         );
  OAI22_X1 DP_mult_208_U2588 ( .A1(DP_mult_208_n2179), .A2(DP_mult_208_n1502), 
        .B1(DP_mult_208_n2051), .B2(DP_mult_208_n1501), .ZN(DP_mult_208_n1213)
         );
  OAI22_X1 DP_mult_208_U2587 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1496), 
        .B1(DP_mult_208_n2200), .B2(DP_mult_208_n1495), .ZN(DP_mult_208_n1207)
         );
  OAI22_X1 DP_mult_208_U2586 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1495), 
        .B1(DP_mult_208_n1494), .B2(DP_mult_208_n2051), .ZN(DP_mult_208_n1206)
         );
  OAI22_X1 DP_mult_208_U2585 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1497), 
        .B1(DP_mult_208_n1496), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1208)
         );
  XNOR2_X1 DP_mult_208_U2584 ( .A(DP_mult_208_n419), .B(DP_mult_208_n309), 
        .ZN(DP_pipe0_coeff_pipe02[15]) );
  OAI22_X1 DP_mult_208_U2583 ( .A1(DP_mult_208_n2191), .A2(DP_mult_208_n1659), 
        .B1(DP_mult_208_n2056), .B2(DP_mult_208_n1658), .ZN(DP_mult_208_n1363)
         );
  OAI22_X1 DP_mult_208_U2582 ( .A1(DP_mult_208_n2191), .A2(DP_mult_208_n1666), 
        .B1(DP_mult_208_n1665), .B2(DP_mult_208_n2035), .ZN(DP_mult_208_n1370)
         );
  OAI22_X1 DP_mult_208_U2581 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1658), 
        .B1(DP_mult_208_n1657), .B2(DP_mult_208_n2056), .ZN(DP_mult_208_n802)
         );
  OAI22_X1 DP_mult_208_U2580 ( .A1(DP_mult_208_n2191), .A2(DP_mult_208_n1662), 
        .B1(DP_mult_208_n1661), .B2(DP_mult_208_n2056), .ZN(DP_mult_208_n1366)
         );
  OAI22_X1 DP_mult_208_U2579 ( .A1(DP_mult_208_n2191), .A2(DP_mult_208_n1665), 
        .B1(DP_mult_208_n1958), .B2(DP_mult_208_n1664), .ZN(DP_mult_208_n1369)
         );
  OAI22_X1 DP_mult_208_U2578 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1667), 
        .B1(DP_mult_208_n2056), .B2(DP_mult_208_n1666), .ZN(DP_mult_208_n1371)
         );
  OAI22_X1 DP_mult_208_U2577 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1664), 
        .B1(DP_mult_208_n1663), .B2(DP_mult_208_n1958), .ZN(DP_mult_208_n1368)
         );
  OAI22_X1 DP_mult_208_U2576 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n2238), 
        .B1(DP_mult_208_n1681), .B2(DP_mult_208_n2035), .ZN(DP_mult_208_n1189)
         );
  OAI22_X1 DP_mult_208_U2575 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1663), 
        .B1(DP_mult_208_n2056), .B2(DP_mult_208_n1662), .ZN(DP_mult_208_n1367)
         );
  OAI22_X1 DP_mult_208_U2574 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1660), 
        .B1(DP_mult_208_n1659), .B2(DP_mult_208_n2056), .ZN(DP_mult_208_n1364)
         );
  OAI22_X1 DP_mult_208_U2573 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1661), 
        .B1(DP_mult_208_n2056), .B2(DP_mult_208_n1660), .ZN(DP_mult_208_n1365)
         );
  NOR2_X1 DP_mult_208_U2572 ( .A1(DP_mult_208_n918), .A2(DP_mult_208_n897), 
        .ZN(DP_mult_208_n534) );
  XNOR2_X1 DP_mult_208_U2571 ( .A(DP_mult_208_n410), .B(DP_mult_208_n308), 
        .ZN(DP_pipe0_coeff_pipe02[16]) );
  OAI22_X1 DP_mult_208_U2570 ( .A1(DP_mult_208_n2181), .A2(DP_mult_208_n1966), 
        .B1(DP_mult_208_n2201), .B2(DP_mult_208_n1526), .ZN(DP_mult_208_n1237)
         );
  OAI22_X1 DP_mult_208_U2569 ( .A1(DP_mult_208_n2181), .A2(DP_mult_208_n1526), 
        .B1(DP_mult_208_n1525), .B2(DP_mult_208_n2202), .ZN(DP_mult_208_n1236)
         );
  OAI22_X1 DP_mult_208_U2568 ( .A1(DP_mult_208_n2181), .A2(DP_mult_208_n1524), 
        .B1(DP_mult_208_n1523), .B2(DP_mult_208_n2202), .ZN(DP_mult_208_n1234)
         );
  OAI22_X1 DP_mult_208_U2567 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1523), 
        .B1(DP_mult_208_n2201), .B2(DP_mult_208_n1522), .ZN(DP_mult_208_n1233)
         );
  OAI22_X1 DP_mult_208_U2566 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1529), 
        .B1(DP_mult_208_n2202), .B2(DP_mult_208_n1528), .ZN(DP_mult_208_n1239)
         );
  OAI22_X1 DP_mult_208_U2565 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1525), 
        .B1(DP_mult_208_n2201), .B2(DP_mult_208_n1524), .ZN(DP_mult_208_n1235)
         );
  OR2_X1 DP_mult_208_U2564 ( .A1(DP_mult_208_n1215), .A2(DP_mult_208_n1237), 
        .ZN(DP_mult_208_n938) );
  OAI22_X1 DP_mult_208_U2563 ( .A1(DP_mult_208_n2044), .A2(DP_mult_208_n1520), 
        .B1(DP_mult_208_n1519), .B2(DP_mult_208_n2201), .ZN(DP_mult_208_n1230)
         );
  OAI22_X1 DP_mult_208_U2562 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1519), 
        .B1(DP_mult_208_n2202), .B2(DP_mult_208_n1518), .ZN(DP_mult_208_n1229)
         );
  XNOR2_X1 DP_mult_208_U2561 ( .A(DP_mult_208_n1237), .B(DP_mult_208_n1215), 
        .ZN(DP_mult_208_n939) );
  OAI22_X1 DP_mult_208_U2560 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1521), 
        .B1(DP_mult_208_n2201), .B2(DP_mult_208_n1520), .ZN(DP_mult_208_n1231)
         );
  OAI22_X1 DP_mult_208_U2559 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1522), 
        .B1(DP_mult_208_n1521), .B2(DP_mult_208_n2201), .ZN(DP_mult_208_n1232)
         );
  XNOR2_X1 DP_mult_208_U2558 ( .A(DP_mult_208_n397), .B(DP_mult_208_n307), 
        .ZN(DP_pipe0_coeff_pipe02[17]) );
  XNOR2_X1 DP_mult_208_U2557 ( .A(DP_pipe02[15]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1515) );
  XNOR2_X1 DP_mult_208_U2556 ( .A(DP_pipe02[13]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1517) );
  XNOR2_X1 DP_mult_208_U2555 ( .A(DP_pipe02[19]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1511) );
  XNOR2_X1 DP_mult_208_U2554 ( .A(DP_pipe02[11]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1519) );
  XNOR2_X1 DP_mult_208_U2553 ( .A(DP_pipe02[21]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1509) );
  OAI22_X1 DP_mult_208_U2552 ( .A1(DP_mult_208_n2179), .A2(DP_mult_208_n2269), 
        .B1(DP_mult_208_n1506), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1182)
         );
  OAI22_X1 DP_mult_208_U2551 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1493), 
        .B1(DP_mult_208_n1492), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1204)
         );
  XNOR2_X1 DP_mult_208_U2550 ( .A(DP_pipe02[17]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1513) );
  OAI22_X1 DP_mult_208_U2549 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1489), 
        .B1(DP_mult_208_n1488), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1200)
         );
  OAI22_X1 DP_mult_208_U2548 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1492), 
        .B1(DP_mult_208_n2051), .B2(DP_mult_208_n1491), .ZN(DP_mult_208_n1203)
         );
  OAI22_X1 DP_mult_208_U2547 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1486), 
        .B1(DP_mult_208_n2200), .B2(DP_mult_208_n1485), .ZN(DP_mult_208_n1197)
         );
  OAI22_X1 DP_mult_208_U2546 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1490), 
        .B1(DP_mult_208_n2051), .B2(DP_mult_208_n1489), .ZN(DP_mult_208_n1201)
         );
  OAI22_X1 DP_mult_208_U2545 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1487), 
        .B1(DP_mult_208_n1486), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1198)
         );
  OAI22_X1 DP_mult_208_U2544 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1488), 
        .B1(DP_mult_208_n2051), .B2(DP_mult_208_n1487), .ZN(DP_mult_208_n1199)
         );
  OAI22_X1 DP_mult_208_U2543 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1491), 
        .B1(DP_mult_208_n1490), .B2(DP_mult_208_n2200), .ZN(DP_mult_208_n1202)
         );
  OAI22_X1 DP_mult_208_U2542 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1485), 
        .B1(DP_mult_208_n1484), .B2(DP_mult_208_n2051), .ZN(DP_mult_208_n1196)
         );
  OAI22_X1 DP_mult_208_U2541 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1484), 
        .B1(DP_mult_208_n2051), .B2(DP_mult_208_n1483), .ZN(DP_mult_208_n1195)
         );
  OAI22_X1 DP_mult_208_U2540 ( .A1(DP_mult_208_n2180), .A2(DP_mult_208_n1483), 
        .B1(DP_mult_208_n1482), .B2(DP_mult_208_n2051), .ZN(DP_mult_208_n676)
         );
  XNOR2_X1 DP_mult_208_U2539 ( .A(DP_mult_208_n370), .B(DP_mult_208_n304), 
        .ZN(DP_pipe0_coeff_pipe02[20]) );
  OAI21_X1 DP_mult_208_U2538 ( .B1(DP_mult_208_n2147), .B2(DP_mult_208_n2176), 
        .A(DP_mult_208_n2275), .ZN(DP_mult_208_n1362) );
  XNOR2_X1 DP_mult_208_U2537 ( .A(DP_mult_208_n388), .B(DP_mult_208_n306), 
        .ZN(DP_pipe0_coeff_pipe02[18]) );
  OAI22_X1 DP_mult_208_U2536 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1680), 
        .B1(DP_mult_208_n1679), .B2(DP_mult_208_n2056), .ZN(DP_mult_208_n1384)
         );
  INV_X1 DP_mult_208_U2535 ( .A(DP_mult_208_n531), .ZN(DP_mult_208_n671) );
  XNOR2_X1 DP_mult_208_U2534 ( .A(DP_mult_208_n379), .B(DP_mult_208_n305), 
        .ZN(DP_pipe0_coeff_pipe02[19]) );
  XNOR2_X1 DP_mult_208_U2533 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2249), .ZN(
        DP_mult_208_n1594) );
  XNOR2_X1 DP_mult_208_U2532 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2249), .ZN(
        DP_mult_208_n1590) );
  XNOR2_X1 DP_mult_208_U2531 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2249), .ZN(
        DP_mult_208_n1592) );
  XNOR2_X1 DP_mult_208_U2530 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2249), .ZN(
        DP_mult_208_n1586) );
  XNOR2_X1 DP_mult_208_U2529 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2249), .ZN(
        DP_mult_208_n1588) );
  XNOR2_X1 DP_mult_208_U2528 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2249), .ZN(
        DP_mult_208_n1584) );
  OAI22_X1 DP_mult_208_U2527 ( .A1(DP_mult_208_n2120), .A2(DP_mult_208_n1568), 
        .B1(DP_mult_208_n1567), .B2(DP_mult_208_n2205), .ZN(DP_mult_208_n1276)
         );
  OAI22_X1 DP_mult_208_U2526 ( .A1(DP_mult_208_n2185), .A2(DP_mult_208_n1558), 
        .B1(DP_mult_208_n1557), .B2(DP_mult_208_n2037), .ZN(DP_mult_208_n706)
         );
  OAI22_X1 DP_mult_208_U2525 ( .A1(DP_mult_208_n2185), .A2(DP_mult_208_n1580), 
        .B1(DP_mult_208_n1579), .B2(DP_mult_208_n2205), .ZN(DP_mult_208_n1288)
         );
  OAI22_X1 DP_mult_208_U2524 ( .A1(DP_mult_208_n2184), .A2(DP_mult_208_n1562), 
        .B1(DP_mult_208_n1561), .B2(DP_mult_208_n2205), .ZN(DP_mult_208_n1270)
         );
  OAI22_X1 DP_mult_208_U2523 ( .A1(DP_mult_208_n2185), .A2(DP_mult_208_n1578), 
        .B1(DP_mult_208_n1577), .B2(DP_mult_208_n2205), .ZN(DP_mult_208_n1286)
         );
  OAI22_X1 DP_mult_208_U2522 ( .A1(DP_mult_208_n2185), .A2(DP_mult_208_n1564), 
        .B1(DP_mult_208_n1563), .B2(DP_mult_208_n2205), .ZN(DP_mult_208_n1272)
         );
  OAI22_X1 DP_mult_208_U2521 ( .A1(DP_mult_208_n2184), .A2(DP_mult_208_n2258), 
        .B1(DP_mult_208_n1581), .B2(DP_mult_208_n2037), .ZN(DP_mult_208_n1185)
         );
  OAI22_X1 DP_mult_208_U2520 ( .A1(DP_mult_208_n2120), .A2(DP_mult_208_n1566), 
        .B1(DP_mult_208_n1565), .B2(DP_mult_208_n2205), .ZN(DP_mult_208_n1274)
         );
  OAI22_X1 DP_mult_208_U2519 ( .A1(DP_mult_208_n2120), .A2(DP_mult_208_n1560), 
        .B1(DP_mult_208_n1559), .B2(DP_mult_208_n2012), .ZN(DP_mult_208_n1268)
         );
  NAND2_X1 DP_mult_208_U2518 ( .A1(DP_mult_208_n2131), .A2(DP_mult_208_n2136), 
        .ZN(DP_mult_208_n364) );
  NAND2_X1 DP_mult_208_U2517 ( .A1(DP_mult_208_n422), .A2(DP_mult_208_n356), 
        .ZN(DP_mult_208_n354) );
  AOI21_X1 DP_mult_208_U2516 ( .B1(DP_mult_208_n423), .B2(DP_mult_208_n356), 
        .A(DP_mult_208_n359), .ZN(DP_mult_208_n355) );
  AOI21_X1 DP_mult_208_U2515 ( .B1(DP_mult_208_n383), .B2(DP_mult_208_n2131), 
        .A(DP_mult_208_n376), .ZN(DP_mult_208_n372) );
  NAND2_X1 DP_mult_208_U2514 ( .A1(DP_mult_208_n382), .A2(DP_mult_208_n2131), 
        .ZN(DP_mult_208_n371) );
  NAND2_X1 DP_mult_208_U2513 ( .A1(DP_mult_208_n2131), .A2(DP_mult_208_n378), 
        .ZN(DP_mult_208_n305) );
  INV_X1 DP_mult_208_U2512 ( .A(DP_mult_208_n325), .ZN(
        DP_pipe0_coeff_pipe02[23]) );
  OAI22_X1 DP_mult_208_U2511 ( .A1(DP_mult_208_n2044), .A2(DP_mult_208_n2268), 
        .B1(DP_mult_208_n1531), .B2(DP_mult_208_n2202), .ZN(DP_mult_208_n1183)
         );
  OAI22_X1 DP_mult_208_U2510 ( .A1(DP_mult_208_n2044), .A2(DP_mult_208_n1516), 
        .B1(DP_mult_208_n1515), .B2(DP_mult_208_n2202), .ZN(DP_mult_208_n1226)
         );
  OAI22_X1 DP_mult_208_U2509 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1512), 
        .B1(DP_mult_208_n1511), .B2(DP_mult_208_n2202), .ZN(DP_mult_208_n1222)
         );
  OAI22_X1 DP_mult_208_U2508 ( .A1(DP_mult_208_n2044), .A2(DP_mult_208_n1514), 
        .B1(DP_mult_208_n1513), .B2(DP_mult_208_n2201), .ZN(DP_mult_208_n1224)
         );
  OAI22_X1 DP_mult_208_U2507 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1518), 
        .B1(DP_mult_208_n1517), .B2(DP_mult_208_n2201), .ZN(DP_mult_208_n1228)
         );
  OAI22_X1 DP_mult_208_U2506 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1510), 
        .B1(DP_mult_208_n1509), .B2(DP_mult_208_n2201), .ZN(DP_mult_208_n1220)
         );
  OAI22_X1 DP_mult_208_U2505 ( .A1(DP_mult_208_n2044), .A2(DP_mult_208_n1508), 
        .B1(DP_mult_208_n1507), .B2(DP_mult_208_n2201), .ZN(DP_mult_208_n682)
         );
  XNOR2_X1 DP_mult_208_U2504 ( .A(DP_mult_208_n353), .B(DP_mult_208_n303), 
        .ZN(DP_pipe0_coeff_pipe02[21]) );
  OAI22_X1 DP_mult_208_U2503 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1705), 
        .B1(DP_mult_208_n1704), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n1408)
         );
  OAI22_X1 DP_mult_208_U2502 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1703), 
        .B1(DP_mult_208_n1702), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n1406)
         );
  NAND2_X1 DP_mult_208_U2501 ( .A1(DP_mult_208_n761), .A2(DP_mult_208_n774), 
        .ZN(DP_mult_208_n461) );
  XNOR2_X1 DP_mult_208_U2500 ( .A(DP_mult_208_n342), .B(DP_mult_208_n302), 
        .ZN(DP_pipe0_coeff_pipe02[22]) );
  OAI22_X1 DP_mult_208_U2499 ( .A1(DP_mult_208_n2183), .A2(DP_mult_208_n1551), 
        .B1(DP_mult_208_n1550), .B2(DP_mult_208_n2204), .ZN(DP_mult_208_n1260)
         );
  OAI22_X1 DP_mult_208_U2498 ( .A1(DP_mult_208_n2023), .A2(DP_mult_208_n1547), 
        .B1(DP_mult_208_n1546), .B2(DP_mult_208_n2204), .ZN(DP_mult_208_n1256)
         );
  OAI22_X1 DP_mult_208_U2497 ( .A1(DP_mult_208_n2023), .A2(DP_mult_208_n1548), 
        .B1(DP_mult_208_n2203), .B2(DP_mult_208_n1547), .ZN(DP_mult_208_n1257)
         );
  OAI22_X1 DP_mult_208_U2496 ( .A1(DP_mult_208_n2183), .A2(DP_mult_208_n1554), 
        .B1(DP_mult_208_n2203), .B2(DP_mult_208_n1553), .ZN(DP_mult_208_n1263)
         );
  OAI22_X1 DP_mult_208_U2495 ( .A1(DP_mult_208_n2183), .A2(DP_mult_208_n1545), 
        .B1(DP_mult_208_n1544), .B2(DP_mult_208_n2203), .ZN(DP_mult_208_n1254)
         );
  OAI22_X1 DP_mult_208_U2494 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1546), 
        .B1(DP_mult_208_n2203), .B2(DP_mult_208_n1545), .ZN(DP_mult_208_n1255)
         );
  OAI22_X1 DP_mult_208_U2493 ( .A1(DP_mult_208_n2023), .A2(DP_mult_208_n1550), 
        .B1(DP_mult_208_n2204), .B2(DP_mult_208_n1549), .ZN(DP_mult_208_n1259)
         );
  OAI22_X1 DP_mult_208_U2492 ( .A1(DP_mult_208_n2023), .A2(DP_mult_208_n1549), 
        .B1(DP_mult_208_n1548), .B2(DP_mult_208_n2203), .ZN(DP_mult_208_n1258)
         );
  OAI22_X1 DP_mult_208_U2491 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1555), 
        .B1(DP_mult_208_n1554), .B2(DP_mult_208_n2204), .ZN(DP_mult_208_n1264)
         );
  OAI22_X1 DP_mult_208_U2490 ( .A1(DP_mult_208_n2183), .A2(DP_mult_208_n1552), 
        .B1(DP_mult_208_n2204), .B2(DP_mult_208_n1551), .ZN(DP_mult_208_n1261)
         );
  OAI22_X1 DP_mult_208_U2489 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1544), 
        .B1(DP_mult_208_n2203), .B2(DP_mult_208_n1543), .ZN(DP_mult_208_n1253)
         );
  NOR2_X1 DP_mult_208_U2488 ( .A1(DP_mult_208_n571), .A2(DP_mult_208_n569), 
        .ZN(DP_mult_208_n567) );
  OAI21_X1 DP_mult_208_U2487 ( .B1(DP_mult_208_n572), .B2(DP_mult_208_n1951), 
        .A(DP_mult_208_n570), .ZN(DP_mult_208_n568) );
  OAI22_X1 DP_mult_208_U2486 ( .A1(DP_mult_208_n2187), .A2(DP_mult_208_n1597), 
        .B1(DP_mult_208_n1596), .B2(DP_mult_208_n2206), .ZN(DP_mult_208_n1304)
         );
  OAI22_X1 DP_mult_208_U2485 ( .A1(DP_mult_208_n2187), .A2(DP_mult_208_n1595), 
        .B1(DP_mult_208_n1594), .B2(DP_mult_208_n2206), .ZN(DP_mult_208_n1302)
         );
  OAI22_X1 DP_mult_208_U2484 ( .A1(DP_mult_208_n2187), .A2(DP_mult_208_n1599), 
        .B1(DP_mult_208_n1598), .B2(DP_mult_208_n2206), .ZN(DP_mult_208_n1306)
         );
  OAI22_X1 DP_mult_208_U2483 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1604), 
        .B1(DP_mult_208_n2206), .B2(DP_mult_208_n1603), .ZN(DP_mult_208_n1311)
         );
  OAI22_X1 DP_mult_208_U2482 ( .A1(DP_mult_208_n2187), .A2(DP_mult_208_n2253), 
        .B1(DP_mult_208_n1606), .B2(DP_mult_208_n2206), .ZN(DP_mult_208_n1186)
         );
  OAI22_X1 DP_mult_208_U2481 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1594), 
        .B1(DP_mult_208_n2207), .B2(DP_mult_208_n1593), .ZN(DP_mult_208_n1301)
         );
  OAI22_X1 DP_mult_208_U2480 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1603), 
        .B1(DP_mult_208_n1602), .B2(DP_mult_208_n2207), .ZN(DP_mult_208_n1310)
         );
  OAI22_X1 DP_mult_208_U2479 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1591), 
        .B1(DP_mult_208_n1590), .B2(DP_mult_208_n2206), .ZN(DP_mult_208_n1298)
         );
  OAI22_X1 DP_mult_208_U2478 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1598), 
        .B1(DP_mult_208_n2206), .B2(DP_mult_208_n1597), .ZN(DP_mult_208_n1305)
         );
  OAI22_X1 DP_mult_208_U2477 ( .A1(DP_mult_208_n2047), .A2(DP_mult_208_n1585), 
        .B1(DP_mult_208_n1584), .B2(DP_mult_208_n2207), .ZN(DP_mult_208_n1292)
         );
  OAI22_X1 DP_mult_208_U2476 ( .A1(DP_mult_208_n2187), .A2(DP_mult_208_n1587), 
        .B1(DP_mult_208_n1586), .B2(DP_mult_208_n2207), .ZN(DP_mult_208_n1294)
         );
  OAI22_X1 DP_mult_208_U2475 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1596), 
        .B1(DP_mult_208_n2207), .B2(DP_mult_208_n1595), .ZN(DP_mult_208_n1303)
         );
  OAI22_X1 DP_mult_208_U2474 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1601), 
        .B1(DP_mult_208_n1600), .B2(DP_mult_208_n2206), .ZN(DP_mult_208_n1308)
         );
  OAI22_X1 DP_mult_208_U2473 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1600), 
        .B1(DP_mult_208_n2206), .B2(DP_mult_208_n1599), .ZN(DP_mult_208_n1307)
         );
  OAI22_X1 DP_mult_208_U2472 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1602), 
        .B1(DP_mult_208_n2206), .B2(DP_mult_208_n1601), .ZN(DP_mult_208_n1309)
         );
  OAI22_X1 DP_mult_208_U2471 ( .A1(DP_mult_208_n2047), .A2(DP_mult_208_n1583), 
        .B1(DP_mult_208_n1582), .B2(DP_mult_208_n2207), .ZN(DP_mult_208_n724)
         );
  OAI22_X1 DP_mult_208_U2470 ( .A1(DP_mult_208_n2047), .A2(DP_mult_208_n1589), 
        .B1(DP_mult_208_n1588), .B2(DP_mult_208_n2207), .ZN(DP_mult_208_n1296)
         );
  OAI22_X1 DP_mult_208_U2469 ( .A1(DP_mult_208_n2047), .A2(DP_mult_208_n1593), 
        .B1(DP_mult_208_n1592), .B2(DP_mult_208_n2206), .ZN(DP_mult_208_n1300)
         );
  AOI21_X1 DP_mult_208_U2468 ( .B1(DP_mult_208_n1947), .B2(DP_mult_208_n1971), 
        .A(DP_mult_208_n1987), .ZN(DP_mult_208_n572) );
  OAI22_X1 DP_mult_208_U2467 ( .A1(DP_mult_208_n2191), .A2(DP_mult_208_n1674), 
        .B1(DP_mult_208_n1673), .B2(DP_mult_208_n1958), .ZN(DP_mult_208_n1378)
         );
  NAND2_X1 DP_mult_208_U2466 ( .A1(DP_mult_208_n1816), .A2(DP_mult_208_n2039), 
        .ZN(DP_mult_208_n277) );
  OAI22_X1 DP_mult_208_U2465 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1755), 
        .B1(DP_mult_208_n1754), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n1456)
         );
  INV_X1 DP_mult_208_U2464 ( .A(DP_mult_208_n2036), .ZN(DP_mult_208_n917) );
  OAI22_X1 DP_mult_208_U2463 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1753), 
        .B1(DP_mult_208_n1752), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n1454)
         );
  OAI21_X1 DP_mult_208_U2462 ( .B1(DP_mult_208_n503), .B2(DP_mult_208_n495), 
        .A(DP_mult_208_n496), .ZN(DP_mult_208_n490) );
  NAND2_X1 DP_mult_208_U2461 ( .A1(DP_mult_208_n489), .A2(DP_mult_208_n454), 
        .ZN(DP_mult_208_n452) );
  INV_X1 DP_mult_208_U2460 ( .A(DP_mult_208_n2063), .ZN(DP_mult_208_n667) );
  NAND2_X1 DP_mult_208_U2459 ( .A1(DP_mult_208_n507), .A2(DP_mult_208_n2116), 
        .ZN(DP_mult_208_n487) );
  AOI21_X1 DP_mult_208_U2458 ( .B1(DP_mult_208_n2130), .B2(DP_mult_208_n1975), 
        .A(DP_mult_208_n1986), .ZN(DP_mult_208_n600) );
  NAND2_X1 DP_mult_208_U2457 ( .A1(DP_mult_208_n1071), .A2(DP_mult_208_n1084), 
        .ZN(DP_mult_208_n591) );
  NAND2_X1 DP_mult_208_U2456 ( .A1(DP_mult_208_n2122), .A2(DP_mult_208_n474), 
        .ZN(DP_mult_208_n314) );
  AOI21_X1 DP_mult_208_U2455 ( .B1(DP_mult_208_n2166), .B2(DP_mult_208_n670), 
        .A(DP_mult_208_n519), .ZN(DP_mult_208_n517) );
  INV_X1 DP_mult_208_U2454 ( .A(DP_mult_208_n2166), .ZN(DP_mult_208_n524) );
  AOI21_X1 DP_mult_208_U2453 ( .B1(DP_mult_208_n490), .B2(DP_mult_208_n454), 
        .A(DP_mult_208_n455), .ZN(DP_mult_208_n453) );
  OAI21_X1 DP_mult_208_U2452 ( .B1(DP_mult_208_n506), .B2(DP_mult_208_n452), 
        .A(DP_mult_208_n453), .ZN(DP_mult_208_n451) );
  OAI22_X1 DP_mult_208_U2451 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1539), 
        .B1(DP_mult_208_n1538), .B2(DP_mult_208_n2203), .ZN(DP_mult_208_n1248)
         );
  OAI22_X1 DP_mult_208_U2450 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1541), 
        .B1(DP_mult_208_n1540), .B2(DP_mult_208_n2204), .ZN(DP_mult_208_n1250)
         );
  OAI22_X1 DP_mult_208_U2449 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1533), 
        .B1(DP_mult_208_n1532), .B2(DP_mult_208_n2204), .ZN(DP_mult_208_n692)
         );
  OAI22_X1 DP_mult_208_U2448 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n2264), 
        .B1(DP_mult_208_n1556), .B2(DP_mult_208_n2203), .ZN(DP_mult_208_n1184)
         );
  OAI22_X1 DP_mult_208_U2447 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1543), 
        .B1(DP_mult_208_n1542), .B2(DP_mult_208_n2203), .ZN(DP_mult_208_n1252)
         );
  OAI22_X1 DP_mult_208_U2446 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1537), 
        .B1(DP_mult_208_n1536), .B2(DP_mult_208_n2204), .ZN(DP_mult_208_n1246)
         );
  OAI22_X1 DP_mult_208_U2445 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1535), 
        .B1(DP_mult_208_n1534), .B2(DP_mult_208_n2203), .ZN(DP_mult_208_n1244)
         );
  OAI21_X1 DP_mult_208_U2444 ( .B1(DP_mult_208_n542), .B2(DP_mult_208_n550), 
        .A(DP_mult_208_n543), .ZN(DP_mult_208_n541) );
  NOR2_X1 DP_mult_208_U2443 ( .A1(DP_mult_208_n547), .A2(DP_mult_208_n542), 
        .ZN(DP_mult_208_n540) );
  INV_X1 DP_mult_208_U2442 ( .A(DP_mult_208_n2091), .ZN(DP_mult_208_n565) );
  OAI22_X1 DP_mult_208_U2441 ( .A1(DP_mult_208_n2189), .A2(DP_mult_208_n1628), 
        .B1(DP_mult_208_n1627), .B2(DP_mult_208_n2003), .ZN(DP_mult_208_n1334)
         );
  OAI22_X1 DP_mult_208_U2440 ( .A1(DP_mult_208_n2108), .A2(DP_mult_208_n1630), 
        .B1(DP_mult_208_n1629), .B2(DP_mult_208_n2003), .ZN(DP_mult_208_n1336)
         );
  NAND2_X1 DP_mult_208_U2439 ( .A1(DP_mult_208_n709), .A2(DP_mult_208_n716), 
        .ZN(DP_mult_208_n409) );
  INV_X1 DP_mult_208_U2438 ( .A(DP_mult_208_n346), .ZN(DP_mult_208_n344) );
  OAI22_X1 DP_mult_208_U2437 ( .A1(DP_mult_208_n2195), .A2(DP_mult_208_n1714), 
        .B1(DP_mult_208_n1713), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n1416)
         );
  OAI22_X1 DP_mult_208_U2436 ( .A1(DP_mult_208_n2195), .A2(DP_mult_208_n1712), 
        .B1(DP_mult_208_n1711), .B2(DP_mult_208_n2213), .ZN(DP_mult_208_n1414)
         );
  OAI22_X1 DP_mult_208_U2435 ( .A1(DP_mult_208_n2194), .A2(DP_mult_208_n1708), 
        .B1(DP_mult_208_n1707), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n874)
         );
  OAI22_X1 DP_mult_208_U2434 ( .A1(DP_mult_208_n2195), .A2(DP_mult_208_n1710), 
        .B1(DP_mult_208_n1709), .B2(DP_mult_208_n2213), .ZN(DP_mult_208_n1412)
         );
  OAI22_X1 DP_mult_208_U2433 ( .A1(DP_mult_208_n2194), .A2(DP_mult_208_n1715), 
        .B1(DP_mult_208_n2213), .B2(DP_mult_208_n1714), .ZN(DP_mult_208_n1417)
         );
  OAI22_X1 DP_mult_208_U2432 ( .A1(DP_mult_208_n2018), .A2(DP_mult_208_n1709), 
        .B1(DP_mult_208_n2212), .B2(DP_mult_208_n1708), .ZN(DP_mult_208_n1411)
         );
  OAI22_X1 DP_mult_208_U2431 ( .A1(DP_mult_208_n2017), .A2(DP_mult_208_n1716), 
        .B1(DP_mult_208_n1715), .B2(DP_mult_208_n2213), .ZN(DP_mult_208_n1418)
         );
  OAI22_X1 DP_mult_208_U2430 ( .A1(DP_mult_208_n2194), .A2(DP_mult_208_n1717), 
        .B1(DP_mult_208_n2213), .B2(DP_mult_208_n1716), .ZN(DP_mult_208_n1419)
         );
  OAI22_X1 DP_mult_208_U2429 ( .A1(DP_mult_208_n2017), .A2(DP_mult_208_n1711), 
        .B1(DP_mult_208_n2213), .B2(DP_mult_208_n1710), .ZN(DP_mult_208_n1413)
         );
  OAI22_X1 DP_mult_208_U2428 ( .A1(DP_mult_208_n2018), .A2(DP_mult_208_n1713), 
        .B1(DP_mult_208_n2212), .B2(DP_mult_208_n1712), .ZN(DP_mult_208_n1415)
         );
  OAI22_X1 DP_mult_208_U2427 ( .A1(DP_mult_208_n2194), .A2(DP_mult_208_n1718), 
        .B1(DP_mult_208_n1717), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n1420)
         );
  OAI22_X1 DP_mult_208_U2426 ( .A1(DP_mult_208_n2194), .A2(DP_mult_208_n2229), 
        .B1(DP_mult_208_n1731), .B2(DP_mult_208_n2212), .ZN(DP_mult_208_n1191)
         );
  NOR2_X1 DP_mult_208_U2425 ( .A1(DP_mult_208_n534), .A2(DP_mult_208_n531), 
        .ZN(DP_mult_208_n525) );
  NAND2_X1 DP_mult_208_U2424 ( .A1(DP_mult_208_n511), .A2(DP_mult_208_n525), 
        .ZN(DP_mult_208_n505) );
  INV_X1 DP_mult_208_U2423 ( .A(DP_mult_208_n534), .ZN(DP_mult_208_n672) );
  NAND2_X1 DP_mult_208_U2422 ( .A1(DP_mult_208_n2057), .A2(DP_mult_208_n670), 
        .ZN(DP_mult_208_n516) );
  INV_X1 DP_mult_208_U2421 ( .A(DP_mult_208_n525), .ZN(DP_mult_208_n523) );
  OAI22_X1 DP_mult_208_U2420 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1653), 
        .B1(DP_mult_208_n1652), .B2(DP_mult_208_n2211), .ZN(DP_mult_208_n1358)
         );
  INV_X1 DP_mult_208_U2419 ( .A(DP_mult_208_n772), .ZN(DP_mult_208_n773) );
  OAI22_X1 DP_mult_208_U2418 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1655), 
        .B1(DP_mult_208_n1654), .B2(DP_mult_208_n2210), .ZN(DP_mult_208_n1360)
         );
  NOR2_X1 DP_mult_208_U2417 ( .A1(DP_mult_208_n749), .A2(DP_mult_208_n760), 
        .ZN(DP_mult_208_n438) );
  XNOR2_X1 DP_mult_208_U2416 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2260), .ZN(
        DP_mult_208_n1540) );
  XNOR2_X1 DP_mult_208_U2415 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2261), .ZN(
        DP_mult_208_n1544) );
  XNOR2_X1 DP_mult_208_U2414 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2262), .ZN(
        DP_mult_208_n1538) );
  XNOR2_X1 DP_mult_208_U2413 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2262), .ZN(
        DP_mult_208_n1542) );
  XNOR2_X1 DP_mult_208_U2412 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2260), .ZN(
        DP_mult_208_n1536) );
  XNOR2_X1 DP_mult_208_U2411 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2262), .ZN(
        DP_mult_208_n1534) );
  INV_X1 DP_mult_208_U2410 ( .A(DP_mult_208_n383), .ZN(DP_mult_208_n381) );
  NOR2_X1 DP_mult_208_U2409 ( .A1(DP_mult_208_n1171), .A2(DP_mult_208_n1174), 
        .ZN(DP_mult_208_n633) );
  NAND2_X1 DP_mult_208_U2408 ( .A1(DP_mult_208_n1171), .A2(DP_mult_208_n1174), 
        .ZN(DP_mult_208_n634) );
  OAI22_X1 DP_mult_208_U2407 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1778), 
        .B1(DP_mult_208_n1777), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1479)
         );
  OAI21_X1 DP_mult_208_U2406 ( .B1(DP_mult_208_n628), .B2(DP_mult_208_n626), 
        .A(DP_mult_208_n627), .ZN(DP_mult_208_n625) );
  NOR2_X1 DP_mult_208_U2405 ( .A1(DP_mult_208_n456), .A2(DP_mult_208_n480), 
        .ZN(DP_mult_208_n454) );
  OAI21_X1 DP_mult_208_U2404 ( .B1(DP_mult_208_n456), .B2(DP_mult_208_n481), 
        .A(DP_mult_208_n457), .ZN(DP_mult_208_n455) );
  OAI21_X1 DP_mult_208_U2403 ( .B1(DP_mult_208_n390), .B2(DP_mult_208_n384), 
        .A(DP_mult_208_n387), .ZN(DP_mult_208_n383) );
  XNOR2_X1 DP_mult_208_U2402 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2231), .ZN(
        DP_mult_208_n1692) );
  XNOR2_X1 DP_mult_208_U2401 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2232), .ZN(
        DP_mult_208_n1684) );
  XNOR2_X1 DP_mult_208_U2400 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2233), .ZN(
        DP_mult_208_n1694) );
  XNOR2_X1 DP_mult_208_U2399 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2232), .ZN(
        DP_mult_208_n1686) );
  XNOR2_X1 DP_mult_208_U2398 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2232), .ZN(
        DP_mult_208_n1690) );
  XNOR2_X1 DP_mult_208_U2397 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2232), .ZN(
        DP_mult_208_n1688) );
  OAI22_X1 DP_mult_208_U2396 ( .A1(DP_mult_208_n2108), .A2(DP_mult_208_n1622), 
        .B1(DP_mult_208_n1621), .B2(DP_mult_208_n2209), .ZN(DP_mult_208_n1328)
         );
  OAI22_X1 DP_mult_208_U2395 ( .A1(DP_mult_208_n2108), .A2(DP_mult_208_n1624), 
        .B1(DP_mult_208_n1623), .B2(DP_mult_208_n2209), .ZN(DP_mult_208_n1330)
         );
  OAI22_X1 DP_mult_208_U2394 ( .A1(DP_mult_208_n2188), .A2(DP_mult_208_n1627), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1626), .ZN(DP_mult_208_n1333)
         );
  OAI22_X1 DP_mult_208_U2393 ( .A1(DP_mult_208_n2189), .A2(DP_mult_208_n1619), 
        .B1(DP_mult_208_n2209), .B2(DP_mult_208_n1618), .ZN(DP_mult_208_n1325)
         );
  OAI22_X1 DP_mult_208_U2392 ( .A1(DP_mult_208_n2109), .A2(DP_mult_208_n1623), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1622), .ZN(DP_mult_208_n1329)
         );
  OAI22_X1 DP_mult_208_U2391 ( .A1(DP_mult_208_n2108), .A2(DP_mult_208_n1629), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1628), .ZN(DP_mult_208_n1335)
         );
  OAI22_X1 DP_mult_208_U2390 ( .A1(DP_mult_208_n2188), .A2(DP_mult_208_n1625), 
        .B1(DP_mult_208_n2038), .B2(DP_mult_208_n1624), .ZN(DP_mult_208_n1331)
         );
  OAI22_X1 DP_mult_208_U2389 ( .A1(DP_mult_208_n2188), .A2(DP_mult_208_n1626), 
        .B1(DP_mult_208_n1625), .B2(DP_mult_208_n2038), .ZN(DP_mult_208_n1332)
         );
  OAI22_X1 DP_mult_208_U2388 ( .A1(DP_mult_208_n2108), .A2(DP_mult_208_n1621), 
        .B1(DP_mult_208_n2209), .B2(DP_mult_208_n1620), .ZN(DP_mult_208_n1327)
         );
  OAI22_X1 DP_mult_208_U2387 ( .A1(DP_mult_208_n2188), .A2(DP_mult_208_n1620), 
        .B1(DP_mult_208_n1619), .B2(DP_mult_208_n2038), .ZN(DP_mult_208_n1326)
         );
  OAI22_X1 DP_mult_208_U2386 ( .A1(DP_mult_208_n2187), .A2(DP_mult_208_n1586), 
        .B1(DP_mult_208_n2207), .B2(DP_mult_208_n1585), .ZN(DP_mult_208_n1293)
         );
  OAI22_X1 DP_mult_208_U2385 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1592), 
        .B1(DP_mult_208_n2206), .B2(DP_mult_208_n1591), .ZN(DP_mult_208_n1299)
         );
  OAI22_X1 DP_mult_208_U2384 ( .A1(DP_mult_208_n2186), .A2(DP_mult_208_n1588), 
        .B1(DP_mult_208_n2207), .B2(DP_mult_208_n1587), .ZN(DP_mult_208_n1295)
         );
  OAI22_X1 DP_mult_208_U2383 ( .A1(DP_mult_208_n2047), .A2(DP_mult_208_n1584), 
        .B1(DP_mult_208_n2207), .B2(DP_mult_208_n1583), .ZN(DP_mult_208_n1291)
         );
  OAI22_X1 DP_mult_208_U2382 ( .A1(DP_mult_208_n2047), .A2(DP_mult_208_n1590), 
        .B1(DP_mult_208_n2206), .B2(DP_mult_208_n1589), .ZN(DP_mult_208_n1297)
         );
  NAND2_X1 DP_mult_208_U2381 ( .A1(DP_mult_208_n727), .A2(DP_mult_208_n736), 
        .ZN(DP_mult_208_n429) );
  NOR2_X2 DP_mult_208_U2380 ( .A1(DP_mult_208_n789), .A2(DP_mult_208_n804), 
        .ZN(DP_mult_208_n480) );
  INV_X1 DP_mult_208_U2379 ( .A(DP_mult_208_n480), .ZN(DP_mult_208_n666) );
  OAI21_X1 DP_mult_208_U2378 ( .B1(DP_mult_208_n492), .B2(DP_mult_208_n480), 
        .A(DP_mult_208_n481), .ZN(DP_mult_208_n479) );
  NOR2_X1 DP_mult_208_U2377 ( .A1(DP_mult_208_n491), .A2(DP_mult_208_n480), 
        .ZN(DP_mult_208_n478) );
  XNOR2_X1 DP_mult_208_U2376 ( .A(DP_mult_208_n462), .B(DP_mult_208_n313), 
        .ZN(DP_pipe0_coeff_pipe02[11]) );
  OAI21_X1 DP_mult_208_U2375 ( .B1(DP_mult_208_n2067), .B2(DP_mult_208_n535), 
        .A(DP_mult_208_n532), .ZN(DP_mult_208_n526) );
  NAND2_X1 DP_mult_208_U2374 ( .A1(DP_mult_208_n805), .A2(DP_mult_208_n820), 
        .ZN(DP_mult_208_n496) );
  AOI21_X1 DP_mult_208_U2373 ( .B1(DP_mult_208_n508), .B2(DP_mult_208_n478), 
        .A(DP_mult_208_n479), .ZN(DP_mult_208_n477) );
  NAND2_X1 DP_mult_208_U2372 ( .A1(DP_mult_208_n478), .A2(DP_mult_208_n507), 
        .ZN(DP_mult_208_n476) );
  XNOR2_X1 DP_mult_208_U2371 ( .A(DP_mult_208_n475), .B(DP_mult_208_n314), 
        .ZN(DP_pipe0_coeff_pipe02[10]) );
  OAI21_X1 DP_mult_208_U2370 ( .B1(DP_mult_208_n2197), .B2(DP_mult_208_n2154), 
        .A(DP_mult_208_n2272), .ZN(DP_mult_208_n1434) );
  OAI22_X1 DP_mult_208_U2369 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1540), 
        .B1(DP_mult_208_n2204), .B2(DP_mult_208_n1539), .ZN(DP_mult_208_n1249)
         );
  OAI22_X1 DP_mult_208_U2368 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1538), 
        .B1(DP_mult_208_n2204), .B2(DP_mult_208_n1537), .ZN(DP_mult_208_n1247)
         );
  OAI22_X1 DP_mult_208_U2367 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1542), 
        .B1(DP_mult_208_n2204), .B2(DP_mult_208_n1541), .ZN(DP_mult_208_n1251)
         );
  OAI22_X1 DP_mult_208_U2366 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1534), 
        .B1(DP_mult_208_n2203), .B2(DP_mult_208_n1533), .ZN(DP_mult_208_n1243)
         );
  OAI22_X1 DP_mult_208_U2365 ( .A1(DP_mult_208_n2024), .A2(DP_mult_208_n1536), 
        .B1(DP_mult_208_n2204), .B2(DP_mult_208_n1535), .ZN(DP_mult_208_n1245)
         );
  INV_X1 DP_mult_208_U2364 ( .A(DP_mult_208_n1954), .ZN(DP_mult_208_n675) );
  NAND2_X1 DP_mult_208_U2363 ( .A1(DP_mult_208_n839), .A2(DP_mult_208_n856), 
        .ZN(DP_mult_208_n514) );
  AOI21_X1 DP_mult_208_U2362 ( .B1(DP_mult_208_n589), .B2(DP_mult_208_n2124), 
        .A(DP_mult_208_n1985), .ZN(DP_mult_208_n583) );
  OAI21_X1 DP_mult_208_U2361 ( .B1(DP_mult_208_n590), .B2(DP_mult_208_n593), 
        .A(DP_mult_208_n591), .ZN(DP_mult_208_n589) );
  NOR2_X1 DP_mult_208_U2360 ( .A1(DP_mult_208_n1071), .A2(DP_mult_208_n1084), 
        .ZN(DP_mult_208_n590) );
  OAI22_X1 DP_mult_208_U2359 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1651), 
        .B1(DP_mult_208_n1650), .B2(DP_mult_208_n2210), .ZN(DP_mult_208_n1356)
         );
  OAI22_X1 DP_mult_208_U2358 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1646), 
        .B1(DP_mult_208_n2210), .B2(DP_mult_208_n1645), .ZN(DP_mult_208_n1351)
         );
  OAI22_X1 DP_mult_208_U2357 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1654), 
        .B1(DP_mult_208_n2210), .B2(DP_mult_208_n1653), .ZN(DP_mult_208_n1359)
         );
  OAI22_X1 DP_mult_208_U2356 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1650), 
        .B1(DP_mult_208_n2210), .B2(DP_mult_208_n1649), .ZN(DP_mult_208_n1355)
         );
  OAI22_X1 DP_mult_208_U2355 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1645), 
        .B1(DP_mult_208_n1644), .B2(DP_mult_208_n2211), .ZN(DP_mult_208_n1350)
         );
  OAI22_X1 DP_mult_208_U2354 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1648), 
        .B1(DP_mult_208_n2211), .B2(DP_mult_208_n1647), .ZN(DP_mult_208_n1353)
         );
  OAI22_X1 DP_mult_208_U2353 ( .A1(DP_mult_208_n2079), .A2(DP_mult_208_n1647), 
        .B1(DP_mult_208_n1646), .B2(DP_mult_208_n2211), .ZN(DP_mult_208_n1352)
         );
  OAI22_X1 DP_mult_208_U2352 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1649), 
        .B1(DP_mult_208_n1648), .B2(DP_mult_208_n2211), .ZN(DP_mult_208_n1354)
         );
  OAI22_X1 DP_mult_208_U2351 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1644), 
        .B1(DP_mult_208_n2210), .B2(DP_mult_208_n1643), .ZN(DP_mult_208_n1349)
         );
  OAI22_X1 DP_mult_208_U2350 ( .A1(DP_mult_208_n2089), .A2(DP_mult_208_n1652), 
        .B1(DP_mult_208_n2210), .B2(DP_mult_208_n1651), .ZN(DP_mult_208_n1357)
         );
  AOI21_X1 DP_mult_208_U2349 ( .B1(DP_mult_208_n537), .B2(DP_mult_208_n450), 
        .A(DP_mult_208_n451), .ZN(DP_mult_208_n301) );
  AOI21_X1 DP_mult_208_U2348 ( .B1(DP_mult_208_n537), .B2(DP_mult_208_n450), 
        .A(DP_mult_208_n451), .ZN(DP_mult_208_n2177) );
  AOI21_X1 DP_mult_208_U2347 ( .B1(DP_mult_208_n2114), .B2(DP_mult_208_n450), 
        .A(DP_mult_208_n451), .ZN(DP_mult_208_n2178) );
  INV_X1 DP_mult_208_U2346 ( .A(DP_mult_208_n1934), .ZN(DP_mult_208_n2231) );
  AOI21_X1 DP_mult_208_U2345 ( .B1(DP_mult_208_n629), .B2(DP_mult_208_n635), 
        .A(DP_mult_208_n630), .ZN(DP_mult_208_n628) );
  XNOR2_X1 DP_mult_208_U2344 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2257), .ZN(
        DP_mult_208_n1561) );
  XNOR2_X1 DP_mult_208_U2343 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2256), .ZN(
        DP_mult_208_n1567) );
  XNOR2_X1 DP_mult_208_U2342 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2257), .ZN(
        DP_mult_208_n1563) );
  XNOR2_X1 DP_mult_208_U2341 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2256), .ZN(
        DP_mult_208_n1569) );
  XNOR2_X1 DP_mult_208_U2340 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2257), .ZN(
        DP_mult_208_n1559) );
  XNOR2_X1 DP_mult_208_U2339 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2257), .ZN(
        DP_mult_208_n1565) );
  INV_X1 DP_mult_208_U2338 ( .A(DP_mult_208_n692), .ZN(DP_mult_208_n693) );
  NAND2_X1 DP_mult_208_U2337 ( .A1(DP_mult_208_n362), .A2(DP_mult_208_n2128), 
        .ZN(DP_mult_208_n360) );
  AOI21_X1 DP_mult_208_U2336 ( .B1(DP_mult_208_n362), .B2(DP_mult_208_n394), 
        .A(DP_mult_208_n363), .ZN(DP_mult_208_n361) );
  INV_X1 DP_mult_208_U2335 ( .A(DP_mult_208_n2118), .ZN(DP_mult_208_n508) );
  AOI21_X1 DP_mult_208_U2334 ( .B1(DP_mult_208_n508), .B2(DP_mult_208_n668), 
        .A(DP_mult_208_n501), .ZN(DP_mult_208_n499) );
  AOI21_X1 DP_mult_208_U2333 ( .B1(DP_mult_208_n508), .B2(DP_mult_208_n465), 
        .A(DP_mult_208_n466), .ZN(DP_mult_208_n464) );
  XNOR2_X1 DP_mult_208_U2332 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1609) );
  XNOR2_X1 DP_mult_208_U2331 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1615) );
  XNOR2_X1 DP_mult_208_U2330 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1613) );
  XNOR2_X1 DP_mult_208_U2329 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1619) );
  XNOR2_X1 DP_mult_208_U2328 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1617) );
  XNOR2_X1 DP_mult_208_U2327 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1611) );
  OAI22_X1 DP_mult_208_U2326 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1694), 
        .B1(DP_mult_208_n2049), .B2(DP_mult_208_n1693), .ZN(DP_mult_208_n1397)
         );
  OAI22_X1 DP_mult_208_U2325 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1699), 
        .B1(DP_mult_208_n1698), .B2(DP_mult_208_n2049), .ZN(DP_mult_208_n1402)
         );
  OAI22_X1 DP_mult_208_U2324 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1697), 
        .B1(DP_mult_208_n1696), .B2(DP_mult_208_n2048), .ZN(DP_mult_208_n1400)
         );
  INV_X1 DP_mult_208_U2323 ( .A(DP_mult_208_n706), .ZN(DP_mult_208_n707) );
  OAI21_X1 DP_mult_208_U2322 ( .B1(DP_mult_208_n405), .B2(DP_mult_208_n360), 
        .A(DP_mult_208_n361), .ZN(DP_mult_208_n359) );
  OAI21_X1 DP_mult_208_U2321 ( .B1(DP_mult_208_n337), .B2(DP_mult_208_n334), 
        .A(DP_mult_208_n335), .ZN(DP_mult_208_n333) );
  AOI21_X1 DP_mult_208_U2320 ( .B1(DP_mult_208_n359), .B2(DP_mult_208_n2135), 
        .A(DP_mult_208_n350), .ZN(DP_mult_208_n348) );
  NAND2_X1 DP_mult_208_U2319 ( .A1(DP_mult_208_n2122), .A2(DP_mult_208_n2123), 
        .ZN(DP_mult_208_n456) );
  NAND2_X1 DP_mult_208_U2318 ( .A1(DP_mult_208_n941), .A2(DP_mult_208_n962), 
        .ZN(DP_mult_208_n550) );
  OAI21_X1 DP_mult_208_U2317 ( .B1(DP_mult_208_n428), .B2(DP_mult_208_n436), 
        .A(DP_mult_208_n429), .ZN(DP_mult_208_n427) );
  AOI21_X2 DP_mult_208_U2316 ( .B1(DP_mult_208_n426), .B2(DP_mult_208_n445), 
        .A(DP_mult_208_n427), .ZN(DP_mult_208_n421) );
  AOI21_X1 DP_mult_208_U2315 ( .B1(DP_mult_208_n401), .B2(DP_mult_208_n2128), 
        .A(DP_mult_208_n394), .ZN(DP_mult_208_n390) );
  OAI22_X1 DP_mult_208_U2314 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1700), 
        .B1(DP_mult_208_n2049), .B2(DP_mult_208_n1699), .ZN(DP_mult_208_n1403)
         );
  OAI22_X1 DP_mult_208_U2313 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1696), 
        .B1(DP_mult_208_n2048), .B2(DP_mult_208_n1695), .ZN(DP_mult_208_n1399)
         );
  OAI22_X1 DP_mult_208_U2312 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1704), 
        .B1(DP_mult_208_n2049), .B2(DP_mult_208_n1703), .ZN(DP_mult_208_n1407)
         );
  OAI22_X1 DP_mult_208_U2311 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1695), 
        .B1(DP_mult_208_n1694), .B2(DP_mult_208_n2049), .ZN(DP_mult_208_n1398)
         );
  OAI22_X1 DP_mult_208_U2310 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1702), 
        .B1(DP_mult_208_n2048), .B2(DP_mult_208_n1701), .ZN(DP_mult_208_n1405)
         );
  OAI22_X1 DP_mult_208_U2309 ( .A1(DP_mult_208_n2077), .A2(DP_mult_208_n1698), 
        .B1(DP_mult_208_n2048), .B2(DP_mult_208_n1697), .ZN(DP_mult_208_n1401)
         );
  OAI22_X1 DP_mult_208_U2308 ( .A1(DP_mult_208_n2192), .A2(DP_mult_208_n1701), 
        .B1(DP_mult_208_n1700), .B2(DP_mult_208_n2049), .ZN(DP_mult_208_n1404)
         );
  AOI21_X1 DP_mult_208_U2307 ( .B1(DP_mult_208_n2123), .B2(DP_mult_208_n2061), 
        .A(DP_mult_208_n459), .ZN(DP_mult_208_n457) );
  AOI21_X1 DP_mult_208_U2306 ( .B1(DP_mult_208_n2122), .B2(DP_mult_208_n483), 
        .A(DP_mult_208_n2061), .ZN(DP_mult_208_n468) );
  OAI22_X1 DP_mult_208_U2305 ( .A1(DP_mult_208_n2119), .A2(DP_mult_208_n1576), 
        .B1(DP_mult_208_n1575), .B2(DP_mult_208_n2012), .ZN(DP_mult_208_n1284)
         );
  OAI22_X1 DP_mult_208_U2304 ( .A1(DP_mult_208_n2119), .A2(DP_mult_208_n1574), 
        .B1(DP_mult_208_n1573), .B2(DP_mult_208_n2012), .ZN(DP_mult_208_n1282)
         );
  OAI22_X1 DP_mult_208_U2303 ( .A1(DP_mult_208_n2119), .A2(DP_mult_208_n1572), 
        .B1(DP_mult_208_n1571), .B2(DP_mult_208_n2205), .ZN(DP_mult_208_n1280)
         );
  OAI22_X1 DP_mult_208_U2302 ( .A1(DP_mult_208_n2120), .A2(DP_mult_208_n1577), 
        .B1(DP_mult_208_n2012), .B2(DP_mult_208_n1576), .ZN(DP_mult_208_n1285)
         );
  OAI22_X1 DP_mult_208_U2301 ( .A1(DP_mult_208_n2185), .A2(DP_mult_208_n1579), 
        .B1(DP_mult_208_n2205), .B2(DP_mult_208_n1578), .ZN(DP_mult_208_n1287)
         );
  OAI22_X1 DP_mult_208_U2300 ( .A1(DP_mult_208_n2184), .A2(DP_mult_208_n1573), 
        .B1(DP_mult_208_n2012), .B2(DP_mult_208_n1572), .ZN(DP_mult_208_n1281)
         );
  OAI22_X1 DP_mult_208_U2299 ( .A1(DP_mult_208_n2119), .A2(DP_mult_208_n1569), 
        .B1(DP_mult_208_n2205), .B2(DP_mult_208_n1568), .ZN(DP_mult_208_n1277)
         );
  OAI22_X1 DP_mult_208_U2298 ( .A1(DP_mult_208_n2185), .A2(DP_mult_208_n1575), 
        .B1(DP_mult_208_n2205), .B2(DP_mult_208_n1574), .ZN(DP_mult_208_n1283)
         );
  OAI22_X1 DP_mult_208_U2297 ( .A1(DP_mult_208_n2185), .A2(DP_mult_208_n1571), 
        .B1(DP_mult_208_n2205), .B2(DP_mult_208_n1570), .ZN(DP_mult_208_n1279)
         );
  OAI22_X1 DP_mult_208_U2296 ( .A1(DP_mult_208_n2120), .A2(DP_mult_208_n1570), 
        .B1(DP_mult_208_n1569), .B2(DP_mult_208_n2012), .ZN(DP_mult_208_n1278)
         );
  OAI22_X1 DP_mult_208_U2295 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1751), 
        .B1(DP_mult_208_n1750), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n1452)
         );
  INV_X1 DP_mult_208_U2294 ( .A(DP_mult_208_n2197), .ZN(DP_mult_208_n2196) );
  XNOR2_X1 DP_mult_208_U2293 ( .A(DP_mult_208_n533), .B(DP_mult_208_n320), 
        .ZN(DP_pipe0_coeff_pipe02[4]) );
  XNOR2_X1 DP_mult_208_U2292 ( .A(DP_mult_208_n504), .B(DP_mult_208_n317), 
        .ZN(DP_pipe0_coeff_pipe02[7]) );
  XNOR2_X1 DP_mult_208_U2291 ( .A(DP_mult_208_n522), .B(DP_mult_208_n319), 
        .ZN(DP_pipe0_coeff_pipe02[5]) );
  XNOR2_X1 DP_mult_208_U2290 ( .A(DP_mult_208_n497), .B(DP_mult_208_n316), 
        .ZN(DP_pipe0_coeff_pipe02[8]) );
  XNOR2_X1 DP_mult_208_U2289 ( .A(DP_mult_208_n486), .B(DP_mult_208_n315), 
        .ZN(DP_pipe0_coeff_pipe02[9]) );
  XNOR2_X1 DP_mult_208_U2288 ( .A(DP_mult_208_n515), .B(DP_mult_208_n318), 
        .ZN(DP_pipe0_coeff_pipe02[6]) );
  AOI21_X1 DP_mult_208_U2287 ( .B1(DP_mult_208_n423), .B2(DP_mult_208_n2127), 
        .A(DP_mult_208_n416), .ZN(DP_mult_208_n412) );
  NAND2_X1 DP_mult_208_U2286 ( .A1(DP_mult_208_n422), .A2(DP_mult_208_n2127), 
        .ZN(DP_mult_208_n411) );
  NAND2_X1 DP_mult_208_U2285 ( .A1(DP_mult_208_n332), .A2(DP_mult_208_n2137), 
        .ZN(DP_mult_208_n326) );
  NAND2_X1 DP_mult_208_U2284 ( .A1(DP_mult_208_n2127), .A2(DP_mult_208_n418), 
        .ZN(DP_mult_208_n309) );
  OAI21_X1 DP_mult_208_U2283 ( .B1(DP_mult_208_n2140), .B2(DP_mult_208_n1994), 
        .A(DP_mult_208_n2276), .ZN(DP_mult_208_n1338) );
  INV_X1 DP_mult_208_U2282 ( .A(DP_mult_208_n435), .ZN(DP_mult_208_n662) );
  CLKBUF_X1 DP_mult_208_U2281 ( .A(DP_mult_208_n2096), .Z(DP_mult_208_n2174)
         );
  NAND3_X1 DP_mult_208_U2280 ( .A1(DP_mult_208_n2171), .A2(DP_mult_208_n2172), 
        .A3(DP_mult_208_n2173), .ZN(DP_mult_208_n820) );
  NAND2_X1 DP_mult_208_U2279 ( .A1(DP_mult_208_n825), .A2(DP_mult_208_n823), 
        .ZN(DP_mult_208_n2173) );
  NAND2_X1 DP_mult_208_U2278 ( .A1(DP_mult_208_n840), .A2(DP_mult_208_n823), 
        .ZN(DP_mult_208_n2172) );
  NAND2_X1 DP_mult_208_U2277 ( .A1(DP_mult_208_n840), .A2(DP_mult_208_n825), 
        .ZN(DP_mult_208_n2171) );
  NAND3_X1 DP_mult_208_U2276 ( .A1(DP_mult_208_n2168), .A2(DP_mult_208_n2169), 
        .A3(DP_mult_208_n2170), .ZN(DP_mult_208_n822) );
  NAND2_X1 DP_mult_208_U2275 ( .A1(DP_mult_208_n844), .A2(DP_mult_208_n842), 
        .ZN(DP_mult_208_n2170) );
  NAND2_X1 DP_mult_208_U2274 ( .A1(DP_mult_208_n827), .A2(DP_mult_208_n842), 
        .ZN(DP_mult_208_n2169) );
  NAND2_X1 DP_mult_208_U2273 ( .A1(DP_mult_208_n827), .A2(DP_mult_208_n844), 
        .ZN(DP_mult_208_n2168) );
  XOR2_X1 DP_mult_208_U2272 ( .A(DP_mult_208_n2167), .B(DP_mult_208_n2115), 
        .Z(DP_mult_208_n823) );
  NOR2_X1 DP_mult_208_U2271 ( .A1(DP_mult_208_n520), .A2(DP_mult_208_n513), 
        .ZN(DP_mult_208_n511) );
  NOR2_X1 DP_mult_208_U2270 ( .A1(DP_mult_208_n857), .A2(DP_mult_208_n876), 
        .ZN(DP_mult_208_n520) );
  XNOR2_X1 DP_mult_208_U2269 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2217), .ZN(
        DP_mult_208_n1771) );
  XNOR2_X1 DP_mult_208_U2268 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2217), .ZN(
        DP_mult_208_n1773) );
  XNOR2_X1 DP_mult_208_U2267 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2217), .ZN(
        DP_mult_208_n1757) );
  XNOR2_X1 DP_mult_208_U2266 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2217), .ZN(
        DP_mult_208_n1777) );
  XNOR2_X1 DP_mult_208_U2265 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2217), .ZN(
        DP_mult_208_n1775) );
  OAI22_X1 DP_mult_208_U2264 ( .A1(DP_mult_208_n1946), .A2(DP_mult_208_n1766), 
        .B1(DP_mult_208_n1765), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1467)
         );
  OAI22_X1 DP_mult_208_U2263 ( .A1(DP_mult_208_n2199), .A2(DP_mult_208_n1762), 
        .B1(DP_mult_208_n1761), .B2(DP_mult_208_n2215), .ZN(DP_mult_208_n1463)
         );
  XNOR2_X1 DP_mult_208_U2262 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2217), .ZN(
        DP_mult_208_n1779) );
  OAI22_X1 DP_mult_208_U2261 ( .A1(DP_mult_208_n2199), .A2(DP_mult_208_n1758), 
        .B1(DP_mult_208_n1757), .B2(DP_mult_208_n2215), .ZN(DP_mult_208_n1459)
         );
  OAI22_X1 DP_mult_208_U2260 ( .A1(DP_mult_208_n2059), .A2(DP_mult_208_n1765), 
        .B1(DP_mult_208_n1764), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1466)
         );
  OAI22_X1 DP_mult_208_U2259 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1763), 
        .B1(DP_mult_208_n1762), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1464)
         );
  OAI22_X1 DP_mult_208_U2258 ( .A1(DP_mult_208_n1946), .A2(DP_mult_208_n1761), 
        .B1(DP_mult_208_n1760), .B2(DP_mult_208_n2215), .ZN(DP_mult_208_n1462)
         );
  OAI22_X1 DP_mult_208_U2257 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1764), 
        .B1(DP_mult_208_n1763), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1465)
         );
  OAI22_X1 DP_mult_208_U2256 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1760), 
        .B1(DP_mult_208_n1759), .B2(DP_mult_208_n2215), .ZN(DP_mult_208_n1461)
         );
  OAI22_X1 DP_mult_208_U2255 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1767), 
        .B1(DP_mult_208_n1766), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1468)
         );
  OAI22_X1 DP_mult_208_U2254 ( .A1(DP_mult_208_n2059), .A2(DP_mult_208_n1768), 
        .B1(DP_mult_208_n1767), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1469)
         );
  OAI22_X1 DP_mult_208_U2253 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1759), 
        .B1(DP_mult_208_n1758), .B2(DP_mult_208_n2215), .ZN(DP_mult_208_n1460)
         );
  OAI22_X1 DP_mult_208_U2252 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n2221), 
        .B1(DP_mult_208_n1781), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1193)
         );
  XNOR2_X1 DP_mult_208_U2251 ( .A(DP_pipe02[3]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1527) );
  XNOR2_X1 DP_mult_208_U2250 ( .A(DP_mult_208_n2266), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1528) );
  OAI21_X1 DP_mult_208_U2249 ( .B1(DP_mult_208_n535), .B2(DP_mult_208_n2067), 
        .A(DP_mult_208_n532), .ZN(DP_mult_208_n2166) );
  NAND2_X1 DP_mult_208_U2248 ( .A1(DP_mult_208_n2164), .A2(DP_mult_208_n2165), 
        .ZN(DP_mult_208_n1238) );
  OR2_X1 DP_mult_208_U2247 ( .A1(DP_mult_208_n1527), .A2(DP_mult_208_n2202), 
        .ZN(DP_mult_208_n2165) );
  OR2_X1 DP_mult_208_U2246 ( .A1(DP_mult_208_n2181), .A2(DP_mult_208_n1528), 
        .ZN(DP_mult_208_n2164) );
  INV_X1 DP_mult_208_U2245 ( .A(DP_mult_208_n508), .ZN(DP_mult_208_n2163) );
  NAND3_X1 DP_mult_208_U2244 ( .A1(DP_mult_208_n2161), .A2(DP_mult_208_n2160), 
        .A3(DP_mult_208_n2162), .ZN(DP_mult_208_n952) );
  NAND2_X1 DP_mult_208_U2243 ( .A1(DP_mult_208_n1326), .A2(DP_mult_208_n1392), 
        .ZN(DP_mult_208_n2162) );
  NAND2_X1 DP_mult_208_U2242 ( .A1(DP_mult_208_n961), .A2(DP_mult_208_n1392), 
        .ZN(DP_mult_208_n2161) );
  NAND2_X1 DP_mult_208_U2241 ( .A1(DP_mult_208_n961), .A2(DP_mult_208_n1326), 
        .ZN(DP_mult_208_n2160) );
  OAI21_X1 DP_mult_208_U2240 ( .B1(DP_mult_208_n2090), .B2(DP_mult_208_n538), 
        .A(DP_mult_208_n539), .ZN(DP_mult_208_n537) );
  INV_X1 DP_mult_208_U2239 ( .A(DP_mult_208_n489), .ZN(DP_mult_208_n491) );
  NAND3_X1 DP_mult_208_U2238 ( .A1(DP_mult_208_n2156), .A2(DP_mult_208_n2157), 
        .A3(DP_mult_208_n2158), .ZN(DP_mult_208_n842) );
  NAND2_X1 DP_mult_208_U2237 ( .A1(DP_mult_208_n849), .A2(DP_mult_208_n864), 
        .ZN(DP_mult_208_n2158) );
  NAND2_X1 DP_mult_208_U2236 ( .A1(DP_mult_208_n862), .A2(DP_mult_208_n864), 
        .ZN(DP_mult_208_n2157) );
  NAND2_X1 DP_mult_208_U2235 ( .A1(DP_mult_208_n1957), .A2(DP_mult_208_n849), 
        .ZN(DP_mult_208_n2156) );
  XOR2_X1 DP_mult_208_U2234 ( .A(DP_mult_208_n862), .B(DP_mult_208_n2155), .Z(
        DP_mult_208_n843) );
  XOR2_X1 DP_mult_208_U2233 ( .A(DP_mult_208_n849), .B(DP_mult_208_n864), .Z(
        DP_mult_208_n2155) );
  INV_X1 DP_mult_208_U2232 ( .A(DP_mult_208_n2220), .ZN(DP_mult_208_n2216) );
  XNOR2_X1 DP_mult_208_U2231 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1657) );
  XNOR2_X1 DP_mult_208_U2230 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1673) );
  XNOR2_X1 DP_mult_208_U2229 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1675) );
  XNOR2_X1 DP_mult_208_U2228 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1679) );
  XNOR2_X1 DP_mult_208_U2227 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1671) );
  XNOR2_X1 DP_mult_208_U2226 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2235), .ZN(
        DP_mult_208_n1677) );
  XNOR2_X1 DP_mult_208_U2225 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2262), .ZN(
        DP_mult_208_n1552) );
  XNOR2_X1 DP_mult_208_U2224 ( .A(DP_mult_208_n2261), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1553) );
  NAND2_X1 DP_mult_208_U2223 ( .A1(DP_mult_208_n2152), .A2(DP_mult_208_n2153), 
        .ZN(DP_mult_208_n1262) );
  OR2_X1 DP_mult_208_U2222 ( .A1(DP_mult_208_n1552), .A2(DP_mult_208_n2204), 
        .ZN(DP_mult_208_n2153) );
  OR2_X1 DP_mult_208_U2221 ( .A1(DP_mult_208_n2183), .A2(DP_mult_208_n1553), 
        .ZN(DP_mult_208_n2152) );
  NAND3_X1 DP_mult_208_U2220 ( .A1(DP_mult_208_n2149), .A2(DP_mult_208_n2150), 
        .A3(DP_mult_208_n2151), .ZN(DP_mult_208_n974) );
  NAND2_X1 DP_mult_208_U2219 ( .A1(DP_mult_208_n1415), .A2(DP_mult_208_n1393), 
        .ZN(DP_mult_208_n2151) );
  NAND2_X1 DP_mult_208_U2218 ( .A1(DP_mult_208_n1979), .A2(DP_mult_208_n1393), 
        .ZN(DP_mult_208_n2150) );
  NAND2_X1 DP_mult_208_U2217 ( .A1(DP_mult_208_n1979), .A2(DP_mult_208_n1415), 
        .ZN(DP_mult_208_n2149) );
  INV_X1 DP_mult_208_U2216 ( .A(DP_mult_208_n2245), .ZN(DP_mult_208_n2240) );
  OAI21_X1 DP_mult_208_U2215 ( .B1(DP_mult_208_n1977), .B2(DP_mult_208_n2139), 
        .A(DP_mult_208_n2273), .ZN(DP_mult_208_n1410) );
  INV_X1 DP_mult_208_U2214 ( .A(DP_mult_208_n382), .ZN(DP_mult_208_n380) );
  OAI21_X1 DP_mult_208_U2213 ( .B1(DP_mult_208_n2098), .B2(DP_mult_208_n2208), 
        .A(DP_mult_208_n2278), .ZN(DP_mult_208_n1290) );
  XNOR2_X1 DP_mult_208_U2212 ( .A(DP_mult_208_n2252), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1605) );
  XNOR2_X1 DP_mult_208_U2211 ( .A(DP_mult_208_n2223), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1755) );
  XNOR2_X1 DP_mult_208_U2210 ( .A(DP_mult_208_n2236), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1680) );
  XNOR2_X1 DP_mult_208_U2209 ( .A(DP_mult_208_n2260), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1555) );
  XNOR2_X1 DP_mult_208_U2208 ( .A(DP_mult_208_n2247), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1630) );
  XNOR2_X1 DP_mult_208_U2207 ( .A(DP_mult_208_n2243), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1655) );
  XNOR2_X1 DP_mult_208_U2206 ( .A(DP_mult_208_n2265), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1530) );
  XNOR2_X1 DP_mult_208_U2205 ( .A(DP_mult_208_n2020), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1505) );
  XNOR2_X1 DP_mult_208_U2204 ( .A(DP_mult_208_n2233), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1705) );
  XNOR2_X1 DP_mult_208_U2203 ( .A(DP_mult_208_n2257), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1580) );
  XNOR2_X1 DP_mult_208_U2202 ( .A(DP_mult_208_n2228), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1730) );
  XNOR2_X1 DP_mult_208_U2201 ( .A(DP_mult_208_n2219), .B(DP_pipe02[0]), .ZN(
        DP_mult_208_n1780) );
  INV_X1 DP_mult_208_U2200 ( .A(DP_mult_208_n2259), .ZN(DP_mult_208_n2256) );
  NAND2_X1 DP_mult_208_U2199 ( .A1(DP_mult_208_n897), .A2(DP_mult_208_n918), 
        .ZN(DP_mult_208_n535) );
  NOR2_X1 DP_mult_208_U2198 ( .A1(DP_mult_208_n554), .A2(DP_mult_208_n1949), 
        .ZN(DP_mult_208_n545) );
  OAI21_X1 DP_mult_208_U2197 ( .B1(DP_mult_208_n555), .B2(DP_mult_208_n1949), 
        .A(DP_mult_208_n1948), .ZN(DP_mult_208_n546) );
  INV_X1 DP_mult_208_U2196 ( .A(DP_mult_208_n1949), .ZN(DP_mult_208_n674) );
  OAI21_X1 DP_mult_208_U2195 ( .B1(DP_mult_208_n2142), .B2(DP_mult_208_n2117), 
        .A(DP_mult_208_n2279), .ZN(DP_mult_208_n1266) );
  OAI22_X1 DP_mult_208_U2194 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1517), 
        .B1(DP_mult_208_n2202), .B2(DP_mult_208_n1516), .ZN(DP_mult_208_n1227)
         );
  OAI22_X1 DP_mult_208_U2193 ( .A1(DP_mult_208_n2044), .A2(DP_mult_208_n1515), 
        .B1(DP_mult_208_n2202), .B2(DP_mult_208_n1514), .ZN(DP_mult_208_n1225)
         );
  OAI22_X1 DP_mult_208_U2192 ( .A1(DP_mult_208_n2044), .A2(DP_mult_208_n1509), 
        .B1(DP_mult_208_n2202), .B2(DP_mult_208_n1508), .ZN(DP_mult_208_n1219)
         );
  OAI22_X1 DP_mult_208_U2191 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1511), 
        .B1(DP_mult_208_n2201), .B2(DP_mult_208_n1510), .ZN(DP_mult_208_n1221)
         );
  OAI22_X1 DP_mult_208_U2190 ( .A1(DP_mult_208_n2044), .A2(DP_mult_208_n1513), 
        .B1(DP_mult_208_n2202), .B2(DP_mult_208_n1512), .ZN(DP_mult_208_n1223)
         );
  INV_X1 DP_mult_208_U2189 ( .A(DP_mult_208_n265), .ZN(DP_mult_208_n2208) );
  INV_X1 DP_mult_208_U2188 ( .A(DP_mult_208_n2015), .ZN(DP_mult_208_n670) );
  XNOR2_X1 DP_mult_208_U2187 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1482) );
  XNOR2_X1 DP_mult_208_U2186 ( .A(DP_mult_208_n448), .B(DP_mult_208_n312), 
        .ZN(DP_pipe0_coeff_pipe02[12]) );
  AOI21_X1 DP_mult_208_U2185 ( .B1(DP_mult_208_n565), .B2(DP_mult_208_n545), 
        .A(DP_mult_208_n546), .ZN(DP_mult_208_n544) );
  AOI21_X1 DP_mult_208_U2184 ( .B1(DP_mult_208_n565), .B2(DP_mult_208_n561), 
        .A(DP_mult_208_n562), .ZN(DP_mult_208_n560) );
  NAND2_X1 DP_mult_208_U2183 ( .A1(DP_mult_208_n667), .A2(DP_mult_208_n496), 
        .ZN(DP_mult_208_n316) );
  NAND2_X1 DP_mult_208_U2182 ( .A1(DP_mult_208_n2123), .A2(DP_mult_208_n461), 
        .ZN(DP_mult_208_n313) );
  INV_X1 DP_mult_208_U2181 ( .A(DP_coeffs_ff_int[71]), .ZN(DP_mult_208_n251)
         );
  AND2_X2 DP_mult_208_U2180 ( .A1(DP_mult_208_n1807), .A2(DP_mult_208_n1935), 
        .ZN(DP_mult_208_n2144) );
  INV_X1 DP_mult_208_U2179 ( .A(DP_mult_208_n1757), .ZN(DP_mult_208_n2271) );
  OAI21_X1 DP_mult_208_U2178 ( .B1(DP_coeffs_ff_int[71]), .B2(
        DP_mult_208_n2052), .A(DP_mult_208_n2271), .ZN(DP_mult_208_n1458) );
  NAND2_X1 DP_mult_208_U2177 ( .A1(DP_mult_208_n666), .A2(DP_mult_208_n481), 
        .ZN(DP_mult_208_n315) );
  NAND2_X1 DP_mult_208_U2176 ( .A1(DP_mult_208_n2019), .A2(DP_mult_208_n514), 
        .ZN(DP_mult_208_n318) );
  NAND2_X1 DP_mult_208_U2175 ( .A1(DP_mult_208_n2013), .A2(DP_mult_208_n670), 
        .ZN(DP_mult_208_n319) );
  NAND2_X1 DP_mult_208_U2174 ( .A1(DP_mult_208_n668), .A2(DP_mult_208_n503), 
        .ZN(DP_mult_208_n317) );
  NAND2_X1 DP_mult_208_U2173 ( .A1(DP_mult_208_n671), .A2(DP_mult_208_n532), 
        .ZN(DP_mult_208_n320) );
  XNOR2_X1 DP_mult_208_U2172 ( .A(DP_pipe02[19]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1486) );
  XNOR2_X1 DP_mult_208_U2171 ( .A(DP_pipe02[13]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1492) );
  XNOR2_X1 DP_mult_208_U2170 ( .A(DP_pipe02[21]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1484) );
  XNOR2_X1 DP_mult_208_U2169 ( .A(DP_pipe02[17]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1488) );
  XNOR2_X1 DP_mult_208_U2168 ( .A(DP_pipe02[11]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1494) );
  XNOR2_X1 DP_mult_208_U2167 ( .A(DP_pipe02[15]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1490) );
  XNOR2_X1 DP_mult_208_U2166 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1727) );
  XNOR2_X1 DP_mult_208_U2165 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2241), .ZN(
        DP_mult_208_n1652) );
  XNOR2_X1 DP_mult_208_U2164 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2232), .ZN(
        DP_mult_208_n1702) );
  XNOR2_X1 DP_mult_208_U2163 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1627) );
  XNOR2_X1 DP_mult_208_U2162 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2250), .ZN(
        DP_mult_208_n1602) );
  XNOR2_X1 DP_mult_208_U2161 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2255), .ZN(
        DP_mult_208_n1577) );
  XNOR2_X1 DP_mult_208_U2160 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1502) );
  OAI22_X1 DP_mult_208_U2159 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1678), 
        .B1(DP_mult_208_n1677), .B2(DP_mult_208_n2035), .ZN(DP_mult_208_n1382)
         );
  XNOR2_X1 DP_mult_208_U2158 ( .A(DP_pipe02[9]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1521) );
  XNOR2_X1 DP_mult_208_U2157 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2232), .ZN(
        DP_mult_208_n1704) );
  XNOR2_X1 DP_mult_208_U2156 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1500) );
  XNOR2_X1 DP_mult_208_U2155 ( .A(DP_pipe02[5]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1525) );
  XNOR2_X1 DP_mult_208_U2154 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1729) );
  XNOR2_X1 DP_mult_208_U2153 ( .A(DP_pipe02[1]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1529) );
  XNOR2_X1 DP_mult_208_U2152 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1629) );
  XNOR2_X1 DP_mult_208_U2151 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2233), .ZN(
        DP_mult_208_n1700) );
  XNOR2_X1 DP_mult_208_U2150 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1725) );
  XNOR2_X1 DP_mult_208_U2149 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2261), .ZN(
        DP_mult_208_n1550) );
  XNOR2_X1 DP_mult_208_U2148 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2241), .ZN(
        DP_mult_208_n1654) );
  XNOR2_X1 DP_mult_208_U2147 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2241), .ZN(
        DP_mult_208_n1650) );
  XNOR2_X1 DP_mult_208_U2146 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2250), .ZN(
        DP_mult_208_n1604) );
  XNOR2_X1 DP_mult_208_U2145 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2232), .ZN(
        DP_mult_208_n1696) );
  XNOR2_X1 DP_mult_208_U2144 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1721) );
  XNOR2_X1 DP_mult_208_U2143 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1625) );
  XNOR2_X1 DP_mult_208_U2142 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2255), .ZN(
        DP_mult_208_n1579) );
  XNOR2_X1 DP_mult_208_U2141 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2241), .ZN(
        DP_mult_208_n1646) );
  XNOR2_X1 DP_mult_208_U2140 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2261), .ZN(
        DP_mult_208_n1554) );
  XNOR2_X1 DP_mult_208_U2139 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2250), .ZN(
        DP_mult_208_n1600) );
  XNOR2_X1 DP_mult_208_U2138 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2250), .ZN(
        DP_mult_208_n1596) );
  XNOR2_X1 DP_mult_208_U2137 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1621) );
  XNOR2_X1 DP_mult_208_U2136 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2255), .ZN(
        DP_mult_208_n1575) );
  XNOR2_X1 DP_mult_208_U2135 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2255), .ZN(
        DP_mult_208_n1571) );
  XNOR2_X1 DP_mult_208_U2134 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2262), .ZN(
        DP_mult_208_n1546) );
  XNOR2_X1 DP_mult_208_U2133 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1496) );
  XNOR2_X1 DP_mult_208_U2132 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2261), .ZN(
        DP_mult_208_n1548) );
  XNOR2_X1 DP_mult_208_U2131 ( .A(DP_pipe02[7]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1523) );
  XNOR2_X1 DP_mult_208_U2130 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2232), .ZN(
        DP_mult_208_n1698) );
  XNOR2_X1 DP_mult_208_U2129 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1723) );
  XNOR2_X1 DP_mult_208_U2128 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2241), .ZN(
        DP_mult_208_n1648) );
  XNOR2_X1 DP_mult_208_U2127 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1623) );
  XNOR2_X1 DP_mult_208_U2126 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2250), .ZN(
        DP_mult_208_n1598) );
  XNOR2_X1 DP_mult_208_U2125 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2255), .ZN(
        DP_mult_208_n1573) );
  XNOR2_X1 DP_mult_208_U2124 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2020), .ZN(
        DP_mult_208_n1498) );
  XNOR2_X1 DP_mult_208_U2123 ( .A(DP_pipe02[3]), .B(DP_mult_208_n2065), .ZN(
        DP_mult_208_n1752) );
  XNOR2_X1 DP_mult_208_U2122 ( .A(DP_pipe02[23]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1507) );
  XNOR2_X1 DP_mult_208_U2121 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2262), .ZN(
        DP_mult_208_n1532) );
  XNOR2_X1 DP_mult_208_U2120 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2065), .ZN(
        DP_mult_208_n1732) );
  XNOR2_X1 DP_mult_208_U2119 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2226), .ZN(
        DP_mult_208_n1707) );
  XNOR2_X1 DP_mult_208_U2118 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2250), .ZN(
        DP_mult_208_n1582) );
  XNOR2_X1 DP_mult_208_U2117 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2008), .ZN(
        DP_mult_208_n1607) );
  XNOR2_X1 DP_mult_208_U2116 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2255), .ZN(
        DP_mult_208_n1557) );
  XNOR2_X1 DP_mult_208_U2115 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2231), .ZN(
        DP_mult_208_n1682) );
  XNOR2_X1 DP_mult_208_U2114 ( .A(DP_pipe02[23]), .B(DP_mult_208_n2241), .ZN(
        DP_mult_208_n1632) );
  XNOR2_X1 DP_mult_208_U2113 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2064), .ZN(
        DP_mult_208_n1754) );
  XNOR2_X1 DP_mult_208_U2112 ( .A(DP_pipe02[5]), .B(DP_mult_208_n2065), .ZN(
        DP_mult_208_n1750) );
  XNOR2_X1 DP_mult_208_U2111 ( .A(DP_pipe02[9]), .B(DP_mult_208_n2064), .ZN(
        DP_mult_208_n1746) );
  XNOR2_X1 DP_mult_208_U2110 ( .A(DP_mult_208_n2227), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1728) );
  XNOR2_X1 DP_mult_208_U2109 ( .A(DP_mult_208_n2242), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1653) );
  XNOR2_X1 DP_mult_208_U2108 ( .A(DP_mult_208_n2232), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1703) );
  XNOR2_X1 DP_mult_208_U2107 ( .A(DP_mult_208_n2246), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1628) );
  XNOR2_X1 DP_mult_208_U2106 ( .A(DP_mult_208_n2251), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1603) );
  XNOR2_X1 DP_mult_208_U2105 ( .A(DP_mult_208_n2256), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1578) );
  XNOR2_X1 DP_mult_208_U2104 ( .A(DP_mult_208_n2020), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1503) );
  XNOR2_X1 DP_mult_208_U2103 ( .A(DP_pipe02[7]), .B(DP_mult_208_n2064), .ZN(
        DP_mult_208_n1748) );
  XNOR2_X1 DP_mult_208_U2102 ( .A(DP_mult_208_n2020), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1483) );
  XNOR2_X1 DP_mult_208_U2101 ( .A(DP_mult_208_n2266), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1522) );
  XNOR2_X1 DP_mult_208_U2100 ( .A(DP_mult_208_n2243), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1639) );
  XNOR2_X1 DP_mult_208_U2099 ( .A(DP_mult_208_n2242), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1637) );
  XNOR2_X1 DP_mult_208_U2098 ( .A(DP_mult_208_n2020), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1501) );
  XNOR2_X1 DP_mult_208_U2097 ( .A(DP_mult_208_n2260), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1547) );
  XNOR2_X1 DP_mult_208_U2096 ( .A(DP_mult_208_n2020), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1493) );
  XNOR2_X1 DP_mult_208_U2095 ( .A(DP_mult_208_n2265), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1524) );
  XNOR2_X1 DP_mult_208_U2094 ( .A(DP_mult_208_n2261), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1549) );
  XNOR2_X1 DP_mult_208_U2093 ( .A(DP_mult_208_n2227), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1722) );
  XNOR2_X1 DP_mult_208_U2092 ( .A(DP_mult_208_n2227), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1726) );
  XNOR2_X1 DP_mult_208_U2091 ( .A(DP_mult_208_n2233), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1701) );
  XNOR2_X1 DP_mult_208_U2090 ( .A(DP_mult_208_n2242), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1651) );
  XNOR2_X1 DP_mult_208_U2089 ( .A(DP_mult_208_n2233), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1697) );
  XNOR2_X1 DP_mult_208_U2088 ( .A(DP_mult_208_n2233), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1699) );
  XNOR2_X1 DP_mult_208_U2087 ( .A(DP_mult_208_n2262), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1551) );
  XNOR2_X1 DP_mult_208_U2086 ( .A(DP_mult_208_n2242), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1643) );
  XNOR2_X1 DP_mult_208_U2085 ( .A(DP_mult_208_n2227), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1724) );
  XNOR2_X1 DP_mult_208_U2084 ( .A(DP_mult_208_n2266), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1520) );
  XNOR2_X1 DP_mult_208_U2083 ( .A(DP_mult_208_n2246), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1612) );
  XNOR2_X1 DP_mult_208_U2082 ( .A(DP_mult_208_n2243), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1635) );
  XNOR2_X1 DP_mult_208_U2081 ( .A(DP_mult_208_n2262), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1543) );
  XNOR2_X1 DP_mult_208_U2080 ( .A(DP_mult_208_n2246), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1626) );
  XNOR2_X1 DP_mult_208_U2079 ( .A(DP_mult_208_n2242), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1649) );
  XNOR2_X1 DP_mult_208_U2078 ( .A(DP_mult_208_n2266), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1518) );
  XNOR2_X1 DP_mult_208_U2077 ( .A(DP_mult_208_n2232), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1695) );
  XNOR2_X1 DP_mult_208_U2076 ( .A(DP_mult_208_n2227), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1718) );
  XNOR2_X1 DP_mult_208_U2075 ( .A(DP_mult_208_n2227), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1720) );
  XNOR2_X1 DP_mult_208_U2074 ( .A(DP_mult_208_n2242), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1645) );
  XNOR2_X1 DP_mult_208_U2073 ( .A(DP_mult_208_n2246), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1624) );
  XNOR2_X1 DP_mult_208_U2072 ( .A(DP_mult_208_n2233), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1693) );
  XNOR2_X1 DP_mult_208_U2071 ( .A(DP_mult_208_n2242), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1647) );
  XNOR2_X1 DP_mult_208_U2070 ( .A(DP_mult_208_n2223), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1739) );
  XNOR2_X1 DP_mult_208_U2069 ( .A(DP_mult_208_n2251), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1601) );
  XNOR2_X1 DP_mult_208_U2068 ( .A(DP_mult_208_n2265), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1508) );
  XNOR2_X1 DP_mult_208_U2067 ( .A(DP_mult_208_n2256), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1576) );
  XNOR2_X1 DP_mult_208_U2066 ( .A(DP_mult_208_n2246), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1622) );
  XNOR2_X1 DP_mult_208_U2065 ( .A(DP_mult_208_n2251), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1599) );
  XNOR2_X1 DP_mult_208_U2064 ( .A(DP_mult_208_n2228), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1714) );
  XNOR2_X1 DP_mult_208_U2063 ( .A(DP_mult_208_n2231), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1683) );
  XNOR2_X1 DP_mult_208_U2062 ( .A(DP_mult_208_n2228), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1708) );
  XNOR2_X1 DP_mult_208_U2061 ( .A(DP_mult_208_n2228), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1710) );
  XNOR2_X1 DP_mult_208_U2060 ( .A(DP_mult_208_n2246), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1618) );
  XNOR2_X1 DP_mult_208_U2059 ( .A(DP_mult_208_n2222), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1737) );
  XNOR2_X1 DP_mult_208_U2058 ( .A(DP_mult_208_n2233), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1687) );
  XNOR2_X1 DP_mult_208_U2057 ( .A(DP_mult_208_n2237), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1664) );
  XNOR2_X1 DP_mult_208_U2056 ( .A(DP_mult_208_n2256), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1572) );
  XNOR2_X1 DP_mult_208_U2055 ( .A(DP_mult_208_n2223), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1735) );
  XNOR2_X1 DP_mult_208_U2054 ( .A(DP_mult_208_n2251), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1597) );
  XNOR2_X1 DP_mult_208_U2053 ( .A(DP_mult_208_n2256), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1574) );
  XNOR2_X1 DP_mult_208_U2052 ( .A(DP_mult_208_n2266), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1514) );
  XNOR2_X1 DP_mult_208_U2051 ( .A(DP_mult_208_n2020), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1499) );
  XNOR2_X1 DP_mult_208_U2050 ( .A(DP_mult_208_n2020), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1497) );
  XNOR2_X1 DP_mult_208_U2049 ( .A(DP_mult_208_n2256), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1568) );
  XNOR2_X1 DP_mult_208_U2048 ( .A(DP_mult_208_n2251), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1595) );
  XNOR2_X1 DP_mult_208_U2047 ( .A(DP_mult_208_n2223), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1733) );
  XNOR2_X1 DP_mult_208_U2046 ( .A(DP_mult_208_n2236), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1662) );
  XNOR2_X1 DP_mult_208_U2045 ( .A(DP_mult_208_n2227), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1712) );
  XNOR2_X1 DP_mult_208_U2044 ( .A(DP_mult_208_n2247), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1610) );
  XNOR2_X1 DP_mult_208_U2043 ( .A(DP_mult_208_n2237), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1658) );
  XNOR2_X1 DP_mult_208_U2042 ( .A(DP_mult_208_n2252), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1583) );
  XNOR2_X1 DP_mult_208_U2041 ( .A(DP_mult_208_n2020), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1485) );
  XNOR2_X1 DP_mult_208_U2040 ( .A(DP_mult_208_n2246), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1620) );
  XNOR2_X1 DP_mult_208_U2039 ( .A(DP_mult_208_n2261), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1545) );
  XNOR2_X1 DP_mult_208_U2038 ( .A(DP_mult_208_n2247), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1614) );
  XNOR2_X1 DP_mult_208_U2037 ( .A(DP_mult_208_n2020), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1489) );
  XNOR2_X1 DP_mult_208_U2036 ( .A(DP_mult_208_n2257), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1570) );
  XNOR2_X1 DP_mult_208_U2035 ( .A(DP_mult_208_n2237), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1660) );
  XNOR2_X1 DP_mult_208_U2034 ( .A(DP_mult_208_n2247), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1608) );
  XNOR2_X1 DP_mult_208_U2033 ( .A(DP_mult_208_n2232), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1685) );
  XNOR2_X1 DP_mult_208_U2032 ( .A(DP_mult_208_n2251), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1593) );
  XNOR2_X1 DP_mult_208_U2031 ( .A(DP_mult_208_n2232), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1689) );
  XNOR2_X1 DP_mult_208_U2030 ( .A(DP_mult_208_n2020), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1487) );
  XNOR2_X1 DP_mult_208_U2029 ( .A(DP_mult_208_n2266), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1510) );
  XNOR2_X1 DP_mult_208_U2028 ( .A(DP_mult_208_n2265), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1512) );
  XNOR2_X1 DP_mult_208_U2027 ( .A(DP_mult_208_n2252), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1585) );
  XNOR2_X1 DP_mult_208_U2026 ( .A(DP_mult_208_n2262), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1539) );
  XNOR2_X1 DP_mult_208_U2025 ( .A(DP_mult_208_n2262), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1537) );
  XNOR2_X1 DP_mult_208_U2024 ( .A(DP_mult_208_n2252), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1589) );
  XNOR2_X1 DP_mult_208_U2023 ( .A(DP_mult_208_n2260), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1533) );
  XNOR2_X1 DP_mult_208_U2022 ( .A(DP_mult_208_n2251), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1587) );
  XNOR2_X1 DP_mult_208_U2021 ( .A(DP_mult_208_n2020), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1495) );
  XNOR2_X1 DP_mult_208_U2020 ( .A(DP_mult_208_n2260), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1535) );
  XNOR2_X1 DP_mult_208_U2019 ( .A(DP_mult_208_n2265), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1526) );
  XNOR2_X1 DP_mult_208_U2018 ( .A(DP_mult_208_n2243), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1633) );
  XNOR2_X1 DP_mult_208_U2017 ( .A(DP_mult_208_n2219), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1764) );
  XNOR2_X1 DP_mult_208_U2016 ( .A(DP_mult_208_n2218), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1762) );
  XNOR2_X1 DP_mult_208_U2015 ( .A(DP_mult_208_n2219), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1760) );
  XNOR2_X1 DP_mult_208_U2014 ( .A(DP_mult_208_n2219), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1758) );
  XNOR2_X1 DP_mult_208_U2013 ( .A(DP_mult_208_n2265), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1516) );
  XNOR2_X1 DP_mult_208_U2012 ( .A(DP_mult_208_n2242), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1641) );
  XNOR2_X1 DP_mult_208_U2011 ( .A(DP_mult_208_n2222), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1741) );
  XNOR2_X1 DP_mult_208_U2010 ( .A(DP_mult_208_n2227), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1716) );
  XNOR2_X1 DP_mult_208_U2009 ( .A(DP_mult_208_n2251), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1591) );
  XNOR2_X1 DP_mult_208_U2008 ( .A(DP_mult_208_n2232), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1691) );
  XNOR2_X1 DP_mult_208_U2007 ( .A(DP_mult_208_n2237), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1666) );
  XNOR2_X1 DP_mult_208_U2006 ( .A(DP_mult_208_n2246), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1616) );
  XNOR2_X1 DP_mult_208_U2005 ( .A(DP_mult_208_n2262), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1541) );
  XNOR2_X1 DP_mult_208_U2004 ( .A(DP_mult_208_n2020), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1491) );
  XNOR2_X1 DP_mult_208_U2003 ( .A(DP_mult_208_n2218), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1766) );
  XNOR2_X1 DP_mult_208_U2002 ( .A(DP_mult_208_n2218), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1778) );
  XNOR2_X1 DP_mult_208_U2001 ( .A(DP_mult_208_n2222), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1753) );
  XNOR2_X1 DP_mult_208_U2000 ( .A(DP_mult_208_n2218), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1768) );
  XNOR2_X1 DP_mult_208_U1999 ( .A(DP_mult_208_n2236), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1674) );
  XNOR2_X1 DP_mult_208_U1998 ( .A(DP_mult_208_n2257), .B(DP_pipe02[18]), .ZN(
        DP_mult_208_n1562) );
  XNOR2_X1 DP_mult_208_U1997 ( .A(DP_mult_208_n2222), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1743) );
  XNOR2_X1 DP_mult_208_U1996 ( .A(DP_mult_208_n2222), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1751) );
  XNOR2_X1 DP_mult_208_U1995 ( .A(DP_mult_208_n2236), .B(DP_pipe02[12]), .ZN(
        DP_mult_208_n1668) );
  XNOR2_X1 DP_mult_208_U1994 ( .A(DP_mult_208_n2257), .B(DP_pipe02[20]), .ZN(
        DP_mult_208_n1560) );
  XNOR2_X1 DP_mult_208_U1993 ( .A(DP_mult_208_n2257), .B(DP_pipe02[22]), .ZN(
        DP_mult_208_n1558) );
  XNOR2_X1 DP_mult_208_U1992 ( .A(DP_mult_208_n2257), .B(DP_pipe02[16]), .ZN(
        DP_mult_208_n1564) );
  XNOR2_X1 DP_mult_208_U1991 ( .A(DP_mult_208_n2257), .B(DP_pipe02[14]), .ZN(
        DP_mult_208_n1566) );
  XNOR2_X1 DP_mult_208_U1990 ( .A(DP_mult_208_n2237), .B(DP_pipe02[2]), .ZN(
        DP_mult_208_n1678) );
  XNOR2_X1 DP_mult_208_U1989 ( .A(DP_mult_208_n2218), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1776) );
  XNOR2_X1 DP_mult_208_U1988 ( .A(DP_mult_208_n2218), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1772) );
  XNOR2_X1 DP_mult_208_U1987 ( .A(DP_mult_208_n2218), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1774) );
  XNOR2_X1 DP_mult_208_U1986 ( .A(DP_mult_208_n2218), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1770) );
  XNOR2_X1 DP_mult_208_U1985 ( .A(DP_mult_208_n2222), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1747) );
  XNOR2_X1 DP_mult_208_U1984 ( .A(DP_mult_208_n2222), .B(DP_pipe02[6]), .ZN(
        DP_mult_208_n1749) );
  XNOR2_X1 DP_mult_208_U1983 ( .A(DP_mult_208_n2222), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1745) );
  XNOR2_X1 DP_mult_208_U1982 ( .A(DP_mult_208_n2236), .B(DP_pipe02[4]), .ZN(
        DP_mult_208_n1676) );
  XNOR2_X1 DP_mult_208_U1981 ( .A(DP_mult_208_n2236), .B(DP_pipe02[8]), .ZN(
        DP_mult_208_n1672) );
  XNOR2_X1 DP_mult_208_U1980 ( .A(DP_mult_208_n2237), .B(DP_pipe02[10]), .ZN(
        DP_mult_208_n1670) );
  OAI22_X1 DP_mult_208_U1979 ( .A1(DP_mult_208_n1950), .A2(DP_mult_208_n1776), 
        .B1(DP_mult_208_n1775), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1477)
         );
  INV_X1 DP_mult_208_U1978 ( .A(DP_mult_208_n1482), .ZN(DP_mult_208_n2282) );
  OAI21_X1 DP_mult_208_U1977 ( .B1(DP_mult_208_n2145), .B2(DP_mult_208_n2159), 
        .A(DP_mult_208_n2282), .ZN(DP_mult_208_n1194) );
  INV_X1 DP_mult_208_U1976 ( .A(DP_mult_208_n1732), .ZN(DP_mult_208_n2272) );
  INV_X1 DP_mult_208_U1975 ( .A(DP_mult_208_n1582), .ZN(DP_mult_208_n2278) );
  INV_X1 DP_mult_208_U1974 ( .A(DP_mult_208_n1657), .ZN(DP_mult_208_n2275) );
  CLKBUF_X1 DP_mult_208_U1973 ( .A(DP_mult_208_n251), .Z(DP_mult_208_n2215) );
  INV_X1 DP_mult_208_U1972 ( .A(DP_mult_208_n802), .ZN(DP_mult_208_n803) );
  NAND2_X1 DP_mult_208_U1971 ( .A1(DP_mult_208_n2218), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1781) );
  OAI22_X1 DP_mult_208_U1970 ( .A1(DP_mult_208_n1950), .A2(DP_mult_208_n1780), 
        .B1(DP_mult_208_n1779), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1481)
         );
  OAI22_X1 DP_mult_208_U1969 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1750), 
        .B1(DP_mult_208_n2011), .B2(DP_mult_208_n1749), .ZN(DP_mult_208_n1451)
         );
  OAI22_X1 DP_mult_208_U1968 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1773), 
        .B1(DP_mult_208_n1772), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1474)
         );
  OAI22_X1 DP_mult_208_U1967 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1747), 
        .B1(DP_mult_208_n1746), .B2(DP_mult_208_n1937), .ZN(DP_mult_208_n1448)
         );
  OAI22_X1 DP_mult_208_U1966 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1676), 
        .B1(DP_mult_208_n1675), .B2(DP_mult_208_n2035), .ZN(DP_mult_208_n1380)
         );
  OAI22_X1 DP_mult_208_U1965 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1671), 
        .B1(DP_mult_208_n2056), .B2(DP_mult_208_n1670), .ZN(DP_mult_208_n1375)
         );
  INV_X1 DP_mult_208_U1964 ( .A(DP_mult_208_n874), .ZN(DP_mult_208_n875) );
  INV_X1 DP_mult_208_U1963 ( .A(DP_mult_208_n1607), .ZN(DP_mult_208_n2277) );
  OAI21_X1 DP_mult_208_U1962 ( .B1(DP_mult_208_n2143), .B2(DP_mult_208_n2148), 
        .A(DP_mult_208_n2277), .ZN(DP_mult_208_n1314) );
  INV_X1 DP_mult_208_U1961 ( .A(DP_mult_208_n1557), .ZN(DP_mult_208_n2279) );
  NOR2_X1 DP_mult_208_U1960 ( .A1(DP_mult_208_n2003), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1337) );
  NOR2_X1 DP_mult_208_U1959 ( .A1(DP_mult_208_n2012), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1289) );
  INV_X1 DP_mult_208_U1958 ( .A(DP_mult_208_n724), .ZN(DP_mult_208_n725) );
  OAI22_X1 DP_mult_208_U1957 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1749), 
        .B1(DP_mult_208_n1748), .B2(DP_mult_208_n2011), .ZN(DP_mult_208_n1450)
         );
  OAI22_X1 DP_mult_208_U1956 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1670), 
        .B1(DP_mult_208_n1669), .B2(DP_mult_208_n1958), .ZN(DP_mult_208_n1374)
         );
  INV_X1 DP_mult_208_U1955 ( .A(DP_mult_208_n1707), .ZN(DP_mult_208_n2273) );
  NOR2_X1 DP_mult_208_U1954 ( .A1(DP_mult_208_n2202), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1241) );
  OAI22_X1 DP_mult_208_U1953 ( .A1(DP_mult_208_n2184), .A2(DP_mult_208_n1565), 
        .B1(DP_mult_208_n2012), .B2(DP_mult_208_n1564), .ZN(DP_mult_208_n1273)
         );
  NOR2_X1 DP_mult_208_U1952 ( .A1(DP_mult_208_n2211), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1361) );
  NOR2_X1 DP_mult_208_U1951 ( .A1(DP_mult_208_n2203), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1265) );
  OAI22_X1 DP_mult_208_U1950 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1752), 
        .B1(DP_mult_208_n1937), .B2(DP_mult_208_n1751), .ZN(DP_mult_208_n1453)
         );
  OAI22_X1 DP_mult_208_U1949 ( .A1(DP_mult_208_n1950), .A2(DP_mult_208_n1775), 
        .B1(DP_mult_208_n1774), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1476)
         );
  OAI22_X1 DP_mult_208_U1948 ( .A1(DP_mult_208_n1950), .A2(DP_mult_208_n1772), 
        .B1(DP_mult_208_n1771), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1473)
         );
  OAI22_X1 DP_mult_208_U1947 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1669), 
        .B1(DP_mult_208_n2056), .B2(DP_mult_208_n1668), .ZN(DP_mult_208_n1373)
         );
  OAI22_X1 DP_mult_208_U1946 ( .A1(DP_mult_208_n1950), .A2(DP_mult_208_n1774), 
        .B1(DP_mult_208_n1773), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1475)
         );
  OAI22_X1 DP_mult_208_U1945 ( .A1(DP_mult_208_n2120), .A2(DP_mult_208_n1567), 
        .B1(DP_mult_208_n2012), .B2(DP_mult_208_n1566), .ZN(DP_mult_208_n1275)
         );
  OAI22_X1 DP_mult_208_U1944 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1771), 
        .B1(DP_mult_208_n1770), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1472)
         );
  OAI22_X1 DP_mult_208_U1943 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1679), 
        .B1(DP_mult_208_n2035), .B2(DP_mult_208_n1678), .ZN(DP_mult_208_n1383)
         );
  OAI22_X1 DP_mult_208_U1942 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1748), 
        .B1(DP_mult_208_n2011), .B2(DP_mult_208_n1747), .ZN(DP_mult_208_n1449)
         );
  OAI22_X1 DP_mult_208_U1941 ( .A1(DP_mult_208_n2059), .A2(DP_mult_208_n1770), 
        .B1(DP_mult_208_n1769), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1471)
         );
  NOR2_X1 DP_mult_208_U1940 ( .A1(DP_mult_208_n2206), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1313) );
  OAI22_X1 DP_mult_208_U1939 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1673), 
        .B1(DP_mult_208_n1958), .B2(DP_mult_208_n1672), .ZN(DP_mult_208_n1377)
         );
  INV_X1 DP_mult_208_U1938 ( .A(DP_mult_208_n1682), .ZN(DP_mult_208_n2274) );
  OAI21_X1 DP_mult_208_U1937 ( .B1(DP_mult_208_n2146), .B2(DP_mult_208_n2175), 
        .A(DP_mult_208_n2274), .ZN(DP_mult_208_n1386) );
  NOR2_X1 DP_mult_208_U1936 ( .A1(DP_mult_208_n2051), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1217) );
  OAI22_X1 DP_mult_208_U1935 ( .A1(DP_mult_208_n2184), .A2(DP_mult_208_n1561), 
        .B1(DP_mult_208_n2037), .B2(DP_mult_208_n1560), .ZN(DP_mult_208_n1269)
         );
  NAND2_X1 DP_mult_208_U1934 ( .A1(DP_mult_208_n2265), .A2(DP_mult_208_n1965), 
        .ZN(DP_mult_208_n1531) );
  NAND2_X1 DP_mult_208_U1933 ( .A1(DP_mult_208_n2236), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1681) );
  NAND2_X1 DP_mult_208_U1932 ( .A1(DP_mult_208_n2251), .A2(DP_mult_208_n1964), 
        .ZN(DP_mult_208_n1606) );
  NAND2_X1 DP_mult_208_U1931 ( .A1(DP_mult_208_n2233), .A2(DP_mult_208_n1965), 
        .ZN(DP_mult_208_n1706) );
  NAND2_X1 DP_mult_208_U1930 ( .A1(DP_mult_208_n2246), .A2(DP_mult_208_n1965), 
        .ZN(DP_mult_208_n1631) );
  NAND2_X1 DP_mult_208_U1929 ( .A1(DP_mult_208_n2020), .A2(DP_mult_208_n1964), 
        .ZN(DP_mult_208_n1506) );
  NAND2_X1 DP_mult_208_U1928 ( .A1(DP_mult_208_n2242), .A2(DP_mult_208_n1964), 
        .ZN(DP_mult_208_n1656) );
  NAND2_X1 DP_mult_208_U1927 ( .A1(DP_mult_208_n2260), .A2(DP_mult_208_n1965), 
        .ZN(DP_mult_208_n1556) );
  OAI22_X1 DP_mult_208_U1926 ( .A1(DP_mult_208_n2184), .A2(DP_mult_208_n1559), 
        .B1(DP_mult_208_n2037), .B2(DP_mult_208_n1558), .ZN(DP_mult_208_n1267)
         );
  OAI22_X1 DP_mult_208_U1925 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1672), 
        .B1(DP_mult_208_n1671), .B2(DP_mult_208_n2035), .ZN(DP_mult_208_n1376)
         );
  INV_X1 DP_mult_208_U1924 ( .A(DP_mult_208_n1632), .ZN(DP_mult_208_n2276) );
  OAI22_X1 DP_mult_208_U1923 ( .A1(DP_mult_208_n2120), .A2(DP_mult_208_n1563), 
        .B1(DP_mult_208_n2037), .B2(DP_mult_208_n1562), .ZN(DP_mult_208_n1271)
         );
  NOR2_X1 DP_mult_208_U1922 ( .A1(DP_mult_208_n1181), .A2(DP_mult_208_n1192), 
        .ZN(DP_mult_208_n644) );
  NAND2_X1 DP_mult_208_U1921 ( .A1(DP_mult_208_n1181), .A2(DP_mult_208_n1192), 
        .ZN(DP_mult_208_n645) );
  NAND2_X1 DP_mult_208_U1920 ( .A1(DP_mult_208_n2257), .A2(DP_mult_208_n1965), 
        .ZN(DP_mult_208_n1581) );
  OAI22_X1 DP_mult_208_U1919 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1754), 
        .B1(DP_mult_208_n2011), .B2(DP_mult_208_n1753), .ZN(DP_mult_208_n1455)
         );
  OAI22_X1 DP_mult_208_U1918 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1777), 
        .B1(DP_mult_208_n1776), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1478)
         );
  OAI22_X1 DP_mult_208_U1917 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1745), 
        .B1(DP_mult_208_n1744), .B2(DP_mult_208_n2011), .ZN(DP_mult_208_n1446)
         );
  INV_X1 DP_mult_208_U1916 ( .A(DP_mult_208_n2054), .ZN(DP_mult_208_n2203) );
  NOR2_X1 DP_mult_208_U1915 ( .A1(DP_mult_208_n2213), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1433) );
  OAI22_X1 DP_mult_208_U1914 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1744), 
        .B1(DP_mult_208_n2011), .B2(DP_mult_208_n1743), .ZN(DP_mult_208_n1445)
         );
  OAI22_X1 DP_mult_208_U1913 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1675), 
        .B1(DP_mult_208_n2035), .B2(DP_mult_208_n1674), .ZN(DP_mult_208_n1379)
         );
  OAI22_X1 DP_mult_208_U1912 ( .A1(DP_mult_208_n2100), .A2(DP_mult_208_n1746), 
        .B1(DP_mult_208_n1937), .B2(DP_mult_208_n1745), .ZN(DP_mult_208_n1447)
         );
  OAI22_X1 DP_mult_208_U1911 ( .A1(DP_mult_208_n2059), .A2(DP_mult_208_n1769), 
        .B1(DP_mult_208_n1768), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1470)
         );
  OAI22_X1 DP_mult_208_U1910 ( .A1(DP_mult_208_n2190), .A2(DP_mult_208_n1677), 
        .B1(DP_mult_208_n2056), .B2(DP_mult_208_n1676), .ZN(DP_mult_208_n1381)
         );
  NOR2_X1 DP_mult_208_U1909 ( .A1(DP_mult_208_n2048), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1409) );
  INV_X1 DP_mult_208_U1908 ( .A(DP_mult_208_n1532), .ZN(DP_mult_208_n2280) );
  OAI21_X1 DP_mult_208_U1907 ( .B1(DP_mult_208_n2066), .B2(DP_mult_208_n2054), 
        .A(DP_mult_208_n2280), .ZN(DP_mult_208_n1242) );
  NOR2_X1 DP_mult_208_U1906 ( .A1(DP_mult_208_n2035), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1385) );
  NAND2_X1 DP_mult_208_U1905 ( .A1(DP_mult_208_n2227), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1731) );
  INV_X1 DP_mult_208_U1904 ( .A(DP_mult_208_n682), .ZN(DP_mult_208_n683) );
  INV_X1 DP_mult_208_U1903 ( .A(DP_mult_208_n1507), .ZN(DP_mult_208_n2281) );
  OAI21_X1 DP_mult_208_U1902 ( .B1(DP_mult_208_n2144), .B2(DP_mult_208_n2045), 
        .A(DP_mult_208_n2281), .ZN(DP_mult_208_n1218) );
  NOR2_X1 DP_mult_208_U1901 ( .A1(DP_mult_208_n2011), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1457) );
  INV_X1 DP_mult_208_U1900 ( .A(DP_mult_208_n2244), .ZN(DP_mult_208_n2242) );
  OAI22_X1 DP_mult_208_U1899 ( .A1(DP_mult_208_n2198), .A2(DP_mult_208_n1779), 
        .B1(DP_mult_208_n1778), .B2(DP_mult_208_n1960), .ZN(DP_mult_208_n1480)
         );
  NAND2_X1 DP_mult_208_U1898 ( .A1(DP_mult_208_n2222), .A2(DP_mult_208_n1955), 
        .ZN(DP_mult_208_n1756) );
  OR2_X1 DP_mult_208_U1897 ( .A1(DP_mult_208_n1194), .A2(DP_mult_208_n676), 
        .ZN(DP_mult_208_n2137) );
  NAND2_X1 DP_mult_208_U1896 ( .A1(DP_mult_208_n678), .A2(DP_mult_208_n677), 
        .ZN(DP_mult_208_n335) );
  NAND2_X1 DP_mult_208_U1895 ( .A1(DP_mult_208_n1159), .A2(DP_mult_208_n1161), 
        .ZN(DP_mult_208_n627) );
  NAND2_X1 DP_mult_208_U1894 ( .A1(DP_mult_208_n1175), .A2(DP_mult_208_n1178), 
        .ZN(DP_mult_208_n637) );
  NAND2_X1 DP_mult_208_U1893 ( .A1(DP_mult_208_n1165), .A2(DP_mult_208_n1170), 
        .ZN(DP_mult_208_n632) );
  NOR2_X1 DP_mult_208_U1892 ( .A1(DP_mult_208_n1159), .A2(DP_mult_208_n1161), 
        .ZN(DP_mult_208_n626) );
  OR2_X1 DP_mult_208_U1891 ( .A1(DP_mult_208_n685), .A2(DP_mult_208_n688), 
        .ZN(DP_mult_208_n2136) );
  NAND2_X1 DP_mult_208_U1890 ( .A1(DP_mult_208_n679), .A2(DP_mult_208_n680), 
        .ZN(DP_mult_208_n341) );
  NAND2_X1 DP_mult_208_U1889 ( .A1(DP_mult_208_n685), .A2(DP_mult_208_n688), 
        .ZN(DP_mult_208_n369) );
  NAND2_X1 DP_mult_208_U1888 ( .A1(DP_mult_208_n681), .A2(DP_mult_208_n684), 
        .ZN(DP_mult_208_n352) );
  NOR2_X1 DP_mult_208_U1887 ( .A1(DP_mult_208_n678), .A2(DP_mult_208_n677), 
        .ZN(DP_mult_208_n334) );
  OR2_X1 DP_mult_208_U1886 ( .A1(DP_mult_208_n679), .A2(DP_mult_208_n680), 
        .ZN(DP_mult_208_n2134) );
  NOR2_X1 DP_mult_208_U1885 ( .A1(DP_mult_208_n1175), .A2(DP_mult_208_n1178), 
        .ZN(DP_mult_208_n636) );
  AOI21_X1 DP_mult_208_U1884 ( .B1(DP_mult_208_n1972), .B2(DP_mult_208_n1970), 
        .A(DP_mult_208_n1981), .ZN(DP_mult_208_n646) );
  OAI21_X1 DP_mult_208_U1883 ( .B1(DP_mult_208_n646), .B2(DP_mult_208_n644), 
        .A(DP_mult_208_n645), .ZN(DP_mult_208_n643) );
  AOI21_X1 DP_mult_208_U1882 ( .B1(DP_mult_208_n643), .B2(DP_mult_208_n1973), 
        .A(DP_mult_208_n1983), .ZN(DP_mult_208_n638) );
  AND2_X1 DP_mult_208_U1881 ( .A1(DP_mult_208_n1194), .A2(DP_mult_208_n676), 
        .ZN(DP_mult_208_n2133) );
  NOR2_X1 DP_mult_208_U1880 ( .A1(DP_mult_208_n1165), .A2(DP_mult_208_n1170), 
        .ZN(DP_mult_208_n631) );
  INV_X1 DP_mult_208_U1879 ( .A(DP_mult_208_n676), .ZN(DP_mult_208_n677) );
  NAND2_X1 DP_mult_208_U1878 ( .A1(DP_mult_208_n2135), .A2(DP_mult_208_n352), 
        .ZN(DP_mult_208_n303) );
  NAND2_X1 DP_mult_208_U1877 ( .A1(DP_mult_208_n2134), .A2(DP_mult_208_n341), 
        .ZN(DP_mult_208_n302) );
  NAND2_X1 DP_mult_208_U1876 ( .A1(DP_mult_208_n2130), .A2(DP_mult_208_n1989), 
        .ZN(DP_mult_208_n599) );
  NAND2_X1 DP_mult_208_U1875 ( .A1(DP_mult_208_n2121), .A2(DP_mult_208_n2132), 
        .ZN(DP_mult_208_n610) );
  NAND2_X1 DP_mult_208_U1874 ( .A1(DP_mult_208_n1085), .A2(DP_mult_208_n1098), 
        .ZN(DP_mult_208_n593) );
  NAND2_X1 DP_mult_208_U1873 ( .A1(DP_mult_208_n2136), .A2(DP_mult_208_n369), 
        .ZN(DP_mult_208_n304) );
  INV_X1 DP_mult_208_U1872 ( .A(DP_mult_208_n369), .ZN(DP_mult_208_n367) );
  NAND2_X1 DP_mult_208_U1871 ( .A1(DP_mult_208_n694), .A2(DP_mult_208_n689), 
        .ZN(DP_mult_208_n378) );
  NAND2_X1 DP_mult_208_U1870 ( .A1(DP_mult_208_n1099), .A2(DP_mult_208_n1110), 
        .ZN(DP_mult_208_n598) );
  NOR2_X1 DP_mult_208_U1869 ( .A1(DP_mult_208_n336), .A2(DP_mult_208_n334), 
        .ZN(DP_mult_208_n332) );
  NAND2_X1 DP_mult_208_U1868 ( .A1(DP_mult_208_n701), .A2(DP_mult_208_n708), 
        .ZN(DP_mult_208_n396) );
  NOR2_X1 DP_mult_208_U1867 ( .A1(DP_mult_208_n1085), .A2(DP_mult_208_n1098), 
        .ZN(DP_mult_208_n592) );
  NOR2_X1 DP_mult_208_U1866 ( .A1(DP_mult_208_n590), .A2(DP_mult_208_n592), 
        .ZN(DP_mult_208_n588) );
  NAND2_X1 DP_mult_208_U1865 ( .A1(DP_mult_208_n588), .A2(DP_mult_208_n2124), 
        .ZN(DP_mult_208_n582) );
  NAND2_X1 DP_mult_208_U1864 ( .A1(DP_mult_208_n695), .A2(DP_mult_208_n700), 
        .ZN(DP_mult_208_n387) );
  OR2_X1 DP_mult_208_U1863 ( .A1(DP_mult_208_n1133), .A2(DP_mult_208_n1142), 
        .ZN(DP_mult_208_n2132) );
  INV_X1 DP_mult_208_U1862 ( .A(DP_mult_208_n341), .ZN(DP_mult_208_n339) );
  AOI21_X1 DP_mult_208_U1861 ( .B1(DP_mult_208_n346), .B2(DP_mult_208_n2134), 
        .A(DP_mult_208_n339), .ZN(DP_mult_208_n337) );
  OR2_X2 DP_mult_208_U1860 ( .A1(DP_mult_208_n694), .A2(DP_mult_208_n689), 
        .ZN(DP_mult_208_n2131) );
  AOI21_X1 DP_mult_208_U1859 ( .B1(DP_mult_208_n2132), .B2(DP_mult_208_n1974), 
        .A(DP_mult_208_n1984), .ZN(DP_mult_208_n611) );
  AOI21_X1 DP_mult_208_U1858 ( .B1(DP_mult_208_n376), .B2(DP_mult_208_n2136), 
        .A(DP_mult_208_n367), .ZN(DP_mult_208_n365) );
  OAI21_X1 DP_mult_208_U1857 ( .B1(DP_mult_208_n364), .B2(DP_mult_208_n387), 
        .A(DP_mult_208_n365), .ZN(DP_mult_208_n363) );
  NAND2_X1 DP_mult_208_U1856 ( .A1(DP_mult_208_n821), .A2(DP_mult_208_n838), 
        .ZN(DP_mult_208_n503) );
  OR2_X1 DP_mult_208_U1855 ( .A1(DP_mult_208_n1111), .A2(DP_mult_208_n1122), 
        .ZN(DP_mult_208_n2130) );
  NOR2_X1 DP_mult_208_U1854 ( .A1(DP_mult_208_n1099), .A2(DP_mult_208_n1110), 
        .ZN(DP_mult_208_n597) );
  OR2_X2 DP_mult_208_U1853 ( .A1(DP_mult_208_n709), .A2(DP_mult_208_n716), 
        .ZN(DP_mult_208_n2129) );
  OR2_X2 DP_mult_208_U1852 ( .A1(DP_mult_208_n701), .A2(DP_mult_208_n708), 
        .ZN(DP_mult_208_n2128) );
  OAI21_X1 DP_mult_208_U1851 ( .B1(DP_mult_208_n638), .B2(DP_mult_208_n636), 
        .A(DP_mult_208_n637), .ZN(DP_mult_208_n635) );
  OAI21_X1 DP_mult_208_U1850 ( .B1(DP_mult_208_n631), .B2(DP_mult_208_n634), 
        .A(DP_mult_208_n632), .ZN(DP_mult_208_n630) );
  NOR2_X1 DP_mult_208_U1849 ( .A1(DP_mult_208_n633), .A2(DP_mult_208_n631), 
        .ZN(DP_mult_208_n629) );
  INV_X1 DP_mult_208_U1848 ( .A(DP_mult_208_n352), .ZN(DP_mult_208_n350) );
  OAI21_X1 DP_mult_208_U1847 ( .B1(DP_mult_208_n421), .B2(DP_mult_208_n347), 
        .A(DP_mult_208_n348), .ZN(DP_mult_208_n346) );
  OR2_X2 DP_mult_208_U1846 ( .A1(DP_mult_208_n717), .A2(DP_mult_208_n726), 
        .ZN(DP_mult_208_n2127) );
  AOI21_X1 DP_mult_208_U1845 ( .B1(DP_mult_208_n625), .B2(DP_mult_208_n1988), 
        .A(DP_mult_208_n1976), .ZN(DP_mult_208_n620) );
  NOR2_X1 DP_mult_208_U1844 ( .A1(DP_mult_208_n695), .A2(DP_mult_208_n700), 
        .ZN(DP_mult_208_n384) );
  XOR2_X1 DP_mult_208_U1843 ( .A(DP_mult_208_n827), .B(DP_mult_208_n844), .Z(
        DP_mult_208_n2167) );
  XNOR2_X1 DP_mult_208_U1842 ( .A(DP_mult_208_n840), .B(DP_mult_208_n825), 
        .ZN(DP_mult_208_n2126) );
  XNOR2_X1 DP_mult_208_U1841 ( .A(DP_mult_208_n2126), .B(DP_mult_208_n823), 
        .ZN(DP_mult_208_n821) );
  NAND2_X1 DP_mult_208_U1840 ( .A1(DP_mult_208_n2125), .A2(DP_mult_208_n1982), 
        .ZN(DP_mult_208_n571) );
  NAND2_X1 DP_mult_208_U1839 ( .A1(DP_mult_208_n2128), .A2(DP_mult_208_n396), 
        .ZN(DP_mult_208_n307) );
  INV_X1 DP_mult_208_U1838 ( .A(DP_mult_208_n384), .ZN(DP_mult_208_n657) );
  NAND2_X1 DP_mult_208_U1837 ( .A1(DP_mult_208_n657), .A2(DP_mult_208_n387), 
        .ZN(DP_mult_208_n306) );
  INV_X1 DP_mult_208_U1836 ( .A(DP_mult_208_n396), .ZN(DP_mult_208_n394) );
  NAND2_X1 DP_mult_208_U1835 ( .A1(DP_mult_208_n2129), .A2(DP_mult_208_n409), 
        .ZN(DP_mult_208_n308) );
  INV_X1 DP_mult_208_U1834 ( .A(DP_mult_208_n428), .ZN(DP_mult_208_n661) );
  NAND2_X1 DP_mult_208_U1833 ( .A1(DP_mult_208_n661), .A2(DP_mult_208_n429), 
        .ZN(DP_mult_208_n310) );
  NAND2_X1 DP_mult_208_U1832 ( .A1(DP_mult_208_n1003), .A2(DP_mult_208_n1020), 
        .ZN(DP_mult_208_n570) );
  NAND2_X1 DP_mult_208_U1831 ( .A1(DP_mult_208_n400), .A2(DP_mult_208_n2128), 
        .ZN(DP_mult_208_n389) );
  OR2_X1 DP_mult_208_U1830 ( .A1(DP_mult_208_n1021), .A2(DP_mult_208_n1038), 
        .ZN(DP_mult_208_n2125) );
  NOR2_X1 DP_mult_208_U1829 ( .A1(DP_mult_208_n389), .A2(DP_mult_208_n384), 
        .ZN(DP_mult_208_n382) );
  OR2_X1 DP_mult_208_U1828 ( .A1(DP_mult_208_n1055), .A2(DP_mult_208_n1070), 
        .ZN(DP_mult_208_n2124) );
  INV_X1 DP_mult_208_U1827 ( .A(DP_mult_208_n378), .ZN(DP_mult_208_n376) );
  NAND2_X1 DP_mult_208_U1826 ( .A1(DP_mult_208_n983), .A2(DP_mult_208_n1002), 
        .ZN(DP_mult_208_n564) );
  INV_X1 DP_mult_208_U1825 ( .A(DP_mult_208_n418), .ZN(DP_mult_208_n416) );
  OR2_X1 DP_mult_208_U1824 ( .A1(DP_mult_208_n761), .A2(DP_mult_208_n774), 
        .ZN(DP_mult_208_n2123) );
  OAI21_X1 DP_mult_208_U1823 ( .B1(DP_mult_208_n620), .B2(DP_mult_208_n610), 
        .A(DP_mult_208_n611), .ZN(DP_mult_208_n609) );
  NOR2_X1 DP_mult_208_U1822 ( .A1(DP_mult_208_n597), .A2(DP_mult_208_n599), 
        .ZN(DP_mult_208_n595) );
  OAI21_X1 DP_mult_208_U1821 ( .B1(DP_mult_208_n600), .B2(DP_mult_208_n597), 
        .A(DP_mult_208_n598), .ZN(DP_mult_208_n596) );
  AOI21_X1 DP_mult_208_U1820 ( .B1(DP_mult_208_n595), .B2(DP_mult_208_n609), 
        .A(DP_mult_208_n596), .ZN(DP_mult_208_n594) );
  NAND2_X1 DP_mult_208_U1819 ( .A1(DP_mult_208_n919), .A2(DP_mult_208_n940), 
        .ZN(DP_mult_208_n543) );
  NOR2_X1 DP_mult_208_U1818 ( .A1(DP_mult_208_n384), .A2(DP_mult_208_n364), 
        .ZN(DP_mult_208_n362) );
  NAND2_X1 DP_mult_208_U1817 ( .A1(DP_mult_208_n963), .A2(DP_mult_208_n982), 
        .ZN(DP_mult_208_n559) );
  NOR2_X1 DP_mult_208_U1816 ( .A1(DP_mult_208_n983), .A2(DP_mult_208_n1002), 
        .ZN(DP_mult_208_n563) );
  NAND2_X1 DP_mult_208_U1815 ( .A1(DP_mult_208_n877), .A2(DP_mult_208_n896), 
        .ZN(DP_mult_208_n532) );
  INV_X1 DP_mult_208_U1814 ( .A(DP_mult_208_n502), .ZN(DP_mult_208_n668) );
  NAND2_X1 DP_mult_208_U1813 ( .A1(DP_mult_208_n857), .A2(DP_mult_208_n876), 
        .ZN(DP_mult_208_n521) );
  NAND2_X1 DP_mult_208_U1812 ( .A1(DP_mult_208_n749), .A2(DP_mult_208_n760), 
        .ZN(DP_mult_208_n439) );
  NAND2_X1 DP_mult_208_U1811 ( .A1(DP_mult_208_n737), .A2(DP_mult_208_n748), 
        .ZN(DP_mult_208_n436) );
  NOR2_X1 DP_mult_208_U1810 ( .A1(DP_mult_208_n737), .A2(DP_mult_208_n748), 
        .ZN(DP_mult_208_n435) );
  NAND2_X1 DP_mult_208_U1809 ( .A1(DP_mult_208_n789), .A2(DP_mult_208_n804), 
        .ZN(DP_mult_208_n481) );
  INV_X1 DP_mult_208_U1808 ( .A(DP_mult_208_n503), .ZN(DP_mult_208_n501) );
  INV_X1 DP_mult_208_U1807 ( .A(DP_mult_208_n409), .ZN(DP_mult_208_n407) );
  AOI21_X1 DP_mult_208_U1806 ( .B1(DP_mult_208_n2129), .B2(DP_mult_208_n416), 
        .A(DP_mult_208_n407), .ZN(DP_mult_208_n405) );
  AOI21_X1 DP_mult_208_U1805 ( .B1(DP_mult_208_n526), .B2(DP_mult_208_n511), 
        .A(DP_mult_208_n2110), .ZN(DP_mult_208_n506) );
  NAND2_X1 DP_mult_208_U1804 ( .A1(DP_mult_208_n507), .A2(DP_mult_208_n668), 
        .ZN(DP_mult_208_n498) );
  INV_X1 DP_mult_208_U1803 ( .A(DP_mult_208_n461), .ZN(DP_mult_208_n459) );
  INV_X1 DP_mult_208_U1802 ( .A(DP_mult_208_n553), .ZN(DP_mult_208_n555) );
  NAND2_X1 DP_mult_208_U1801 ( .A1(DP_mult_208_n663), .A2(DP_mult_208_n439), 
        .ZN(DP_mult_208_n312) );
  INV_X1 DP_mult_208_U1800 ( .A(DP_mult_208_n564), .ZN(DP_mult_208_n562) );
  INV_X1 DP_mult_208_U1799 ( .A(DP_mult_208_n563), .ZN(DP_mult_208_n561) );
  NAND2_X1 DP_mult_208_U1798 ( .A1(DP_mult_208_n662), .A2(DP_mult_208_n436), 
        .ZN(DP_mult_208_n311) );
  INV_X1 DP_mult_208_U1797 ( .A(DP_mult_208_n421), .ZN(DP_mult_208_n423) );
  NAND2_X1 DP_mult_208_U1796 ( .A1(DP_mult_208_n666), .A2(DP_mult_208_n2122), 
        .ZN(DP_mult_208_n467) );
  NAND2_X1 DP_mult_208_U1795 ( .A1(DP_mult_208_n426), .A2(DP_mult_208_n663), 
        .ZN(DP_mult_208_n420) );
  INV_X1 DP_mult_208_U1794 ( .A(DP_mult_208_n439), .ZN(DP_mult_208_n445) );
  NOR2_X1 DP_mult_208_U1793 ( .A1(DP_mult_208_n402), .A2(DP_mult_208_n360), 
        .ZN(DP_mult_208_n356) );
  OAI21_X1 DP_mult_208_U1792 ( .B1(DP_mult_208_n421), .B2(DP_mult_208_n402), 
        .A(DP_mult_208_n405), .ZN(DP_mult_208_n401) );
  NOR2_X1 DP_mult_208_U1791 ( .A1(DP_mult_208_n420), .A2(DP_mult_208_n402), 
        .ZN(DP_mult_208_n400) );
  INV_X1 DP_mult_208_U1790 ( .A(DP_mult_208_n521), .ZN(DP_mult_208_n519) );
  INV_X1 DP_mult_208_U1789 ( .A(DP_mult_208_n481), .ZN(DP_mult_208_n483) );
  OAI21_X1 DP_mult_208_U1788 ( .B1(DP_mult_208_n492), .B2(DP_mult_208_n467), 
        .A(DP_mult_208_n468), .ZN(DP_mult_208_n466) );
  INV_X1 DP_mult_208_U1787 ( .A(DP_mult_208_n436), .ZN(DP_mult_208_n434) );
  AOI21_X1 DP_mult_208_U1786 ( .B1(DP_mult_208_n662), .B2(DP_mult_208_n445), 
        .A(DP_mult_208_n434), .ZN(DP_mult_208_n432) );
  NAND2_X1 DP_mult_208_U1785 ( .A1(DP_mult_208_n663), .A2(DP_mult_208_n662), 
        .ZN(DP_mult_208_n431) );
  INV_X1 DP_mult_208_U1784 ( .A(DP_mult_208_n438), .ZN(DP_mult_208_n663) );
  OAI21_X1 DP_mult_208_U1783 ( .B1(DP_mult_208_n1954), .B2(DP_mult_208_n564), 
        .A(DP_mult_208_n559), .ZN(DP_mult_208_n553) );
  INV_X1 DP_mult_208_U1782 ( .A(DP_mult_208_n552), .ZN(DP_mult_208_n554) );
  INV_X1 DP_mult_208_U1781 ( .A(DP_mult_208_n420), .ZN(DP_mult_208_n422) );
  NOR2_X1 DP_mult_208_U1780 ( .A1(DP_mult_208_n491), .A2(DP_mult_208_n467), 
        .ZN(DP_mult_208_n465) );
  AOI21_X1 DP_mult_208_U1779 ( .B1(DP_mult_208_n565), .B2(DP_mult_208_n552), 
        .A(DP_mult_208_n2009), .ZN(DP_mult_208_n551) );
  INV_X1 DP_mult_208_U1778 ( .A(DP_mult_208_n505), .ZN(DP_mult_208_n507) );
  INV_X1 DP_mult_208_U1777 ( .A(DP_mult_208_n401), .ZN(DP_mult_208_n399) );
  INV_X1 DP_mult_208_U1776 ( .A(DP_mult_208_n400), .ZN(DP_mult_208_n398) );
  NAND2_X1 DP_mult_208_U1775 ( .A1(DP_mult_208_n465), .A2(DP_mult_208_n507), 
        .ZN(DP_mult_208_n463) );
  INV_X2 DP_mult_208_U1774 ( .A(DP_mult_208_n2238), .ZN(DP_mult_208_n2236) );
  INV_X2 DP_mult_208_U1773 ( .A(DP_mult_208_n2248), .ZN(DP_mult_208_n2246) );
  INV_X2 DP_mult_208_U1772 ( .A(DP_mult_208_n2253), .ZN(DP_mult_208_n2251) );
  INV_X2 DP_mult_208_U1771 ( .A(DP_mult_208_n2112), .ZN(DP_mult_208_n2210) );
  OR2_X1 DP_mult_208_U1770 ( .A1(DP_mult_208_n681), .A2(DP_mult_208_n684), 
        .ZN(DP_mult_208_n2135) );
  OR2_X1 DP_mult_208_U1769 ( .A1(DP_mult_208_n1143), .A2(DP_mult_208_n1150), 
        .ZN(DP_mult_208_n2121) );
  NOR2_X2 DP_mult_208_U1768 ( .A1(DP_mult_208_n727), .A2(DP_mult_208_n736), 
        .ZN(DP_mult_208_n428) );
  INV_X1 DP_mult_208_U1767 ( .A(DP_mult_208_n2142), .ZN(DP_mult_208_n2184) );
  AOI21_X1 DP_mult_208_U1766 ( .B1(DP_mult_208_n2166), .B2(DP_mult_208_n2010), 
        .A(DP_mult_208_n2078), .ZN(DP_mult_208_n2118) );
  INV_X1 DP_mult_208_U1765 ( .A(DP_mult_208_n2254), .ZN(DP_mult_208_n2249) );
  INV_X2 DP_mult_208_U1764 ( .A(DP_mult_208_n2114), .ZN(DP_mult_208_n536) );
  NOR2_X1 DP_mult_208_U1763 ( .A1(DP_mult_208_n495), .A2(DP_mult_208_n502), 
        .ZN(DP_mult_208_n489) );
  INV_X1 DP_mult_208_U1762 ( .A(DP_mult_208_n491), .ZN(DP_mult_208_n2116) );
  NAND3_X1 DP_mult_208_U1761 ( .A1(DP_mult_208_n2156), .A2(DP_mult_208_n2157), 
        .A3(DP_mult_208_n2158), .ZN(DP_mult_208_n2115) );
  OAI21_X1 DP_mult_208_U1760 ( .B1(DP_mult_208_n566), .B2(DP_mult_208_n538), 
        .A(DP_mult_208_n2046), .ZN(DP_mult_208_n2114) );
  INV_X2 DP_mult_208_U1759 ( .A(DP_mult_208_n2146), .ZN(DP_mult_208_n2192) );
  INV_X1 DP_mult_208_U1758 ( .A(DP_mult_208_n507), .ZN(DP_mult_208_n2113) );
  CLKBUF_X1 DP_mult_208_U1757 ( .A(DP_mult_208_n535), .Z(DP_mult_208_n2111) );
  OAI21_X1 DP_mult_208_U1756 ( .B1(DP_mult_208_n1933), .B2(DP_mult_208_n521), 
        .A(DP_mult_208_n514), .ZN(DP_mult_208_n2110) );
  INV_X2 DP_mult_208_U1755 ( .A(DP_mult_208_n2245), .ZN(DP_mult_208_n2241) );
  INV_X2 DP_mult_208_U1754 ( .A(DP_mult_208_n2229), .ZN(DP_mult_208_n2226) );
  INV_X1 DP_mult_208_U1753 ( .A(DP_mult_208_n2016), .ZN(DP_mult_208_n2201) );
  INV_X1 DP_mult_208_U1752 ( .A(DP_mult_208_n2143), .ZN(DP_mult_208_n2189) );
  NOR2_X1 DP_mult_208_U1751 ( .A1(DP_mult_208_n505), .A2(DP_mult_208_n452), 
        .ZN(DP_mult_208_n450) );
  NAND2_X1 DP_mult_208_U1750 ( .A1(DP_mult_208_n2106), .A2(DP_mult_208_n2107), 
        .ZN(DP_mult_208_n1372) );
  OR2_X1 DP_mult_208_U1749 ( .A1(DP_mult_208_n1667), .A2(DP_mult_208_n2035), 
        .ZN(DP_mult_208_n2107) );
  OR2_X1 DP_mult_208_U1748 ( .A1(DP_mult_208_n2191), .A2(DP_mult_208_n1668), 
        .ZN(DP_mult_208_n2106) );
  NAND3_X1 DP_mult_208_U1747 ( .A1(DP_mult_208_n2103), .A2(DP_mult_208_n2104), 
        .A3(DP_mult_208_n2105), .ZN(DP_mult_208_n972) );
  NAND2_X1 DP_mult_208_U1746 ( .A1(DP_mult_208_n994), .A2(DP_mult_208_n1217), 
        .ZN(DP_mult_208_n2105) );
  NAND2_X1 DP_mult_208_U1745 ( .A1(DP_mult_208_n996), .A2(DP_mult_208_n1217), 
        .ZN(DP_mult_208_n2104) );
  NAND2_X1 DP_mult_208_U1744 ( .A1(DP_mult_208_n996), .A2(DP_mult_208_n994), 
        .ZN(DP_mult_208_n2103) );
  XOR2_X1 DP_mult_208_U1743 ( .A(DP_mult_208_n2055), .B(DP_mult_208_n2102), 
        .Z(DP_mult_208_n973) );
  XOR2_X1 DP_mult_208_U1742 ( .A(DP_mult_208_n994), .B(DP_mult_208_n1217), .Z(
        DP_mult_208_n2102) );
  INV_X2 DP_mult_208_U1741 ( .A(DP_mult_208_n2159), .ZN(DP_mult_208_n2200) );
  OR2_X1 DP_mult_208_U1740 ( .A1(DP_mult_208_n919), .A2(DP_mult_208_n940), 
        .ZN(DP_mult_208_n2099) );
  AND2_X1 DP_mult_208_U1739 ( .A1(DP_mult_208_n1810), .A2(DP_mult_208_n265), 
        .ZN(DP_mult_208_n2098) );
  AND2_X1 DP_mult_208_U1738 ( .A1(DP_mult_208_n1810), .A2(DP_mult_208_n265), 
        .ZN(DP_mult_208_n2097) );
  OAI21_X1 DP_mult_208_U1737 ( .B1(DP_mult_208_n503), .B2(DP_mult_208_n2063), 
        .A(DP_mult_208_n496), .ZN(DP_mult_208_n2096) );
  NAND3_X1 DP_mult_208_U1736 ( .A1(DP_mult_208_n2093), .A2(DP_mult_208_n2094), 
        .A3(DP_mult_208_n2095), .ZN(DP_mult_208_n862) );
  NAND2_X1 DP_mult_208_U1735 ( .A1(DP_mult_208_n873), .A2(DP_mult_208_n888), 
        .ZN(DP_mult_208_n2095) );
  NAND2_X1 DP_mult_208_U1734 ( .A1(DP_mult_208_n886), .A2(DP_mult_208_n888), 
        .ZN(DP_mult_208_n2094) );
  NAND2_X1 DP_mult_208_U1733 ( .A1(DP_mult_208_n886), .A2(DP_mult_208_n873), 
        .ZN(DP_mult_208_n2093) );
  XOR2_X1 DP_mult_208_U1732 ( .A(DP_mult_208_n886), .B(DP_mult_208_n2092), .Z(
        DP_mult_208_n863) );
  XOR2_X1 DP_mult_208_U1731 ( .A(DP_mult_208_n873), .B(DP_mult_208_n888), .Z(
        DP_mult_208_n2092) );
  NOR2_X1 DP_mult_208_U1730 ( .A1(DP_mult_208_n941), .A2(DP_mult_208_n962), 
        .ZN(DP_mult_208_n547) );
  NOR2_X1 DP_mult_208_U1729 ( .A1(DP_mult_208_n919), .A2(DP_mult_208_n940), 
        .ZN(DP_mult_208_n542) );
  AOI21_X1 DP_mult_208_U1728 ( .B1(DP_mult_208_n1956), .B2(DP_mult_208_n1961), 
        .A(DP_mult_208_n568), .ZN(DP_mult_208_n2090) );
  AOI21_X1 DP_mult_208_U1727 ( .B1(DP_mult_208_n1956), .B2(DP_mult_208_n1961), 
        .A(DP_mult_208_n568), .ZN(DP_mult_208_n2091) );
  INV_X1 DP_mult_208_U1726 ( .A(DP_mult_208_n2146), .ZN(DP_mult_208_n2193) );
  INV_X1 DP_mult_208_U1725 ( .A(DP_mult_208_n2089), .ZN(DP_mult_208_n2140) );
  NAND3_X1 DP_mult_208_U1724 ( .A1(DP_mult_208_n2085), .A2(DP_mult_208_n2086), 
        .A3(DP_mult_208_n2087), .ZN(DP_mult_208_n860) );
  NAND2_X1 DP_mult_208_U1723 ( .A1(DP_mult_208_n865), .A2(DP_mult_208_n884), 
        .ZN(DP_mult_208_n2087) );
  NAND2_X1 DP_mult_208_U1722 ( .A1(DP_mult_208_n867), .A2(DP_mult_208_n884), 
        .ZN(DP_mult_208_n2086) );
  NAND2_X1 DP_mult_208_U1721 ( .A1(DP_mult_208_n867), .A2(DP_mult_208_n865), 
        .ZN(DP_mult_208_n2085) );
  XOR2_X1 DP_mult_208_U1720 ( .A(DP_mult_208_n2084), .B(DP_mult_208_n884), .Z(
        DP_mult_208_n861) );
  XOR2_X1 DP_mult_208_U1719 ( .A(DP_mult_208_n867), .B(DP_mult_208_n865), .Z(
        DP_mult_208_n2084) );
  NAND2_X1 DP_mult_208_U1718 ( .A1(DP_mult_208_n908), .A2(DP_mult_208_n895), 
        .ZN(DP_mult_208_n2083) );
  NAND2_X1 DP_mult_208_U1717 ( .A1(DP_mult_208_n891), .A2(DP_mult_208_n895), 
        .ZN(DP_mult_208_n2082) );
  NAND2_X1 DP_mult_208_U1716 ( .A1(DP_mult_208_n891), .A2(DP_mult_208_n908), 
        .ZN(DP_mult_208_n2081) );
  XOR2_X1 DP_mult_208_U1715 ( .A(DP_mult_208_n2080), .B(DP_mult_208_n895), .Z(
        DP_mult_208_n885) );
  XOR2_X1 DP_mult_208_U1714 ( .A(DP_mult_208_n891), .B(DP_mult_208_n908), .Z(
        DP_mult_208_n2080) );
  CLKBUF_X1 DP_mult_208_U1713 ( .A(DP_mult_208_n2110), .Z(DP_mult_208_n2078)
         );
  XOR2_X1 DP_mult_208_U1712 ( .A(DP_mult_208_n1216), .B(DP_mult_208_n1238), 
        .Z(DP_mult_208_n961) );
  INV_X2 DP_mult_208_U1711 ( .A(DP_mult_208_n2221), .ZN(DP_mult_208_n2217) );
  INV_X2 DP_mult_208_U1710 ( .A(DP_mult_208_n2053), .ZN(DP_mult_208_n2198) );
  NAND3_X1 DP_mult_208_U1709 ( .A1(DP_mult_208_n2074), .A2(DP_mult_208_n2075), 
        .A3(DP_mult_208_n2076), .ZN(DP_mult_208_n954) );
  NAND2_X1 DP_mult_208_U1708 ( .A1(DP_mult_208_n1304), .A2(DP_mult_208_n1414), 
        .ZN(DP_mult_208_n2076) );
  NAND2_X1 DP_mult_208_U1707 ( .A1(DP_mult_208_n1282), .A2(DP_mult_208_n1414), 
        .ZN(DP_mult_208_n2075) );
  NAND2_X1 DP_mult_208_U1706 ( .A1(DP_mult_208_n1282), .A2(DP_mult_208_n1304), 
        .ZN(DP_mult_208_n2074) );
  XOR2_X1 DP_mult_208_U1705 ( .A(DP_mult_208_n2073), .B(DP_mult_208_n2014), 
        .Z(DP_mult_208_n955) );
  XOR2_X1 DP_mult_208_U1704 ( .A(DP_mult_208_n1304), .B(DP_mult_208_n1414), 
        .Z(DP_mult_208_n2073) );
  INV_X2 DP_mult_208_U1703 ( .A(DP_mult_208_n2208), .ZN(DP_mult_208_n2207) );
  INV_X2 DP_mult_208_U1702 ( .A(DP_mult_208_n2147), .ZN(DP_mult_208_n2190) );
  INV_X2 DP_mult_208_U1701 ( .A(DP_mult_208_n2239), .ZN(DP_mult_208_n2235) );
  INV_X2 DP_mult_208_U1700 ( .A(DP_mult_208_n2144), .ZN(DP_mult_208_n2182) );
  INV_X2 DP_mult_208_U1699 ( .A(DP_mult_208_n2139), .ZN(DP_mult_208_n2212) );
  INV_X1 DP_mult_208_U1698 ( .A(DP_mult_208_n2072), .ZN(DP_mult_208_n2139) );
  XOR2_X1 DP_mult_208_U1697 ( .A(DP_coeffs_ff_int[61]), .B(DP_mult_208_n2244), 
        .Z(DP_mult_208_n2141) );
  INV_X2 DP_mult_208_U1696 ( .A(DP_mult_208_n2117), .ZN(DP_mult_208_n2205) );
  OAI22_X1 DP_mult_208_U1695 ( .A1(DP_mult_208_n2193), .A2(DP_mult_208_n1683), 
        .B1(DP_mult_208_n1682), .B2(DP_mult_208_n2050), .ZN(DP_mult_208_n2069)
         );
  INV_X1 DP_mult_208_U1694 ( .A(DP_mult_208_n2138), .ZN(DP_mult_208_n2199) );
  NOR2_X1 DP_mult_208_U1693 ( .A1(DP_mult_208_n896), .A2(DP_mult_208_n877), 
        .ZN(DP_mult_208_n531) );
  NOR2_X1 DP_mult_208_U1692 ( .A1(DP_mult_208_n877), .A2(DP_mult_208_n896), 
        .ZN(DP_mult_208_n2067) );
  INV_X1 DP_mult_208_U1691 ( .A(DP_mult_208_n2088), .ZN(DP_mult_208_n2176) );
  NOR2_X1 DP_mult_208_U1690 ( .A1(DP_mult_208_n805), .A2(DP_mult_208_n820), 
        .ZN(DP_mult_208_n495) );
  INV_X1 DP_mult_208_U1689 ( .A(DP_mult_208_n2224), .ZN(DP_mult_208_n2064) );
  INV_X1 DP_mult_208_U1688 ( .A(DP_mult_208_n2225), .ZN(DP_mult_208_n2065) );
  NOR2_X1 DP_mult_208_U1687 ( .A1(DP_mult_208_n805), .A2(DP_mult_208_n820), 
        .ZN(DP_mult_208_n2063) );
  INV_X1 DP_mult_208_U1686 ( .A(DP_mult_208_n2197), .ZN(DP_mult_208_n2062) );
  INV_X1 DP_mult_208_U1685 ( .A(DP_mult_208_n2146), .ZN(DP_mult_208_n2077) );
  OR2_X2 DP_mult_208_U1684 ( .A1(DP_mult_208_n775), .A2(DP_mult_208_n788), 
        .ZN(DP_mult_208_n2122) );
  XNOR2_X1 DP_mult_208_U1683 ( .A(DP_coeffs_ff_int[65]), .B(DP_mult_208_n2234), 
        .ZN(DP_mult_208_n1814) );
  XNOR2_X1 DP_mult_208_U1682 ( .A(DP_mult_208_n1415), .B(DP_mult_208_n1393), 
        .ZN(DP_mult_208_n2060) );
  XNOR2_X1 DP_mult_208_U1681 ( .A(DP_mult_208_n1979), .B(DP_mult_208_n2060), 
        .ZN(DP_mult_208_n975) );
  INV_X1 DP_mult_208_U1680 ( .A(DP_mult_208_n672), .ZN(DP_mult_208_n2058) );
  INV_X1 DP_mult_208_U1679 ( .A(DP_mult_208_n523), .ZN(DP_mult_208_n2057) );
  XOR2_X1 DP_mult_208_U1678 ( .A(DP_mult_208_n1240), .B(DP_mult_208_n1262), 
        .Z(DP_mult_208_n1001) );
  INV_X1 DP_mult_208_U1677 ( .A(DP_mult_208_n2101), .ZN(DP_mult_208_n2159) );
  INV_X1 DP_mult_208_U1676 ( .A(DP_mult_208_n2258), .ZN(DP_mult_208_n2255) );
  BUF_X4 DP_mult_208_U1675 ( .A(DP_mult_208_n277), .Z(DP_mult_208_n2100) );
  XOR2_X1 DP_mult_208_U1674 ( .A(DP_coeffs_ff_int[53]), .B(
        DP_coeffs_ff_int[54]), .Z(DP_mult_208_n2054) );
  OAI22_X1 DP_mult_208_U1673 ( .A1(DP_mult_208_n2182), .A2(DP_mult_208_n1530), 
        .B1(DP_mult_208_n1529), .B2(DP_mult_208_n2201), .ZN(DP_mult_208_n1240)
         );
  INV_X1 DP_mult_208_U1672 ( .A(DP_mult_208_n2071), .ZN(DP_mult_208_n2175) );
  INV_X1 DP_mult_208_U1671 ( .A(DP_mult_208_n2068), .ZN(DP_mult_208_n2148) );
  AND2_X1 DP_mult_208_U1670 ( .A1(DP_mult_208_n1817), .A2(DP_mult_208_n1959), 
        .ZN(DP_mult_208_n2138) );
  AND2_X1 DP_mult_208_U1669 ( .A1(DP_mult_208_n1817), .A2(DP_mult_208_n1959), 
        .ZN(DP_mult_208_n2052) );
  AND2_X1 DP_mult_208_U1668 ( .A1(DP_mult_208_n1817), .A2(DP_mult_208_n1959), 
        .ZN(DP_mult_208_n2053) );
  AND2_X1 DP_mult_208_U1667 ( .A1(DP_mult_208_n1808), .A2(DP_mult_208_n1978), 
        .ZN(DP_mult_208_n2066) );
  XNOR2_X1 DP_mult_208_U1666 ( .A(DP_coeffs_ff_int[50]), .B(
        DP_coeffs_ff_int[49]), .ZN(DP_mult_208_n2101) );
  INV_X1 DP_mult_208_U1665 ( .A(DP_mult_208_n2016), .ZN(DP_mult_208_n2202) );
  AND2_X2 DP_mult_208_U1664 ( .A1(DP_mult_208_n1806), .A2(DP_mult_208_n2101), 
        .ZN(DP_mult_208_n2145) );
  XNOR2_X1 DP_mult_208_U1663 ( .A(DP_coeffs_ff_int[71]), .B(DP_mult_208_n2220), 
        .ZN(DP_mult_208_n1817) );
  INV_X2 DP_mult_208_U1662 ( .A(DP_mult_208_n2176), .ZN(DP_mult_208_n2056) );
  XNOR2_X1 DP_mult_208_U1661 ( .A(DP_coeffs_ff_int[65]), .B(
        DP_coeffs_ff_int[66]), .ZN(DP_mult_208_n2071) );
  INV_X2 DP_mult_208_U1660 ( .A(DP_mult_208_n2175), .ZN(DP_mult_208_n2050) );
  INV_X1 DP_mult_208_U1659 ( .A(DP_mult_208_n2175), .ZN(DP_mult_208_n2048) );
  INV_X1 DP_mult_208_U1658 ( .A(DP_mult_208_n2175), .ZN(DP_mult_208_n2049) );
  INV_X1 DP_mult_208_U1657 ( .A(DP_mult_208_n2097), .ZN(DP_mult_208_n2047) );
  AOI21_X1 DP_mult_208_U1656 ( .B1(DP_mult_208_n553), .B2(DP_mult_208_n540), 
        .A(DP_mult_208_n541), .ZN(DP_mult_208_n2046) );
  INV_X1 DP_mult_208_U1655 ( .A(DP_mult_208_n2144), .ZN(DP_mult_208_n2181) );
  INV_X1 DP_mult_208_U1654 ( .A(DP_mult_208_n2201), .ZN(DP_mult_208_n2045) );
  INV_X1 DP_mult_208_U1653 ( .A(DP_mult_208_n2144), .ZN(DP_mult_208_n2044) );
  NAND3_X1 DP_mult_208_U1652 ( .A1(DP_mult_208_n2041), .A2(DP_mult_208_n2042), 
        .A3(DP_mult_208_n2043), .ZN(DP_mult_208_n796) );
  NAND2_X1 DP_mult_208_U1651 ( .A1(DP_mult_208_n1274), .A2(DP_mult_208_n1296), 
        .ZN(DP_mult_208_n2043) );
  NAND2_X1 DP_mult_208_U1650 ( .A1(DP_mult_208_n818), .A2(DP_mult_208_n1296), 
        .ZN(DP_mult_208_n2042) );
  NAND2_X1 DP_mult_208_U1649 ( .A1(DP_mult_208_n818), .A2(DP_mult_208_n1274), 
        .ZN(DP_mult_208_n2041) );
  XOR2_X1 DP_mult_208_U1648 ( .A(DP_mult_208_n818), .B(DP_mult_208_n2040), .Z(
        DP_mult_208_n797) );
  XOR2_X1 DP_mult_208_U1647 ( .A(DP_mult_208_n1274), .B(DP_mult_208_n1296), 
        .Z(DP_mult_208_n2040) );
  INV_X1 DP_mult_208_U1646 ( .A(DP_mult_208_n2070), .ZN(DP_mult_208_n2117) );
  OR2_X2 DP_mult_208_U1645 ( .A1(DP_mult_208_n2141), .A2(DP_mult_208_n2112), 
        .ZN(DP_mult_208_n2089) );
  OR2_X2 DP_mult_208_U1644 ( .A1(DP_mult_208_n2141), .A2(DP_mult_208_n1994), 
        .ZN(DP_mult_208_n2079) );
  INV_X1 DP_mult_208_U1643 ( .A(DP_mult_208_n1994), .ZN(DP_mult_208_n2211) );
  XNOR2_X1 DP_mult_208_U1642 ( .A(DP_coeffs_ff_int[69]), .B(
        DP_coeffs_ff_int[70]), .ZN(DP_mult_208_n2039) );
  XNOR2_X1 DP_mult_208_U1641 ( .A(DP_coeffs_ff_int[68]), .B(
        DP_coeffs_ff_int[67]), .ZN(DP_mult_208_n2072) );
  AND2_X2 DP_mult_208_U1640 ( .A1(DP_mult_208_n1811), .A2(DP_mult_208_n2068), 
        .ZN(DP_mult_208_n2143) );
  INV_X1 DP_mult_208_U1639 ( .A(DP_mult_208_n2148), .ZN(DP_mult_208_n2209) );
  INV_X2 DP_mult_208_U1638 ( .A(DP_mult_208_n2148), .ZN(DP_mult_208_n2038) );
  XNOR2_X1 DP_mult_208_U1637 ( .A(DP_coeffs_ff_int[57]), .B(
        DP_coeffs_ff_int[58]), .ZN(DP_mult_208_n265) );
  INV_X1 DP_mult_208_U1636 ( .A(DP_mult_208_n2117), .ZN(DP_mult_208_n2037) );
  XNOR2_X1 DP_mult_208_U1635 ( .A(DP_coeffs_ff_int[51]), .B(DP_mult_208_n2267), 
        .ZN(DP_mult_208_n1807) );
  OAI22_X1 DP_mult_208_U1634 ( .A1(DP_mult_208_n2196), .A2(DP_mult_208_n1733), 
        .B1(DP_mult_208_n1732), .B2(DP_mult_208_n2011), .ZN(DP_mult_208_n2036)
         );
  NAND3_X1 DP_mult_208_U1633 ( .A1(DP_mult_208_n2032), .A2(DP_mult_208_n2033), 
        .A3(DP_mult_208_n2034), .ZN(DP_mult_208_n958) );
  NAND2_X1 DP_mult_208_U1632 ( .A1(DP_mult_208_n1182), .A2(DP_mult_208_n1260), 
        .ZN(DP_mult_208_n2034) );
  NAND2_X1 DP_mult_208_U1631 ( .A1(DP_mult_208_n1348), .A2(DP_mult_208_n1182), 
        .ZN(DP_mult_208_n2033) );
  NAND2_X1 DP_mult_208_U1630 ( .A1(DP_mult_208_n1260), .A2(DP_mult_208_n1348), 
        .ZN(DP_mult_208_n2032) );
  XOR2_X1 DP_mult_208_U1629 ( .A(DP_mult_208_n2031), .B(DP_mult_208_n1348), 
        .Z(DP_mult_208_n959) );
  XOR2_X1 DP_mult_208_U1628 ( .A(DP_mult_208_n1182), .B(DP_mult_208_n1260), 
        .Z(DP_mult_208_n2031) );
  XNOR2_X1 DP_mult_208_U1627 ( .A(DP_coeffs_ff_int[63]), .B(DP_mult_208_n2239), 
        .ZN(DP_mult_208_n1813) );
  INV_X1 DP_mult_208_U1626 ( .A(DP_coeffs_ff_int[48]), .ZN(DP_mult_208_n2269)
         );
  INV_X2 DP_mult_208_U1625 ( .A(DP_mult_208_n2098), .ZN(DP_mult_208_n2187) );
  INV_X1 DP_mult_208_U1624 ( .A(DP_mult_208_n2264), .ZN(DP_mult_208_n2260) );
  INV_X2 DP_mult_208_U1623 ( .A(DP_mult_208_n1934), .ZN(DP_mult_208_n2232) );
  XNOR2_X1 DP_mult_208_U1622 ( .A(DP_coeffs_ff_int[53]), .B(DP_mult_208_n2263), 
        .ZN(DP_mult_208_n1808) );
  NAND3_X1 DP_mult_208_U1621 ( .A1(DP_mult_208_n2028), .A2(DP_mult_208_n2029), 
        .A3(DP_mult_208_n2030), .ZN(DP_mult_208_n918) );
  NAND2_X1 DP_mult_208_U1620 ( .A1(DP_mult_208_n923), .A2(DP_mult_208_n921), 
        .ZN(DP_mult_208_n2030) );
  NAND2_X1 DP_mult_208_U1619 ( .A1(DP_mult_208_n942), .A2(DP_mult_208_n921), 
        .ZN(DP_mult_208_n2029) );
  NAND2_X1 DP_mult_208_U1618 ( .A1(DP_mult_208_n942), .A2(DP_mult_208_n923), 
        .ZN(DP_mult_208_n2028) );
  NAND3_X1 DP_mult_208_U1617 ( .A1(DP_mult_208_n2025), .A2(DP_mult_208_n2026), 
        .A3(DP_mult_208_n2027), .ZN(DP_mult_208_n920) );
  NAND2_X1 DP_mult_208_U1616 ( .A1(DP_mult_208_n927), .A2(DP_mult_208_n944), 
        .ZN(DP_mult_208_n2027) );
  NAND2_X1 DP_mult_208_U1615 ( .A1(DP_mult_208_n944), .A2(DP_mult_208_n925), 
        .ZN(DP_mult_208_n2026) );
  NAND2_X1 DP_mult_208_U1614 ( .A1(DP_mult_208_n925), .A2(DP_mult_208_n927), 
        .ZN(DP_mult_208_n2025) );
  AND2_X2 DP_mult_208_U1613 ( .A1(DP_mult_208_n1809), .A2(DP_mult_208_n2070), 
        .ZN(DP_mult_208_n2142) );
  NAND2_X2 DP_mult_208_U1612 ( .A1(DP_mult_208_n1808), .A2(DP_mult_208_n1978), 
        .ZN(DP_mult_208_n2024) );
  NAND2_X1 DP_mult_208_U1611 ( .A1(DP_mult_208_n1808), .A2(DP_mult_208_n1978), 
        .ZN(DP_mult_208_n2023) );
  XNOR2_X1 DP_mult_208_U1610 ( .A(DP_mult_208_n942), .B(DP_mult_208_n923), 
        .ZN(DP_mult_208_n2022) );
  XNOR2_X1 DP_mult_208_U1609 ( .A(DP_mult_208_n2022), .B(DP_mult_208_n921), 
        .ZN(DP_mult_208_n919) );
  XNOR2_X1 DP_mult_208_U1608 ( .A(DP_mult_208_n925), .B(DP_mult_208_n927), 
        .ZN(DP_mult_208_n2021) );
  XNOR2_X1 DP_mult_208_U1607 ( .A(DP_mult_208_n2021), .B(DP_mult_208_n944), 
        .ZN(DP_mult_208_n921) );
  BUF_X4 DP_mult_208_U1606 ( .A(DP_coeffs_ff_int[48]), .Z(DP_mult_208_n2020)
         );
  INV_X1 DP_mult_208_U1605 ( .A(DP_mult_208_n1977), .ZN(DP_mult_208_n2194) );
  INV_X1 DP_mult_208_U1604 ( .A(DP_mult_208_n1936), .ZN(DP_mult_208_n2154) );
  XNOR2_X1 DP_mult_208_U1603 ( .A(DP_coeffs_ff_int[59]), .B(DP_mult_208_n2248), 
        .ZN(DP_mult_208_n1811) );
  OR2_X1 DP_mult_208_U1602 ( .A1(DP_mult_208_n839), .A2(DP_mult_208_n856), 
        .ZN(DP_mult_208_n2019) );
  INV_X2 DP_mult_208_U1601 ( .A(DP_mult_208_n2139), .ZN(DP_mult_208_n2213) );
  INV_X1 DP_mult_208_U1600 ( .A(DP_mult_208_n1977), .ZN(DP_mult_208_n2195) );
  INV_X1 DP_mult_208_U1599 ( .A(DP_mult_208_n1977), .ZN(DP_mult_208_n2017) );
  INV_X1 DP_mult_208_U1598 ( .A(DP_mult_208_n1977), .ZN(DP_mult_208_n2018) );
  XOR2_X1 DP_mult_208_U1597 ( .A(DP_coeffs_ff_int[51]), .B(
        DP_coeffs_ff_int[52]), .Z(DP_mult_208_n2016) );
  CLKBUF_X1 DP_mult_208_U1596 ( .A(DP_mult_208_n520), .Z(DP_mult_208_n2015) );
  BUF_X1 DP_mult_208_U1595 ( .A(DP_mult_208_n1282), .Z(DP_mult_208_n2014) );
  INV_X1 DP_mult_208_U1594 ( .A(DP_mult_208_n519), .ZN(DP_mult_208_n2013) );
  XNOR2_X1 DP_mult_208_U1593 ( .A(DP_coeffs_ff_int[55]), .B(
        DP_coeffs_ff_int[56]), .ZN(DP_mult_208_n2070) );
  BUF_X2 DP_mult_208_U1592 ( .A(DP_mult_208_n2070), .Z(DP_mult_208_n2012) );
  NOR2_X1 DP_mult_208_U1591 ( .A1(DP_mult_208_n839), .A2(DP_mult_208_n856), 
        .ZN(DP_mult_208_n513) );
  CLKBUF_X1 DP_mult_208_U1590 ( .A(DP_mult_208_n511), .Z(DP_mult_208_n2010) );
  AND2_X2 DP_mult_208_U1589 ( .A1(DP_mult_208_n1814), .A2(DP_mult_208_n2071), 
        .ZN(DP_mult_208_n2146) );
  INV_X1 DP_mult_208_U1588 ( .A(DP_mult_208_n555), .ZN(DP_mult_208_n2009) );
  XOR2_X1 DP_mult_208_U1587 ( .A(DP_coeffs_ff_int[67]), .B(
        DP_coeffs_ff_int[66]), .Z(DP_mult_208_n1815) );
  NAND3_X1 DP_mult_208_U1586 ( .A1(DP_mult_208_n2005), .A2(DP_mult_208_n2006), 
        .A3(DP_mult_208_n2007), .ZN(DP_mult_208_n994) );
  NAND2_X1 DP_mult_208_U1585 ( .A1(DP_mult_208_n1416), .A2(DP_mult_208_n1306), 
        .ZN(DP_mult_208_n2007) );
  NAND2_X1 DP_mult_208_U1584 ( .A1(DP_mult_208_n1328), .A2(DP_mult_208_n1306), 
        .ZN(DP_mult_208_n2006) );
  NAND2_X1 DP_mult_208_U1583 ( .A1(DP_mult_208_n1328), .A2(DP_mult_208_n1416), 
        .ZN(DP_mult_208_n2005) );
  XOR2_X1 DP_mult_208_U1582 ( .A(DP_mult_208_n1328), .B(DP_mult_208_n2004), 
        .Z(DP_mult_208_n995) );
  XOR2_X1 DP_mult_208_U1581 ( .A(DP_mult_208_n1306), .B(DP_mult_208_n1416), 
        .Z(DP_mult_208_n2004) );
  XNOR2_X1 DP_mult_208_U1580 ( .A(DP_coeffs_ff_int[59]), .B(
        DP_coeffs_ff_int[60]), .ZN(DP_mult_208_n2068) );
  BUF_X2 DP_mult_208_U1579 ( .A(DP_mult_208_n2068), .Z(DP_mult_208_n2003) );
  NAND3_X1 DP_mult_208_U1578 ( .A1(DP_mult_208_n2000), .A2(DP_mult_208_n2001), 
        .A3(DP_mult_208_n2002), .ZN(DP_mult_208_n1038) );
  NAND2_X1 DP_mult_208_U1577 ( .A1(DP_mult_208_n1056), .A2(DP_mult_208_n1043), 
        .ZN(DP_mult_208_n2002) );
  NAND2_X1 DP_mult_208_U1576 ( .A1(DP_mult_208_n1041), .A2(DP_mult_208_n1043), 
        .ZN(DP_mult_208_n2001) );
  NAND2_X1 DP_mult_208_U1575 ( .A1(DP_mult_208_n1041), .A2(DP_mult_208_n1056), 
        .ZN(DP_mult_208_n2000) );
  XOR2_X1 DP_mult_208_U1574 ( .A(DP_mult_208_n1041), .B(DP_mult_208_n1999), 
        .Z(DP_mult_208_n1039) );
  XOR2_X1 DP_mult_208_U1573 ( .A(DP_mult_208_n1056), .B(DP_mult_208_n1043), 
        .Z(DP_mult_208_n1999) );
  INV_X2 DP_mult_208_U1572 ( .A(DP_mult_208_n2259), .ZN(DP_mult_208_n2257) );
  NAND3_X1 DP_mult_208_U1571 ( .A1(DP_mult_208_n1996), .A2(DP_mult_208_n1997), 
        .A3(DP_mult_208_n1998), .ZN(DP_mult_208_n1032) );
  NAND2_X1 DP_mult_208_U1570 ( .A1(DP_mult_208_n1330), .A2(DP_mult_208_n1463), 
        .ZN(DP_mult_208_n1998) );
  NAND2_X1 DP_mult_208_U1569 ( .A1(DP_mult_208_n1463), .A2(DP_mult_208_n1396), 
        .ZN(DP_mult_208_n1997) );
  NAND2_X1 DP_mult_208_U1568 ( .A1(DP_mult_208_n1330), .A2(DP_mult_208_n1396), 
        .ZN(DP_mult_208_n1996) );
  XOR2_X1 DP_mult_208_U1567 ( .A(DP_mult_208_n1995), .B(DP_mult_208_n1396), 
        .Z(DP_mult_208_n1033) );
  XOR2_X1 DP_mult_208_U1566 ( .A(DP_mult_208_n1330), .B(DP_mult_208_n1463), 
        .Z(DP_mult_208_n1995) );
  XNOR2_X1 DP_mult_208_U1565 ( .A(DP_coeffs_ff_int[61]), .B(DP_mult_208_n2238), 
        .ZN(DP_mult_208_n2112) );
  XNOR2_X1 DP_mult_208_U1564 ( .A(DP_coeffs_ff_int[61]), .B(DP_mult_208_n2238), 
        .ZN(DP_mult_208_n1994) );
  INV_X1 DP_mult_208_U1563 ( .A(DP_mult_208_n2142), .ZN(DP_mult_208_n2119) );
  AND2_X1 DP_mult_208_U1562 ( .A1(DP_mult_208_n672), .A2(DP_mult_208_n2111), 
        .ZN(DP_mult_208_n1993) );
  XNOR2_X1 DP_mult_208_U1561 ( .A(DP_mult_208_n536), .B(DP_mult_208_n1993), 
        .ZN(DP_pipe0_coeff_pipe02[3]) );
  AND2_X1 DP_mult_208_U1560 ( .A1(DP_mult_208_n675), .A2(DP_mult_208_n559), 
        .ZN(DP_mult_208_n1992) );
  XNOR2_X1 DP_mult_208_U1559 ( .A(DP_mult_208_n560), .B(DP_mult_208_n1992), 
        .ZN(DP_pipe0_coeff_pipe02[0]) );
  AND2_X1 DP_mult_208_U1558 ( .A1(DP_mult_208_n2099), .A2(DP_mult_208_n543), 
        .ZN(DP_mult_208_n1991) );
  XNOR2_X1 DP_mult_208_U1557 ( .A(DP_mult_208_n544), .B(DP_mult_208_n1991), 
        .ZN(DP_pipe0_coeff_pipe02[2]) );
  AND2_X1 DP_mult_208_U1556 ( .A1(DP_mult_208_n1948), .A2(DP_mult_208_n674), 
        .ZN(DP_mult_208_n1990) );
  XNOR2_X1 DP_mult_208_U1555 ( .A(DP_mult_208_n551), .B(DP_mult_208_n1990), 
        .ZN(DP_pipe0_coeff_pipe02[1]) );
  OR2_X1 DP_mult_208_U1554 ( .A1(DP_mult_208_n1123), .A2(DP_mult_208_n1132), 
        .ZN(DP_mult_208_n1989) );
  OR2_X1 DP_mult_208_U1553 ( .A1(DP_mult_208_n1151), .A2(DP_mult_208_n1158), 
        .ZN(DP_mult_208_n1988) );
  AND2_X1 DP_mult_208_U1552 ( .A1(DP_mult_208_n1021), .A2(DP_mult_208_n1038), 
        .ZN(DP_mult_208_n1987) );
  AND2_X1 DP_mult_208_U1551 ( .A1(DP_mult_208_n1111), .A2(DP_mult_208_n1122), 
        .ZN(DP_mult_208_n1986) );
  AND2_X1 DP_mult_208_U1550 ( .A1(DP_mult_208_n1055), .A2(DP_mult_208_n1070), 
        .ZN(DP_mult_208_n1985) );
  AND2_X1 DP_mult_208_U1549 ( .A1(DP_mult_208_n1133), .A2(DP_mult_208_n1142), 
        .ZN(DP_mult_208_n1984) );
  AND2_X1 DP_mult_208_U1548 ( .A1(DP_mult_208_n1179), .A2(DP_mult_208_n1433), 
        .ZN(DP_mult_208_n1983) );
  OR2_X1 DP_mult_208_U1547 ( .A1(DP_mult_208_n1039), .A2(DP_mult_208_n1054), 
        .ZN(DP_mult_208_n1982) );
  AND2_X1 DP_mult_208_U1546 ( .A1(DP_mult_208_n1457), .A2(DP_mult_208_n1480), 
        .ZN(DP_mult_208_n1981) );
  AND2_X1 DP_mult_208_U1545 ( .A1(DP_mult_208_n1216), .A2(DP_mult_208_n1238), 
        .ZN(DP_mult_208_n1980) );
  AND2_X1 DP_mult_208_U1544 ( .A1(DP_mult_208_n1240), .A2(DP_mult_208_n1262), 
        .ZN(DP_mult_208_n1979) );
  XNOR2_X1 DP_mult_208_U1543 ( .A(DP_coeffs_ff_int[53]), .B(
        DP_coeffs_ff_int[54]), .ZN(DP_mult_208_n1978) );
  BUF_X1 DP_mult_208_U1542 ( .A(DP_mult_208_n2088), .Z(DP_mult_208_n2035) );
  AND2_X1 DP_mult_208_U1541 ( .A1(DP_mult_208_n1815), .A2(DP_mult_208_n2072), 
        .ZN(DP_mult_208_n1977) );
  AND2_X1 DP_mult_208_U1540 ( .A1(DP_mult_208_n1151), .A2(DP_mult_208_n1158), 
        .ZN(DP_mult_208_n1976) );
  AND2_X1 DP_mult_208_U1539 ( .A1(DP_mult_208_n1123), .A2(DP_mult_208_n1132), 
        .ZN(DP_mult_208_n1975) );
  AND2_X1 DP_mult_208_U1538 ( .A1(DP_mult_208_n1143), .A2(DP_mult_208_n1150), 
        .ZN(DP_mult_208_n1974) );
  OR2_X1 DP_mult_208_U1537 ( .A1(DP_mult_208_n1179), .A2(DP_mult_208_n1433), 
        .ZN(DP_mult_208_n1973) );
  OR2_X1 DP_mult_208_U1536 ( .A1(DP_mult_208_n1457), .A2(DP_mult_208_n1480), 
        .ZN(DP_mult_208_n1972) );
  AND2_X1 DP_mult_208_U1535 ( .A1(DP_mult_208_n1039), .A2(DP_mult_208_n1054), 
        .ZN(DP_mult_208_n1971) );
  AND2_X1 DP_mult_208_U1534 ( .A1(DP_mult_208_n1193), .A2(DP_mult_208_n1481), 
        .ZN(DP_mult_208_n1970) );
  INV_X1 DP_mult_208_U1533 ( .A(DP_mult_208_n2061), .ZN(DP_mult_208_n474) );
  AND2_X1 DP_mult_208_U1532 ( .A1(DP_mult_208_n775), .A2(DP_mult_208_n788), 
        .ZN(DP_mult_208_n2061) );
  NOR2_X1 DP_mult_208_U1531 ( .A1(DP_mult_208_n821), .A2(DP_mult_208_n838), 
        .ZN(DP_mult_208_n502) );
  NAND2_X1 DP_mult_208_U1530 ( .A1(DP_mult_208_n2127), .A2(DP_mult_208_n2129), 
        .ZN(DP_mult_208_n402) );
  NOR2_X1 DP_mult_208_U1529 ( .A1(DP_mult_208_n435), .A2(DP_mult_208_n428), 
        .ZN(DP_mult_208_n426) );
  NAND3_X1 DP_mult_208_U1528 ( .A1(DP_mult_208_n2081), .A2(DP_mult_208_n2082), 
        .A3(DP_mult_208_n2083), .ZN(DP_mult_208_n884) );
  INV_X1 DP_mult_208_U1527 ( .A(DP_mult_208_n2066), .ZN(DP_mult_208_n2183) );
  NOR2_X1 DP_mult_208_U1526 ( .A1(DP_mult_208_n1969), .A2(DP_mult_208_n568), 
        .ZN(DP_mult_208_n566) );
  AND2_X1 DP_mult_208_U1525 ( .A1(DP_mult_208_n581), .A2(DP_mult_208_n567), 
        .ZN(DP_mult_208_n1969) );
  XNOR2_X1 DP_mult_208_U1524 ( .A(DP_mult_208_n1326), .B(DP_mult_208_n1392), 
        .ZN(DP_mult_208_n1968) );
  XNOR2_X1 DP_mult_208_U1523 ( .A(DP_mult_208_n961), .B(DP_mult_208_n1968), 
        .ZN(DP_mult_208_n953) );
  AND2_X2 DP_mult_208_U1522 ( .A1(DP_mult_208_n1813), .A2(DP_mult_208_n2088), 
        .ZN(DP_mult_208_n2147) );
  INV_X1 DP_mult_208_U1521 ( .A(DP_mult_208_n2234), .ZN(DP_mult_208_n2233) );
  CLKBUF_X3 DP_mult_208_U1520 ( .A(DP_coeffs_ff_int[50]), .Z(DP_mult_208_n1967) );
  XNOR2_X1 DP_mult_208_U1519 ( .A(DP_pipe02[3]), .B(DP_mult_208_n1967), .ZN(
        DP_mult_208_n1966) );
  INV_X1 DP_mult_208_U1518 ( .A(DP_mult_208_n1963), .ZN(DP_mult_208_n1964) );
  INV_X1 DP_mult_208_U1517 ( .A(DP_mult_208_n2270), .ZN(DP_mult_208_n1963) );
  INV_X1 DP_mult_208_U1516 ( .A(DP_coeffs_ff_int[64]), .ZN(DP_mult_208_n2234)
         );
  INV_X1 DP_mult_208_U1515 ( .A(DP_mult_208_n2231), .ZN(DP_mult_208_n1962) );
  INV_X2 DP_mult_208_U1514 ( .A(DP_mult_208_n2147), .ZN(DP_mult_208_n2191) );
  INV_X2 DP_mult_208_U1513 ( .A(DP_mult_208_n2224), .ZN(DP_mult_208_n2222) );
  NOR2_X1 DP_mult_208_U1512 ( .A1(DP_mult_208_n571), .A2(DP_mult_208_n1952), 
        .ZN(DP_mult_208_n1961) );
  BUF_X1 DP_mult_208_U1511 ( .A(DP_mult_208_n251), .Z(DP_mult_208_n2214) );
  BUF_X2 DP_mult_208_U1510 ( .A(DP_mult_208_n2214), .Z(DP_mult_208_n1960) );
  CLKBUF_X1 DP_mult_208_U1509 ( .A(DP_mult_208_n2214), .Z(DP_mult_208_n1959)
         );
  NOR2_X1 DP_mult_208_U1508 ( .A1(DP_mult_208_n558), .A2(DP_mult_208_n563), 
        .ZN(DP_mult_208_n552) );
  INV_X1 DP_mult_208_U1507 ( .A(DP_mult_208_n2143), .ZN(DP_mult_208_n2109) );
  INV_X1 DP_mult_208_U1506 ( .A(DP_mult_208_n2143), .ZN(DP_mult_208_n2188) );
  XNOR2_X1 DP_mult_208_U1505 ( .A(DP_coeffs_ff_int[63]), .B(
        DP_coeffs_ff_int[64]), .ZN(DP_mult_208_n2088) );
  INV_X1 DP_mult_208_U1504 ( .A(DP_mult_208_n2176), .ZN(DP_mult_208_n1958) );
  XOR2_X1 DP_mult_208_U1503 ( .A(DP_coeffs_ff_int[49]), .B(
        DP_coeffs_ff_int[48]), .Z(DP_mult_208_n1806) );
  INV_X2 DP_mult_208_U1502 ( .A(DP_mult_208_n2264), .ZN(DP_mult_208_n2262) );
  XOR2_X1 DP_mult_208_U1501 ( .A(DP_coeffs_ff_int[57]), .B(
        DP_coeffs_ff_int[56]), .Z(DP_mult_208_n1810) );
  CLKBUF_X2 DP_mult_208_U1500 ( .A(DP_coeffs_ff_int[58]), .Z(DP_mult_208_n2008) );
  INV_X2 DP_mult_208_U1499 ( .A(DP_mult_208_n2142), .ZN(DP_mult_208_n2120) );
  NAND3_X1 DP_mult_208_U1498 ( .A1(DP_mult_208_n2093), .A2(DP_mult_208_n2094), 
        .A3(DP_mult_208_n2095), .ZN(DP_mult_208_n1957) );
  INV_X2 DP_mult_208_U1497 ( .A(DP_mult_208_n2142), .ZN(DP_mult_208_n2185) );
  INV_X1 DP_mult_208_U1496 ( .A(DP_mult_208_n1963), .ZN(DP_mult_208_n1965) );
  INV_X1 DP_mult_208_U1495 ( .A(DP_pipe02[0]), .ZN(DP_mult_208_n1955) );
  NOR2_X1 DP_mult_208_U1494 ( .A1(DP_mult_208_n963), .A2(DP_mult_208_n982), 
        .ZN(DP_mult_208_n558) );
  NOR2_X1 DP_mult_208_U1493 ( .A1(DP_mult_208_n963), .A2(DP_mult_208_n982), 
        .ZN(DP_mult_208_n1954) );
  INV_X2 DP_mult_208_U1492 ( .A(DP_mult_208_n2253), .ZN(DP_mult_208_n2250) );
  INV_X1 DP_mult_208_U1491 ( .A(DP_mult_208_n2246), .ZN(DP_mult_208_n1953) );
  NOR2_X1 DP_mult_208_U1490 ( .A1(DP_mult_208_n1003), .A2(DP_mult_208_n1020), 
        .ZN(DP_mult_208_n569) );
  NOR2_X1 DP_mult_208_U1489 ( .A1(DP_mult_208_n1003), .A2(DP_mult_208_n1020), 
        .ZN(DP_mult_208_n1951) );
  NOR2_X1 DP_mult_208_U1488 ( .A1(DP_mult_208_n1003), .A2(DP_mult_208_n1020), 
        .ZN(DP_mult_208_n1952) );
  INV_X1 DP_mult_208_U1487 ( .A(DP_mult_208_n2052), .ZN(DP_mult_208_n2059) );
  INV_X1 DP_mult_208_U1486 ( .A(DP_mult_208_n2052), .ZN(DP_mult_208_n1950) );
  CLKBUF_X1 DP_mult_208_U1485 ( .A(DP_mult_208_n547), .Z(DP_mult_208_n1949) );
  INV_X2 DP_mult_208_U1484 ( .A(DP_mult_208_n2230), .ZN(DP_mult_208_n2227) );
  INV_X1 DP_mult_208_U1483 ( .A(DP_mult_208_n2143), .ZN(DP_mult_208_n2108) );
  CLKBUF_X1 DP_mult_208_U1482 ( .A(DP_mult_208_n550), .Z(DP_mult_208_n1948) );
  OR2_X1 DP_mult_208_U1481 ( .A1(DP_mult_208_n1021), .A2(DP_mult_208_n1038), 
        .ZN(DP_mult_208_n1947) );
  BUF_X1 DP_mult_208_U1480 ( .A(DP_mult_208_n581), .Z(DP_mult_208_n1956) );
  INV_X1 DP_mult_208_U1479 ( .A(DP_mult_208_n2138), .ZN(DP_mult_208_n1946) );
  NAND3_X1 DP_mult_208_U1478 ( .A1(DP_mult_208_n1943), .A2(DP_mult_208_n1944), 
        .A3(DP_mult_208_n1945), .ZN(DP_mult_208_n928) );
  NAND2_X1 DP_mult_208_U1477 ( .A1(DP_mult_208_n954), .A2(DP_mult_208_n956), 
        .ZN(DP_mult_208_n1945) );
  NAND2_X1 DP_mult_208_U1476 ( .A1(DP_mult_208_n958), .A2(DP_mult_208_n956), 
        .ZN(DP_mult_208_n1944) );
  NAND2_X1 DP_mult_208_U1475 ( .A1(DP_mult_208_n958), .A2(DP_mult_208_n954), 
        .ZN(DP_mult_208_n1943) );
  XOR2_X1 DP_mult_208_U1474 ( .A(DP_mult_208_n1942), .B(DP_mult_208_n956), .Z(
        DP_mult_208_n929) );
  XOR2_X1 DP_mult_208_U1473 ( .A(DP_mult_208_n958), .B(DP_mult_208_n954), .Z(
        DP_mult_208_n1942) );
  NAND3_X1 DP_mult_208_U1472 ( .A1(DP_mult_208_n1939), .A2(DP_mult_208_n1940), 
        .A3(DP_mult_208_n1941), .ZN(DP_mult_208_n956) );
  NAND2_X1 DP_mult_208_U1471 ( .A1(DP_mult_208_n1370), .A2(DP_mult_208_n1436), 
        .ZN(DP_mult_208_n1941) );
  NAND2_X1 DP_mult_208_U1470 ( .A1(DP_mult_208_n1459), .A2(DP_mult_208_n1436), 
        .ZN(DP_mult_208_n1940) );
  NAND2_X1 DP_mult_208_U1469 ( .A1(DP_mult_208_n1459), .A2(DP_mult_208_n1370), 
        .ZN(DP_mult_208_n1939) );
  XOR2_X1 DP_mult_208_U1468 ( .A(DP_mult_208_n1938), .B(DP_mult_208_n1436), 
        .Z(DP_mult_208_n957) );
  XOR2_X1 DP_mult_208_U1467 ( .A(DP_mult_208_n1459), .B(DP_mult_208_n1370), 
        .Z(DP_mult_208_n1938) );
  CLKBUF_X3 DP_mult_208_U1466 ( .A(DP_mult_208_n2039), .Z(DP_mult_208_n2011)
         );
  CLKBUF_X3 DP_mult_208_U1465 ( .A(DP_mult_208_n1936), .Z(DP_mult_208_n1937)
         );
  XNOR2_X1 DP_mult_208_U1464 ( .A(DP_coeffs_ff_int[69]), .B(
        DP_coeffs_ff_int[70]), .ZN(DP_mult_208_n1936) );
  XNOR2_X1 DP_mult_208_U1463 ( .A(DP_coeffs_ff_int[51]), .B(
        DP_coeffs_ff_int[52]), .ZN(DP_mult_208_n1935) );
  XOR2_X1 DP_mult_208_U1462 ( .A(DP_pipe02[1]), .B(DP_mult_208_n2269), .Z(
        DP_mult_208_n1504) );
  INV_X1 DP_mult_208_U1461 ( .A(DP_coeffs_ff_int[64]), .ZN(DP_mult_208_n1934)
         );
  XOR2_X1 DP_mult_208_U1460 ( .A(DP_coeffs_ff_int[69]), .B(
        DP_coeffs_ff_int[68]), .Z(DP_mult_208_n1816) );
  INV_X1 DP_mult_208_U1459 ( .A(DP_mult_208_n2145), .ZN(DP_mult_208_n2179) );
  CLKBUF_X2 DP_mult_208_U1458 ( .A(DP_mult_208_n2101), .Z(DP_mult_208_n2051)
         );
  NOR2_X1 DP_mult_208_U1457 ( .A1(DP_mult_208_n839), .A2(DP_mult_208_n856), 
        .ZN(DP_mult_208_n1933) );
  BUF_X1 DP_mult_208_U1456 ( .A(DP_mult_208_n996), .Z(DP_mult_208_n2055) );
  NAND3_X1 DP_mult_208_U1455 ( .A1(DP_mult_208_n1930), .A2(DP_mult_208_n1931), 
        .A3(DP_mult_208_n1932), .ZN(DP_mult_208_n996) );
  NAND2_X1 DP_mult_208_U1454 ( .A1(DP_mult_208_n1372), .A2(DP_mult_208_n1438), 
        .ZN(DP_mult_208_n1932) );
  NAND2_X1 DP_mult_208_U1453 ( .A1(DP_mult_208_n1284), .A2(DP_mult_208_n1438), 
        .ZN(DP_mult_208_n1931) );
  NAND2_X1 DP_mult_208_U1452 ( .A1(DP_mult_208_n1284), .A2(DP_mult_208_n1372), 
        .ZN(DP_mult_208_n1930) );
  XOR2_X1 DP_mult_208_U1451 ( .A(DP_mult_208_n1929), .B(DP_mult_208_n1284), 
        .Z(DP_mult_208_n997) );
  XOR2_X1 DP_mult_208_U1450 ( .A(DP_mult_208_n1372), .B(DP_mult_208_n1438), 
        .Z(DP_mult_208_n1929) );
  INV_X2 DP_mult_208_U1449 ( .A(DP_mult_208_n2221), .ZN(DP_mult_208_n2218) );
  XOR2_X1 DP_mult_208_U1448 ( .A(DP_coeffs_ff_int[55]), .B(
        DP_coeffs_ff_int[54]), .Z(DP_mult_208_n1809) );
  HA_X1 DP_mult_208_U798 ( .A(DP_mult_208_n1456), .B(DP_mult_208_n1479), .CO(
        DP_mult_208_n1180), .S(DP_mult_208_n1181) );
  FA_X1 DP_mult_208_U797 ( .A(DP_mult_208_n1455), .B(DP_mult_208_n1478), .CI(
        DP_mult_208_n1180), .CO(DP_mult_208_n1178), .S(DP_mult_208_n1179) );
  HA_X1 DP_mult_208_U796 ( .A(DP_mult_208_n1432), .B(DP_mult_208_n1477), .CO(
        DP_mult_208_n1176), .S(DP_mult_208_n1177) );
  FA_X1 DP_mult_208_U795 ( .A(DP_mult_208_n1191), .B(DP_mult_208_n1454), .CI(
        DP_mult_208_n1177), .CO(DP_mult_208_n1174), .S(DP_mult_208_n1175) );
  FA_X1 DP_mult_208_U794 ( .A(DP_mult_208_n1476), .B(DP_mult_208_n1453), .CI(
        DP_mult_208_n1431), .CO(DP_mult_208_n1172), .S(DP_mult_208_n1173) );
  FA_X1 DP_mult_208_U793 ( .A(DP_mult_208_n1409), .B(DP_mult_208_n1176), .CI(
        DP_mult_208_n1173), .CO(DP_mult_208_n1170), .S(DP_mult_208_n1171) );
  HA_X1 DP_mult_208_U792 ( .A(DP_mult_208_n1408), .B(DP_mult_208_n1430), .CO(
        DP_mult_208_n1168), .S(DP_mult_208_n1169) );
  FA_X1 DP_mult_208_U791 ( .A(DP_mult_208_n1452), .B(DP_mult_208_n1475), .CI(
        DP_mult_208_n1190), .CO(DP_mult_208_n1166), .S(DP_mult_208_n1167) );
  FA_X1 DP_mult_208_U790 ( .A(DP_mult_208_n1172), .B(DP_mult_208_n1169), .CI(
        DP_mult_208_n1167), .CO(DP_mult_208_n1164), .S(DP_mult_208_n1165) );
  FA_X1 DP_mult_208_U789 ( .A(DP_mult_208_n1451), .B(DP_mult_208_n1474), .CI(
        DP_mult_208_n1407), .CO(DP_mult_208_n1162), .S(DP_mult_208_n1163) );
  FA_X1 DP_mult_208_U788 ( .A(DP_mult_208_n1168), .B(DP_mult_208_n1429), .CI(
        DP_mult_208_n1166), .CO(DP_mult_208_n1160), .S(DP_mult_208_n1161) );
  FA_X1 DP_mult_208_U787 ( .A(DP_mult_208_n1163), .B(DP_mult_208_n1385), .CI(
        DP_mult_208_n1164), .CO(DP_mult_208_n1158), .S(DP_mult_208_n1159) );
  HA_X1 DP_mult_208_U786 ( .A(DP_mult_208_n1384), .B(DP_mult_208_n1406), .CO(
        DP_mult_208_n1156), .S(DP_mult_208_n1157) );
  FA_X1 DP_mult_208_U785 ( .A(DP_mult_208_n1450), .B(DP_mult_208_n1428), .CI(
        DP_mult_208_n1189), .CO(DP_mult_208_n1154), .S(DP_mult_208_n1155) );
  FA_X1 DP_mult_208_U784 ( .A(DP_mult_208_n1157), .B(DP_mult_208_n1473), .CI(
        DP_mult_208_n1162), .CO(DP_mult_208_n1152), .S(DP_mult_208_n1153) );
  FA_X1 DP_mult_208_U783 ( .A(DP_mult_208_n1160), .B(DP_mult_208_n1155), .CI(
        DP_mult_208_n1153), .CO(DP_mult_208_n1150), .S(DP_mult_208_n1151) );
  FA_X1 DP_mult_208_U782 ( .A(DP_mult_208_n1383), .B(DP_mult_208_n1472), .CI(
        DP_mult_208_n1405), .CO(DP_mult_208_n1148), .S(DP_mult_208_n1149) );
  FA_X1 DP_mult_208_U781 ( .A(DP_mult_208_n1427), .B(DP_mult_208_n1449), .CI(
        DP_mult_208_n1156), .CO(DP_mult_208_n1146), .S(DP_mult_208_n1147) );
  FA_X1 DP_mult_208_U780 ( .A(DP_mult_208_n1361), .B(DP_mult_208_n1154), .CI(
        DP_mult_208_n1149), .CO(DP_mult_208_n1144), .S(DP_mult_208_n1145) );
  FA_X1 DP_mult_208_U779 ( .A(DP_mult_208_n1152), .B(DP_mult_208_n1147), .CI(
        DP_mult_208_n1145), .CO(DP_mult_208_n1142), .S(DP_mult_208_n1143) );
  HA_X1 DP_mult_208_U778 ( .A(DP_mult_208_n1360), .B(DP_mult_208_n1382), .CO(
        DP_mult_208_n1140), .S(DP_mult_208_n1141) );
  FA_X1 DP_mult_208_U777 ( .A(DP_mult_208_n1188), .B(DP_mult_208_n1426), .CI(
        DP_mult_208_n1471), .CO(DP_mult_208_n1138), .S(DP_mult_208_n1139) );
  FA_X1 DP_mult_208_U776 ( .A(DP_mult_208_n1404), .B(DP_mult_208_n1448), .CI(
        DP_mult_208_n1141), .CO(DP_mult_208_n1136), .S(DP_mult_208_n1137) );
  FA_X1 DP_mult_208_U775 ( .A(DP_mult_208_n1146), .B(DP_mult_208_n1148), .CI(
        DP_mult_208_n1139), .CO(DP_mult_208_n1134), .S(DP_mult_208_n1135) );
  FA_X1 DP_mult_208_U774 ( .A(DP_mult_208_n1144), .B(DP_mult_208_n1137), .CI(
        DP_mult_208_n1135), .CO(DP_mult_208_n1132), .S(DP_mult_208_n1133) );
  FA_X1 DP_mult_208_U773 ( .A(DP_mult_208_n1359), .B(DP_mult_208_n1470), .CI(
        DP_mult_208_n1381), .CO(DP_mult_208_n1130), .S(DP_mult_208_n1131) );
  FA_X1 DP_mult_208_U772 ( .A(DP_mult_208_n1403), .B(DP_mult_208_n1447), .CI(
        DP_mult_208_n1425), .CO(DP_mult_208_n1128), .S(DP_mult_208_n1129) );
  FA_X1 DP_mult_208_U771 ( .A(DP_mult_208_n1138), .B(DP_mult_208_n1140), .CI(
        DP_mult_208_n1337), .CO(DP_mult_208_n1126), .S(DP_mult_208_n1127) );
  FA_X1 DP_mult_208_U770 ( .A(DP_mult_208_n1131), .B(DP_mult_208_n1129), .CI(
        DP_mult_208_n1136), .CO(DP_mult_208_n1124), .S(DP_mult_208_n1125) );
  FA_X1 DP_mult_208_U769 ( .A(DP_mult_208_n1127), .B(DP_mult_208_n1134), .CI(
        DP_mult_208_n1125), .CO(DP_mult_208_n1122), .S(DP_mult_208_n1123) );
  HA_X1 DP_mult_208_U768 ( .A(DP_mult_208_n1336), .B(DP_mult_208_n1358), .CO(
        DP_mult_208_n1120), .S(DP_mult_208_n1121) );
  FA_X1 DP_mult_208_U767 ( .A(DP_mult_208_n1380), .B(DP_mult_208_n1402), .CI(
        DP_mult_208_n1187), .CO(DP_mult_208_n1118), .S(DP_mult_208_n1119) );
  FA_X1 DP_mult_208_U766 ( .A(DP_mult_208_n1424), .B(DP_mult_208_n1469), .CI(
        DP_mult_208_n1446), .CO(DP_mult_208_n1116), .S(DP_mult_208_n1117) );
  FA_X1 DP_mult_208_U765 ( .A(DP_mult_208_n1130), .B(DP_mult_208_n1121), .CI(
        DP_mult_208_n1128), .CO(DP_mult_208_n1114), .S(DP_mult_208_n1115) );
  FA_X1 DP_mult_208_U764 ( .A(DP_mult_208_n1119), .B(DP_mult_208_n1117), .CI(
        DP_mult_208_n1126), .CO(DP_mult_208_n1112), .S(DP_mult_208_n1113) );
  FA_X1 DP_mult_208_U763 ( .A(DP_mult_208_n1124), .B(DP_mult_208_n1115), .CI(
        DP_mult_208_n1113), .CO(DP_mult_208_n1110), .S(DP_mult_208_n1111) );
  FA_X1 DP_mult_208_U762 ( .A(DP_mult_208_n1335), .B(DP_mult_208_n1468), .CI(
        DP_mult_208_n1357), .CO(DP_mult_208_n1108), .S(DP_mult_208_n1109) );
  FA_X1 DP_mult_208_U761 ( .A(DP_mult_208_n1379), .B(DP_mult_208_n1445), .CI(
        DP_mult_208_n1401), .CO(DP_mult_208_n1106), .S(DP_mult_208_n1107) );
  FA_X1 DP_mult_208_U760 ( .A(DP_mult_208_n1120), .B(DP_mult_208_n1423), .CI(
        DP_mult_208_n1118), .CO(DP_mult_208_n1104), .S(DP_mult_208_n1105) );
  FA_X1 DP_mult_208_U759 ( .A(DP_mult_208_n1313), .B(DP_mult_208_n1116), .CI(
        DP_mult_208_n1107), .CO(DP_mult_208_n1102), .S(DP_mult_208_n1103) );
  FA_X1 DP_mult_208_U758 ( .A(DP_mult_208_n1114), .B(DP_mult_208_n1109), .CI(
        DP_mult_208_n1105), .CO(DP_mult_208_n1100), .S(DP_mult_208_n1101) );
  FA_X1 DP_mult_208_U757 ( .A(DP_mult_208_n1103), .B(DP_mult_208_n1112), .CI(
        DP_mult_208_n1101), .CO(DP_mult_208_n1098), .S(DP_mult_208_n1099) );
  HA_X1 DP_mult_208_U756 ( .A(DP_mult_208_n1312), .B(DP_mult_208_n1334), .CO(
        DP_mult_208_n1096), .S(DP_mult_208_n1097) );
  FA_X1 DP_mult_208_U755 ( .A(DP_mult_208_n1467), .B(DP_mult_208_n1186), .CI(
        DP_mult_208_n1400), .CO(DP_mult_208_n1094), .S(DP_mult_208_n1095) );
  FA_X1 DP_mult_208_U754 ( .A(DP_mult_208_n1356), .B(DP_mult_208_n1444), .CI(
        DP_mult_208_n1378), .CO(DP_mult_208_n1092), .S(DP_mult_208_n1093) );
  FA_X1 DP_mult_208_U753 ( .A(DP_mult_208_n1097), .B(DP_mult_208_n1422), .CI(
        DP_mult_208_n1108), .CO(DP_mult_208_n1090), .S(DP_mult_208_n1091) );
  FA_X1 DP_mult_208_U752 ( .A(DP_mult_208_n1093), .B(DP_mult_208_n1106), .CI(
        DP_mult_208_n1095), .CO(DP_mult_208_n1088), .S(DP_mult_208_n1089) );
  FA_X1 DP_mult_208_U751 ( .A(DP_mult_208_n1102), .B(DP_mult_208_n1104), .CI(
        DP_mult_208_n1091), .CO(DP_mult_208_n1086), .S(DP_mult_208_n1087) );
  FA_X1 DP_mult_208_U750 ( .A(DP_mult_208_n1100), .B(DP_mult_208_n1089), .CI(
        DP_mult_208_n1087), .CO(DP_mult_208_n1084), .S(DP_mult_208_n1085) );
  FA_X1 DP_mult_208_U749 ( .A(DP_mult_208_n1311), .B(DP_mult_208_n1333), .CI(
        DP_mult_208_n1466), .CO(DP_mult_208_n1082), .S(DP_mult_208_n1083) );
  FA_X1 DP_mult_208_U748 ( .A(DP_mult_208_n1355), .B(DP_mult_208_n1443), .CI(
        DP_mult_208_n1377), .CO(DP_mult_208_n1080), .S(DP_mult_208_n1081) );
  FA_X1 DP_mult_208_U747 ( .A(DP_mult_208_n1399), .B(DP_mult_208_n1421), .CI(
        DP_mult_208_n1096), .CO(DP_mult_208_n1078), .S(DP_mult_208_n1079) );
  FA_X1 DP_mult_208_U746 ( .A(DP_mult_208_n1092), .B(DP_mult_208_n1094), .CI(
        DP_mult_208_n1289), .CO(DP_mult_208_n1076), .S(DP_mult_208_n1077) );
  FA_X1 DP_mult_208_U745 ( .A(DP_mult_208_n1083), .B(DP_mult_208_n1081), .CI(
        DP_mult_208_n1079), .CO(DP_mult_208_n1074), .S(DP_mult_208_n1075) );
  FA_X1 DP_mult_208_U744 ( .A(DP_mult_208_n1088), .B(DP_mult_208_n1090), .CI(
        DP_mult_208_n1077), .CO(DP_mult_208_n1072), .S(DP_mult_208_n1073) );
  FA_X1 DP_mult_208_U743 ( .A(DP_mult_208_n1086), .B(DP_mult_208_n1075), .CI(
        DP_mult_208_n1073), .CO(DP_mult_208_n1070), .S(DP_mult_208_n1071) );
  HA_X1 DP_mult_208_U742 ( .A(DP_mult_208_n1288), .B(DP_mult_208_n1310), .CO(
        DP_mult_208_n1068), .S(DP_mult_208_n1069) );
  FA_X1 DP_mult_208_U741 ( .A(DP_mult_208_n1465), .B(DP_mult_208_n1376), .CI(
        DP_mult_208_n1185), .CO(DP_mult_208_n1066), .S(DP_mult_208_n1067) );
  FA_X1 DP_mult_208_U740 ( .A(DP_mult_208_n1442), .B(DP_mult_208_n1354), .CI(
        DP_mult_208_n1332), .CO(DP_mult_208_n1064), .S(DP_mult_208_n1065) );
  FA_X1 DP_mult_208_U739 ( .A(DP_mult_208_n1398), .B(DP_mult_208_n1420), .CI(
        DP_mult_208_n1069), .CO(DP_mult_208_n1062), .S(DP_mult_208_n1063) );
  FA_X1 DP_mult_208_U738 ( .A(DP_mult_208_n1080), .B(DP_mult_208_n1082), .CI(
        DP_mult_208_n1078), .CO(DP_mult_208_n1060), .S(DP_mult_208_n1061) );
  FA_X1 DP_mult_208_U737 ( .A(DP_mult_208_n1067), .B(DP_mult_208_n1065), .CI(
        DP_mult_208_n1076), .CO(DP_mult_208_n1058), .S(DP_mult_208_n1059) );
  FA_X1 DP_mult_208_U736 ( .A(DP_mult_208_n1061), .B(DP_mult_208_n1063), .CI(
        DP_mult_208_n1074), .CO(DP_mult_208_n1056), .S(DP_mult_208_n1057) );
  FA_X1 DP_mult_208_U735 ( .A(DP_mult_208_n1072), .B(DP_mult_208_n1059), .CI(
        DP_mult_208_n1057), .CO(DP_mult_208_n1054), .S(DP_mult_208_n1055) );
  FA_X1 DP_mult_208_U734 ( .A(DP_mult_208_n1309), .B(DP_mult_208_n1464), .CI(
        DP_mult_208_n1287), .CO(DP_mult_208_n1052), .S(DP_mult_208_n1053) );
  FA_X1 DP_mult_208_U733 ( .A(DP_mult_208_n1331), .B(DP_mult_208_n1353), .CI(
        DP_mult_208_n1375), .CO(DP_mult_208_n1050), .S(DP_mult_208_n1051) );
  FA_X1 DP_mult_208_U732 ( .A(DP_mult_208_n1397), .B(DP_mult_208_n1441), .CI(
        DP_mult_208_n1419), .CO(DP_mult_208_n1048), .S(DP_mult_208_n1049) );
  FA_X1 DP_mult_208_U731 ( .A(DP_mult_208_n1064), .B(DP_mult_208_n1068), .CI(
        DP_mult_208_n1066), .CO(DP_mult_208_n1046), .S(DP_mult_208_n1047) );
  FA_X1 DP_mult_208_U730 ( .A(DP_mult_208_n1049), .B(DP_mult_208_n1265), .CI(
        DP_mult_208_n1051), .CO(DP_mult_208_n1044), .S(DP_mult_208_n1045) );
  FA_X1 DP_mult_208_U729 ( .A(DP_mult_208_n1062), .B(DP_mult_208_n1053), .CI(
        DP_mult_208_n1060), .CO(DP_mult_208_n1042), .S(DP_mult_208_n1043) );
  FA_X1 DP_mult_208_U728 ( .A(DP_mult_208_n1058), .B(DP_mult_208_n1047), .CI(
        DP_mult_208_n1045), .CO(DP_mult_208_n1040), .S(DP_mult_208_n1041) );
  HA_X1 DP_mult_208_U726 ( .A(DP_mult_208_n1264), .B(DP_mult_208_n1286), .CO(
        DP_mult_208_n1036), .S(DP_mult_208_n1037) );
  FA_X1 DP_mult_208_U725 ( .A(DP_mult_208_n1308), .B(DP_mult_208_n1374), .CI(
        DP_mult_208_n1184), .CO(DP_mult_208_n1034), .S(DP_mult_208_n1035) );
  FA_X1 DP_mult_208_U723 ( .A(DP_mult_208_n1352), .B(DP_mult_208_n1440), .CI(
        DP_mult_208_n1418), .CO(DP_mult_208_n1030), .S(DP_mult_208_n1031) );
  FA_X1 DP_mult_208_U722 ( .A(DP_mult_208_n1052), .B(DP_mult_208_n1037), .CI(
        DP_mult_208_n1050), .CO(DP_mult_208_n1028), .S(DP_mult_208_n1029) );
  FA_X1 DP_mult_208_U721 ( .A(DP_mult_208_n1031), .B(DP_mult_208_n1048), .CI(
        DP_mult_208_n1033), .CO(DP_mult_208_n1026), .S(DP_mult_208_n1027) );
  FA_X1 DP_mult_208_U720 ( .A(DP_mult_208_n1046), .B(DP_mult_208_n1035), .CI(
        DP_mult_208_n1029), .CO(DP_mult_208_n1024), .S(DP_mult_208_n1025) );
  FA_X1 DP_mult_208_U719 ( .A(DP_mult_208_n1027), .B(DP_mult_208_n1044), .CI(
        DP_mult_208_n1042), .CO(DP_mult_208_n1022), .S(DP_mult_208_n1023) );
  FA_X1 DP_mult_208_U718 ( .A(DP_mult_208_n1040), .B(DP_mult_208_n1025), .CI(
        DP_mult_208_n1023), .CO(DP_mult_208_n1020), .S(DP_mult_208_n1021) );
  FA_X1 DP_mult_208_U717 ( .A(DP_mult_208_n1263), .B(DP_mult_208_n1351), .CI(
        DP_mult_208_n1285), .CO(DP_mult_208_n1018), .S(DP_mult_208_n1019) );
  FA_X1 DP_mult_208_U716 ( .A(DP_mult_208_n1307), .B(DP_mult_208_n1373), .CI(
        DP_mult_208_n1329), .CO(DP_mult_208_n1016), .S(DP_mult_208_n1017) );
  FA_X1 DP_mult_208_U715 ( .A(DP_mult_208_n1395), .B(DP_mult_208_n1462), .CI(
        DP_mult_208_n1417), .CO(DP_mult_208_n1014), .S(DP_mult_208_n1015) );
  FA_X1 DP_mult_208_U714 ( .A(DP_mult_208_n1036), .B(DP_mult_208_n1439), .CI(
        DP_mult_208_n1032), .CO(DP_mult_208_n1012), .S(DP_mult_208_n1013) );
  FA_X1 DP_mult_208_U713 ( .A(DP_mult_208_n1030), .B(DP_mult_208_n1034), .CI(
        DP_mult_208_n1241), .CO(DP_mult_208_n1010), .S(DP_mult_208_n1011) );
  FA_X1 DP_mult_208_U712 ( .A(DP_mult_208_n1019), .B(DP_mult_208_n1015), .CI(
        DP_mult_208_n1017), .CO(DP_mult_208_n1008), .S(DP_mult_208_n1009) );
  FA_X1 DP_mult_208_U711 ( .A(DP_mult_208_n1013), .B(DP_mult_208_n1028), .CI(
        DP_mult_208_n1026), .CO(DP_mult_208_n1006), .S(DP_mult_208_n1007) );
  FA_X1 DP_mult_208_U710 ( .A(DP_mult_208_n1009), .B(DP_mult_208_n1011), .CI(
        DP_mult_208_n1024), .CO(DP_mult_208_n1004), .S(DP_mult_208_n1005) );
  FA_X1 DP_mult_208_U709 ( .A(DP_mult_208_n1022), .B(DP_mult_208_n1007), .CI(
        DP_mult_208_n1005), .CO(DP_mult_208_n1002), .S(DP_mult_208_n1003) );
  FA_X1 DP_mult_208_U707 ( .A(DP_mult_208_n1461), .B(DP_mult_208_n1350), .CI(
        DP_mult_208_n1183), .CO(DP_mult_208_n998), .S(DP_mult_208_n999) );
  FA_X1 DP_mult_208_U704 ( .A(DP_mult_208_n1018), .B(DP_mult_208_n1394), .CI(
        DP_mult_208_n1001), .CO(DP_mult_208_n992), .S(DP_mult_208_n993) );
  FA_X1 DP_mult_208_U703 ( .A(DP_mult_208_n1014), .B(DP_mult_208_n1016), .CI(
        DP_mult_208_n995), .CO(DP_mult_208_n990), .S(DP_mult_208_n991) );
  FA_X1 DP_mult_208_U702 ( .A(DP_mult_208_n999), .B(DP_mult_208_n997), .CI(
        DP_mult_208_n1012), .CO(DP_mult_208_n988), .S(DP_mult_208_n989) );
  FA_X1 DP_mult_208_U701 ( .A(DP_mult_208_n993), .B(DP_mult_208_n1010), .CI(
        DP_mult_208_n1008), .CO(DP_mult_208_n986), .S(DP_mult_208_n987) );
  FA_X1 DP_mult_208_U700 ( .A(DP_mult_208_n989), .B(DP_mult_208_n991), .CI(
        DP_mult_208_n1006), .CO(DP_mult_208_n984), .S(DP_mult_208_n985) );
  FA_X1 DP_mult_208_U699 ( .A(DP_mult_208_n1004), .B(DP_mult_208_n987), .CI(
        DP_mult_208_n985), .CO(DP_mult_208_n982), .S(DP_mult_208_n983) );
  FA_X1 DP_mult_208_U698 ( .A(DP_mult_208_n1239), .B(DP_mult_208_n1349), .CI(
        DP_mult_208_n1261), .CO(DP_mult_208_n980), .S(DP_mult_208_n981) );
  FA_X1 DP_mult_208_U697 ( .A(DP_mult_208_n1460), .B(DP_mult_208_n1283), .CI(
        DP_mult_208_n1371), .CO(DP_mult_208_n978), .S(DP_mult_208_n979) );
  FA_X1 DP_mult_208_U696 ( .A(DP_mult_208_n1327), .B(DP_mult_208_n1437), .CI(
        DP_mult_208_n1305), .CO(DP_mult_208_n976), .S(DP_mult_208_n977) );
  FA_X1 DP_mult_208_U693 ( .A(DP_mult_208_n977), .B(DP_mult_208_n998), .CI(
        DP_mult_208_n979), .CO(DP_mult_208_n970), .S(DP_mult_208_n971) );
  FA_X1 DP_mult_208_U692 ( .A(DP_mult_208_n975), .B(DP_mult_208_n981), .CI(
        DP_mult_208_n992), .CO(DP_mult_208_n968), .S(DP_mult_208_n969) );
  FA_X1 DP_mult_208_U691 ( .A(DP_mult_208_n973), .B(DP_mult_208_n990), .CI(
        DP_mult_208_n988), .CO(DP_mult_208_n966), .S(DP_mult_208_n967) );
  FA_X1 DP_mult_208_U690 ( .A(DP_mult_208_n969), .B(DP_mult_208_n971), .CI(
        DP_mult_208_n986), .CO(DP_mult_208_n964), .S(DP_mult_208_n965) );
  FA_X1 DP_mult_208_U689 ( .A(DP_mult_208_n984), .B(DP_mult_208_n967), .CI(
        DP_mult_208_n965), .CO(DP_mult_208_n962), .S(DP_mult_208_n963) );
  FA_X1 DP_mult_208_U683 ( .A(DP_mult_208_n976), .B(DP_mult_208_n980), .CI(
        DP_mult_208_n978), .CO(DP_mult_208_n950), .S(DP_mult_208_n951) );
  FA_X1 DP_mult_208_U682 ( .A(DP_mult_208_n955), .B(DP_mult_208_n974), .CI(
        DP_mult_208_n957), .CO(DP_mult_208_n948), .S(DP_mult_208_n949) );
  FA_X1 DP_mult_208_U681 ( .A(DP_mult_208_n972), .B(DP_mult_208_n959), .CI(
        DP_mult_208_n953), .CO(DP_mult_208_n946), .S(DP_mult_208_n947) );
  FA_X1 DP_mult_208_U680 ( .A(DP_mult_208_n970), .B(DP_mult_208_n951), .CI(
        DP_mult_208_n968), .CO(DP_mult_208_n944), .S(DP_mult_208_n945) );
  FA_X1 DP_mult_208_U679 ( .A(DP_mult_208_n947), .B(DP_mult_208_n949), .CI(
        DP_mult_208_n966), .CO(DP_mult_208_n942), .S(DP_mult_208_n943) );
  FA_X1 DP_mult_208_U678 ( .A(DP_mult_208_n964), .B(DP_mult_208_n945), .CI(
        DP_mult_208_n943), .CO(DP_mult_208_n940), .S(DP_mult_208_n941) );
  FA_X1 DP_mult_208_U675 ( .A(DP_mult_208_n1259), .B(DP_mult_208_n1347), .CI(
        DP_mult_208_n1303), .CO(DP_mult_208_n936), .S(DP_mult_208_n937) );
  FA_X1 DP_mult_208_U674 ( .A(DP_mult_208_n1281), .B(DP_mult_208_n1369), .CI(
        DP_mult_208_n1391), .CO(DP_mult_208_n934), .S(DP_mult_208_n935) );
  FA_X1 DP_mult_208_U673 ( .A(DP_mult_208_n1325), .B(DP_mult_208_n1413), .CI(
        DP_mult_208_n1435), .CO(DP_mult_208_n932), .S(DP_mult_208_n933) );
  FA_X1 DP_mult_208_U672 ( .A(DP_mult_208_n1458), .B(DP_mult_208_n1980), .CI(
        DP_mult_208_n939), .CO(DP_mult_208_n930), .S(DP_mult_208_n931) );
  FA_X1 DP_mult_208_U670 ( .A(DP_mult_208_n933), .B(DP_mult_208_n937), .CI(
        DP_mult_208_n952), .CO(DP_mult_208_n926), .S(DP_mult_208_n927) );
  FA_X1 DP_mult_208_U669 ( .A(DP_mult_208_n950), .B(DP_mult_208_n935), .CI(
        DP_mult_208_n931), .CO(DP_mult_208_n924), .S(DP_mult_208_n925) );
  FA_X1 DP_mult_208_U668 ( .A(DP_mult_208_n929), .B(DP_mult_208_n948), .CI(
        DP_mult_208_n946), .CO(DP_mult_208_n922), .S(DP_mult_208_n923) );
  FA_X1 DP_mult_208_U664 ( .A(DP_mult_208_n1214), .B(DP_mult_208_n1302), .CI(
        DP_mult_208_n917), .CO(DP_mult_208_n914), .S(DP_mult_208_n915) );
  FA_X1 DP_mult_208_U663 ( .A(DP_mult_208_n1236), .B(DP_mult_208_n1412), .CI(
        DP_mult_208_n1258), .CO(DP_mult_208_n912), .S(DP_mult_208_n913) );
  FA_X1 DP_mult_208_U662 ( .A(DP_mult_208_n1280), .B(DP_mult_208_n1346), .CI(
        DP_mult_208_n1324), .CO(DP_mult_208_n910), .S(DP_mult_208_n911) );
  FA_X1 DP_mult_208_U661 ( .A(DP_mult_208_n1368), .B(DP_mult_208_n1390), .CI(
        DP_mult_208_n938), .CO(DP_mult_208_n908), .S(DP_mult_208_n909) );
  FA_X1 DP_mult_208_U660 ( .A(DP_mult_208_n932), .B(DP_mult_208_n936), .CI(
        DP_mult_208_n934), .CO(DP_mult_208_n906), .S(DP_mult_208_n907) );
  FA_X1 DP_mult_208_U659 ( .A(DP_mult_208_n913), .B(DP_mult_208_n911), .CI(
        DP_mult_208_n915), .CO(DP_mult_208_n904), .S(DP_mult_208_n905) );
  FA_X1 DP_mult_208_U658 ( .A(DP_mult_208_n909), .B(DP_mult_208_n930), .CI(
        DP_mult_208_n928), .CO(DP_mult_208_n902), .S(DP_mult_208_n903) );
  FA_X1 DP_mult_208_U657 ( .A(DP_mult_208_n926), .B(DP_mult_208_n907), .CI(
        DP_mult_208_n905), .CO(DP_mult_208_n900), .S(DP_mult_208_n901) );
  FA_X1 DP_mult_208_U656 ( .A(DP_mult_208_n903), .B(DP_mult_208_n924), .CI(
        DP_mult_208_n922), .CO(DP_mult_208_n898), .S(DP_mult_208_n899) );
  FA_X1 DP_mult_208_U655 ( .A(DP_mult_208_n920), .B(DP_mult_208_n901), .CI(
        DP_mult_208_n899), .CO(DP_mult_208_n896), .S(DP_mult_208_n897) );
  FA_X1 DP_mult_208_U654 ( .A(DP_mult_208_n1411), .B(DP_mult_208_n1213), .CI(
        DP_mult_208_n1235), .CO(DP_mult_208_n894), .S(DP_mult_208_n895) );
  FA_X1 DP_mult_208_U653 ( .A(DP_mult_208_n1323), .B(DP_mult_208_n1279), .CI(
        DP_mult_208_n916), .CO(DP_mult_208_n892), .S(DP_mult_208_n893) );
  FA_X1 DP_mult_208_U652 ( .A(DP_mult_208_n1257), .B(DP_mult_208_n1345), .CI(
        DP_mult_208_n1301), .CO(DP_mult_208_n890), .S(DP_mult_208_n891) );
  FA_X1 DP_mult_208_U651 ( .A(DP_mult_208_n1367), .B(DP_mult_208_n1389), .CI(
        DP_mult_208_n1434), .CO(DP_mult_208_n888), .S(DP_mult_208_n889) );
  FA_X1 DP_mult_208_U650 ( .A(DP_mult_208_n910), .B(DP_mult_208_n914), .CI(
        DP_mult_208_n912), .CO(DP_mult_208_n886), .S(DP_mult_208_n887) );
  FA_X1 DP_mult_208_U648 ( .A(DP_mult_208_n906), .B(DP_mult_208_n893), .CI(
        DP_mult_208_n889), .CO(DP_mult_208_n882), .S(DP_mult_208_n883) );
  FA_X1 DP_mult_208_U647 ( .A(DP_mult_208_n887), .B(DP_mult_208_n904), .CI(
        DP_mult_208_n902), .CO(DP_mult_208_n880), .S(DP_mult_208_n881) );
  FA_X1 DP_mult_208_U646 ( .A(DP_mult_208_n883), .B(DP_mult_208_n885), .CI(
        DP_mult_208_n900), .CO(DP_mult_208_n878), .S(DP_mult_208_n879) );
  FA_X1 DP_mult_208_U645 ( .A(DP_mult_208_n898), .B(DP_mult_208_n881), .CI(
        DP_mult_208_n879), .CO(DP_mult_208_n876), .S(DP_mult_208_n877) );
  FA_X1 DP_mult_208_U643 ( .A(DP_mult_208_n1388), .B(DP_mult_208_n1278), .CI(
        DP_mult_208_n875), .CO(DP_mult_208_n872), .S(DP_mult_208_n873) );
  FA_X1 DP_mult_208_U642 ( .A(DP_mult_208_n1212), .B(DP_mult_208_n1366), .CI(
        DP_mult_208_n1344), .CO(DP_mult_208_n870), .S(DP_mult_208_n871) );
  FA_X1 DP_mult_208_U641 ( .A(DP_mult_208_n1234), .B(DP_mult_208_n1322), .CI(
        DP_mult_208_n1256), .CO(DP_mult_208_n868), .S(DP_mult_208_n869) );
  FA_X1 DP_mult_208_U640 ( .A(DP_mult_208_n894), .B(DP_mult_208_n1300), .CI(
        DP_mult_208_n892), .CO(DP_mult_208_n866), .S(DP_mult_208_n867) );
  FA_X1 DP_mult_208_U639 ( .A(DP_mult_208_n871), .B(DP_mult_208_n890), .CI(
        DP_mult_208_n869), .CO(DP_mult_208_n864), .S(DP_mult_208_n865) );
  FA_X1 DP_mult_208_U636 ( .A(DP_mult_208_n863), .B(DP_mult_208_n882), .CI(
        DP_mult_208_n880), .CO(DP_mult_208_n858), .S(DP_mult_208_n859) );
  FA_X1 DP_mult_208_U635 ( .A(DP_mult_208_n878), .B(DP_mult_208_n861), .CI(
        DP_mult_208_n859), .CO(DP_mult_208_n856), .S(DP_mult_208_n857) );
  FA_X1 DP_mult_208_U634 ( .A(DP_mult_208_n1387), .B(DP_mult_208_n1211), .CI(
        DP_mult_208_n1233), .CO(DP_mult_208_n854), .S(DP_mult_208_n855) );
  FA_X1 DP_mult_208_U633 ( .A(DP_mult_208_n1255), .B(DP_mult_208_n1321), .CI(
        DP_mult_208_n874), .CO(DP_mult_208_n852), .S(DP_mult_208_n853) );
  FA_X1 DP_mult_208_U632 ( .A(DP_mult_208_n1343), .B(DP_mult_208_n1277), .CI(
        DP_mult_208_n1299), .CO(DP_mult_208_n850), .S(DP_mult_208_n851) );
  FA_X1 DP_mult_208_U631 ( .A(DP_mult_208_n1410), .B(DP_mult_208_n1365), .CI(
        DP_mult_208_n872), .CO(DP_mult_208_n848), .S(DP_mult_208_n849) );
  FA_X1 DP_mult_208_U630 ( .A(DP_mult_208_n868), .B(DP_mult_208_n870), .CI(
        DP_mult_208_n851), .CO(DP_mult_208_n846), .S(DP_mult_208_n847) );
  FA_X1 DP_mult_208_U629 ( .A(DP_mult_208_n855), .B(DP_mult_208_n853), .CI(
        DP_mult_208_n866), .CO(DP_mult_208_n844), .S(DP_mult_208_n845) );
  FA_X1 DP_mult_208_U627 ( .A(DP_mult_208_n845), .B(DP_mult_208_n847), .CI(
        DP_mult_208_n860), .CO(DP_mult_208_n840), .S(DP_mult_208_n841) );
  FA_X1 DP_mult_208_U626 ( .A(DP_mult_208_n858), .B(DP_mult_208_n843), .CI(
        DP_mult_208_n841), .CO(DP_mult_208_n838), .S(DP_mult_208_n839) );
  FA_X1 DP_mult_208_U624 ( .A(DP_mult_208_n1210), .B(DP_mult_208_n837), .CI(
        DP_mult_208_n1276), .CO(DP_mult_208_n834), .S(DP_mult_208_n835) );
  FA_X1 DP_mult_208_U623 ( .A(DP_mult_208_n1232), .B(DP_mult_208_n1364), .CI(
        DP_mult_208_n1342), .CO(DP_mult_208_n832), .S(DP_mult_208_n833) );
  FA_X1 DP_mult_208_U622 ( .A(DP_mult_208_n1254), .B(DP_mult_208_n1298), .CI(
        DP_mult_208_n1320), .CO(DP_mult_208_n830), .S(DP_mult_208_n831) );
  FA_X1 DP_mult_208_U621 ( .A(DP_mult_208_n850), .B(DP_mult_208_n854), .CI(
        DP_mult_208_n852), .CO(DP_mult_208_n828), .S(DP_mult_208_n829) );
  FA_X1 DP_mult_208_U620 ( .A(DP_mult_208_n835), .B(DP_mult_208_n831), .CI(
        DP_mult_208_n833), .CO(DP_mult_208_n826), .S(DP_mult_208_n827) );
  FA_X1 DP_mult_208_U619 ( .A(DP_mult_208_n846), .B(DP_mult_208_n848), .CI(
        DP_mult_208_n829), .CO(DP_mult_208_n824), .S(DP_mult_208_n825) );
  FA_X1 DP_mult_208_U616 ( .A(DP_mult_208_n1363), .B(DP_mult_208_n1209), .CI(
        DP_mult_208_n2069), .CO(DP_mult_208_n818), .S(DP_mult_208_n819) );
  FA_X1 DP_mult_208_U615 ( .A(DP_mult_208_n1231), .B(DP_mult_208_n1297), .CI(
        DP_mult_208_n1275), .CO(DP_mult_208_n816), .S(DP_mult_208_n817) );
  FA_X1 DP_mult_208_U614 ( .A(DP_mult_208_n1319), .B(DP_mult_208_n1253), .CI(
        DP_mult_208_n1341), .CO(DP_mult_208_n814), .S(DP_mult_208_n815) );
  FA_X1 DP_mult_208_U613 ( .A(DP_mult_208_n1386), .B(DP_mult_208_n830), .CI(
        DP_mult_208_n834), .CO(DP_mult_208_n812), .S(DP_mult_208_n813) );
  FA_X1 DP_mult_208_U612 ( .A(DP_mult_208_n815), .B(DP_mult_208_n832), .CI(
        DP_mult_208_n817), .CO(DP_mult_208_n810), .S(DP_mult_208_n811) );
  FA_X1 DP_mult_208_U611 ( .A(DP_mult_208_n828), .B(DP_mult_208_n819), .CI(
        DP_mult_208_n813), .CO(DP_mult_208_n808), .S(DP_mult_208_n809) );
  FA_X1 DP_mult_208_U610 ( .A(DP_mult_208_n811), .B(DP_mult_208_n826), .CI(
        DP_mult_208_n824), .CO(DP_mult_208_n806), .S(DP_mult_208_n807) );
  FA_X1 DP_mult_208_U609 ( .A(DP_mult_208_n822), .B(DP_mult_208_n809), .CI(
        DP_mult_208_n807), .CO(DP_mult_208_n804), .S(DP_mult_208_n805) );
  FA_X1 DP_mult_208_U607 ( .A(DP_mult_208_n1340), .B(DP_mult_208_n1252), .CI(
        DP_mult_208_n803), .CO(DP_mult_208_n800), .S(DP_mult_208_n801) );
  FA_X1 DP_mult_208_U606 ( .A(DP_mult_208_n1208), .B(DP_mult_208_n1318), .CI(
        DP_mult_208_n1230), .CO(DP_mult_208_n798), .S(DP_mult_208_n799) );
  FA_X1 DP_mult_208_U604 ( .A(DP_mult_208_n814), .B(DP_mult_208_n816), .CI(
        DP_mult_208_n799), .CO(DP_mult_208_n794), .S(DP_mult_208_n795) );
  FA_X1 DP_mult_208_U603 ( .A(DP_mult_208_n797), .B(DP_mult_208_n801), .CI(
        DP_mult_208_n812), .CO(DP_mult_208_n792), .S(DP_mult_208_n793) );
  FA_X1 DP_mult_208_U602 ( .A(DP_mult_208_n795), .B(DP_mult_208_n810), .CI(
        DP_mult_208_n808), .CO(DP_mult_208_n790), .S(DP_mult_208_n791) );
  FA_X1 DP_mult_208_U601 ( .A(DP_mult_208_n806), .B(DP_mult_208_n793), .CI(
        DP_mult_208_n791), .CO(DP_mult_208_n788), .S(DP_mult_208_n789) );
  FA_X1 DP_mult_208_U600 ( .A(DP_mult_208_n1251), .B(DP_mult_208_n1207), .CI(
        DP_mult_208_n802), .CO(DP_mult_208_n786), .S(DP_mult_208_n787) );
  FA_X1 DP_mult_208_U599 ( .A(DP_mult_208_n1273), .B(DP_mult_208_n1317), .CI(
        DP_mult_208_n1295), .CO(DP_mult_208_n784), .S(DP_mult_208_n785) );
  FA_X1 DP_mult_208_U598 ( .A(DP_mult_208_n1339), .B(DP_mult_208_n1229), .CI(
        DP_mult_208_n1362), .CO(DP_mult_208_n782), .S(DP_mult_208_n783) );
  FA_X1 DP_mult_208_U597 ( .A(DP_mult_208_n798), .B(DP_mult_208_n800), .CI(
        DP_mult_208_n785), .CO(DP_mult_208_n780), .S(DP_mult_208_n781) );
  FA_X1 DP_mult_208_U596 ( .A(DP_mult_208_n796), .B(DP_mult_208_n787), .CI(
        DP_mult_208_n783), .CO(DP_mult_208_n778), .S(DP_mult_208_n779) );
  FA_X1 DP_mult_208_U595 ( .A(DP_mult_208_n781), .B(DP_mult_208_n794), .CI(
        DP_mult_208_n792), .CO(DP_mult_208_n776), .S(DP_mult_208_n777) );
  FA_X1 DP_mult_208_U594 ( .A(DP_mult_208_n790), .B(DP_mult_208_n779), .CI(
        DP_mult_208_n777), .CO(DP_mult_208_n774), .S(DP_mult_208_n775) );
  FA_X1 DP_mult_208_U592 ( .A(DP_mult_208_n1316), .B(DP_mult_208_n1250), .CI(
        DP_mult_208_n773), .CO(DP_mult_208_n770), .S(DP_mult_208_n771) );
  FA_X1 DP_mult_208_U591 ( .A(DP_mult_208_n1294), .B(DP_mult_208_n1206), .CI(
        DP_mult_208_n1272), .CO(DP_mult_208_n768), .S(DP_mult_208_n769) );
  FA_X1 DP_mult_208_U590 ( .A(DP_mult_208_n786), .B(DP_mult_208_n1228), .CI(
        DP_mult_208_n784), .CO(DP_mult_208_n766), .S(DP_mult_208_n767) );
  FA_X1 DP_mult_208_U589 ( .A(DP_mult_208_n771), .B(DP_mult_208_n769), .CI(
        DP_mult_208_n782), .CO(DP_mult_208_n764), .S(DP_mult_208_n765) );
  FA_X1 DP_mult_208_U588 ( .A(DP_mult_208_n767), .B(DP_mult_208_n780), .CI(
        DP_mult_208_n778), .CO(DP_mult_208_n762), .S(DP_mult_208_n763) );
  FA_X1 DP_mult_208_U587 ( .A(DP_mult_208_n776), .B(DP_mult_208_n765), .CI(
        DP_mult_208_n763), .CO(DP_mult_208_n760), .S(DP_mult_208_n761) );
  FA_X1 DP_mult_208_U586 ( .A(DP_mult_208_n772), .B(DP_mult_208_n1205), .CI(
        DP_mult_208_n1227), .CO(DP_mult_208_n758), .S(DP_mult_208_n759) );
  FA_X1 DP_mult_208_U585 ( .A(DP_mult_208_n1249), .B(DP_mult_208_n1293), .CI(
        DP_mult_208_n1315), .CO(DP_mult_208_n756), .S(DP_mult_208_n757) );
  FA_X1 DP_mult_208_U584 ( .A(DP_mult_208_n1338), .B(DP_mult_208_n1271), .CI(
        DP_mult_208_n770), .CO(DP_mult_208_n754), .S(DP_mult_208_n755) );
  FA_X1 DP_mult_208_U583 ( .A(DP_mult_208_n757), .B(DP_mult_208_n768), .CI(
        DP_mult_208_n759), .CO(DP_mult_208_n752), .S(DP_mult_208_n753) );
  FA_X1 DP_mult_208_U582 ( .A(DP_mult_208_n755), .B(DP_mult_208_n766), .CI(
        DP_mult_208_n764), .CO(DP_mult_208_n750), .S(DP_mult_208_n751) );
  FA_X1 DP_mult_208_U581 ( .A(DP_mult_208_n762), .B(DP_mult_208_n753), .CI(
        DP_mult_208_n751), .CO(DP_mult_208_n748), .S(DP_mult_208_n749) );
  FA_X1 DP_mult_208_U579 ( .A(DP_mult_208_n1292), .B(DP_mult_208_n1248), .CI(
        DP_mult_208_n747), .CO(DP_mult_208_n744), .S(DP_mult_208_n745) );
  FA_X1 DP_mult_208_U578 ( .A(DP_mult_208_n1226), .B(DP_mult_208_n1204), .CI(
        DP_mult_208_n1270), .CO(DP_mult_208_n742), .S(DP_mult_208_n743) );
  FA_X1 DP_mult_208_U577 ( .A(DP_mult_208_n756), .B(DP_mult_208_n758), .CI(
        DP_mult_208_n743), .CO(DP_mult_208_n740), .S(DP_mult_208_n741) );
  FA_X1 DP_mult_208_U576 ( .A(DP_mult_208_n754), .B(DP_mult_208_n745), .CI(
        DP_mult_208_n752), .CO(DP_mult_208_n738), .S(DP_mult_208_n739) );
  FA_X1 DP_mult_208_U575 ( .A(DP_mult_208_n750), .B(DP_mult_208_n741), .CI(
        DP_mult_208_n739), .CO(DP_mult_208_n736), .S(DP_mult_208_n737) );
  FA_X1 DP_mult_208_U574 ( .A(DP_mult_208_n746), .B(DP_mult_208_n1203), .CI(
        DP_mult_208_n1247), .CO(DP_mult_208_n734), .S(DP_mult_208_n735) );
  FA_X1 DP_mult_208_U573 ( .A(DP_mult_208_n1225), .B(DP_mult_208_n1291), .CI(
        DP_mult_208_n1269), .CO(DP_mult_208_n732), .S(DP_mult_208_n733) );
  FA_X1 DP_mult_208_U572 ( .A(DP_mult_208_n744), .B(DP_mult_208_n1314), .CI(
        DP_mult_208_n742), .CO(DP_mult_208_n730), .S(DP_mult_208_n731) );
  FA_X1 DP_mult_208_U571 ( .A(DP_mult_208_n735), .B(DP_mult_208_n733), .CI(
        DP_mult_208_n740), .CO(DP_mult_208_n728), .S(DP_mult_208_n729) );
  FA_X1 DP_mult_208_U570 ( .A(DP_mult_208_n738), .B(DP_mult_208_n731), .CI(
        DP_mult_208_n729), .CO(DP_mult_208_n726), .S(DP_mult_208_n727) );
  FA_X1 DP_mult_208_U568 ( .A(DP_mult_208_n1268), .B(DP_mult_208_n1224), .CI(
        DP_mult_208_n725), .CO(DP_mult_208_n722), .S(DP_mult_208_n723) );
  FA_X1 DP_mult_208_U567 ( .A(DP_mult_208_n1202), .B(DP_mult_208_n1246), .CI(
        DP_mult_208_n734), .CO(DP_mult_208_n720), .S(DP_mult_208_n721) );
  FA_X1 DP_mult_208_U566 ( .A(DP_mult_208_n723), .B(DP_mult_208_n732), .CI(
        DP_mult_208_n730), .CO(DP_mult_208_n718), .S(DP_mult_208_n719) );
  FA_X1 DP_mult_208_U565 ( .A(DP_mult_208_n728), .B(DP_mult_208_n721), .CI(
        DP_mult_208_n719), .CO(DP_mult_208_n716), .S(DP_mult_208_n717) );
  FA_X1 DP_mult_208_U564 ( .A(DP_mult_208_n1267), .B(DP_mult_208_n1201), .CI(
        DP_mult_208_n724), .CO(DP_mult_208_n714), .S(DP_mult_208_n715) );
  FA_X1 DP_mult_208_U563 ( .A(DP_mult_208_n1245), .B(DP_mult_208_n1223), .CI(
        DP_mult_208_n1290), .CO(DP_mult_208_n712), .S(DP_mult_208_n713) );
  FA_X1 DP_mult_208_U562 ( .A(DP_mult_208_n715), .B(DP_mult_208_n722), .CI(
        DP_mult_208_n720), .CO(DP_mult_208_n710), .S(DP_mult_208_n711) );
  FA_X1 DP_mult_208_U561 ( .A(DP_mult_208_n718), .B(DP_mult_208_n713), .CI(
        DP_mult_208_n711), .CO(DP_mult_208_n708), .S(DP_mult_208_n709) );
  FA_X1 DP_mult_208_U559 ( .A(DP_mult_208_n1222), .B(DP_mult_208_n1200), .CI(
        DP_mult_208_n707), .CO(DP_mult_208_n704), .S(DP_mult_208_n705) );
  FA_X1 DP_mult_208_U558 ( .A(DP_mult_208_n714), .B(DP_mult_208_n1244), .CI(
        DP_mult_208_n705), .CO(DP_mult_208_n702), .S(DP_mult_208_n703) );
  FA_X1 DP_mult_208_U557 ( .A(DP_mult_208_n710), .B(DP_mult_208_n712), .CI(
        DP_mult_208_n703), .CO(DP_mult_208_n700), .S(DP_mult_208_n701) );
  FA_X1 DP_mult_208_U556 ( .A(DP_mult_208_n1221), .B(DP_mult_208_n1199), .CI(
        DP_mult_208_n706), .CO(DP_mult_208_n698), .S(DP_mult_208_n699) );
  FA_X1 DP_mult_208_U555 ( .A(DP_mult_208_n1266), .B(DP_mult_208_n1243), .CI(
        DP_mult_208_n704), .CO(DP_mult_208_n696), .S(DP_mult_208_n697) );
  FA_X1 DP_mult_208_U554 ( .A(DP_mult_208_n702), .B(DP_mult_208_n699), .CI(
        DP_mult_208_n697), .CO(DP_mult_208_n694), .S(DP_mult_208_n695) );
  FA_X1 DP_mult_208_U552 ( .A(DP_mult_208_n1198), .B(DP_mult_208_n1220), .CI(
        DP_mult_208_n693), .CO(DP_mult_208_n690), .S(DP_mult_208_n691) );
  FA_X1 DP_mult_208_U551 ( .A(DP_mult_208_n691), .B(DP_mult_208_n698), .CI(
        DP_mult_208_n696), .CO(DP_mult_208_n688), .S(DP_mult_208_n689) );
  FA_X1 DP_mult_208_U550 ( .A(DP_mult_208_n1219), .B(DP_mult_208_n692), .CI(
        DP_mult_208_n1197), .CO(DP_mult_208_n686), .S(DP_mult_208_n687) );
  FA_X1 DP_mult_208_U549 ( .A(DP_mult_208_n690), .B(DP_mult_208_n1242), .CI(
        DP_mult_208_n687), .CO(DP_mult_208_n684), .S(DP_mult_208_n685) );
  FA_X1 DP_mult_208_U547 ( .A(DP_mult_208_n683), .B(DP_mult_208_n1196), .CI(
        DP_mult_208_n686), .CO(DP_mult_208_n680), .S(DP_mult_208_n681) );
  FA_X1 DP_mult_208_U546 ( .A(DP_mult_208_n1195), .B(DP_mult_208_n682), .CI(
        DP_mult_208_n1218), .CO(DP_mult_208_n678), .S(DP_mult_208_n679) );
  INV_X1 DP_mult_209_U2793 ( .A(DP_coeffs_ff_int[74]), .ZN(DP_mult_209_n2302)
         );
  INV_X1 DP_mult_209_U2792 ( .A(DP_coeffs_ff_int[74]), .ZN(DP_mult_209_n2301)
         );
  INV_X1 DP_mult_209_U2791 ( .A(DP_mult_209_n2302), .ZN(DP_mult_209_n2300) );
  INV_X1 DP_mult_209_U2790 ( .A(DP_coeffs_ff_int[76]), .ZN(DP_mult_209_n2297)
         );
  INV_X1 DP_mult_209_U2789 ( .A(DP_coeffs_ff_int[76]), .ZN(DP_mult_209_n2296)
         );
  INV_X1 DP_mult_209_U2788 ( .A(DP_mult_209_n2296), .ZN(DP_mult_209_n2295) );
  INV_X1 DP_mult_209_U2787 ( .A(DP_coeffs_ff_int[78]), .ZN(DP_mult_209_n2293)
         );
  INV_X1 DP_mult_209_U2786 ( .A(DP_coeffs_ff_int[78]), .ZN(DP_mult_209_n2292)
         );
  INV_X1 DP_mult_209_U2785 ( .A(DP_coeffs_ff_int[80]), .ZN(DP_mult_209_n2289)
         );
  INV_X1 DP_mult_209_U2784 ( .A(DP_coeffs_ff_int[80]), .ZN(DP_mult_209_n2288)
         );
  INV_X1 DP_mult_209_U2783 ( .A(DP_mult_209_n2289), .ZN(DP_mult_209_n2287) );
  INV_X1 DP_mult_209_U2782 ( .A(DP_coeffs_ff_int[82]), .ZN(DP_mult_209_n2283)
         );
  INV_X1 DP_mult_209_U2781 ( .A(DP_coeffs_ff_int[82]), .ZN(DP_mult_209_n2282)
         );
  INV_X1 DP_mult_209_U2780 ( .A(DP_mult_209_n2283), .ZN(DP_mult_209_n2281) );
  INV_X1 DP_mult_209_U2779 ( .A(DP_coeffs_ff_int[84]), .ZN(DP_mult_209_n2279)
         );
  INV_X1 DP_mult_209_U2778 ( .A(DP_coeffs_ff_int[84]), .ZN(DP_mult_209_n2278)
         );
  INV_X1 DP_mult_209_U2777 ( .A(DP_mult_209_n2279), .ZN(DP_mult_209_n2277) );
  INV_X1 DP_mult_209_U2776 ( .A(DP_coeffs_ff_int[86]), .ZN(DP_mult_209_n2274)
         );
  INV_X1 DP_mult_209_U2775 ( .A(DP_mult_209_n1988), .ZN(DP_mult_209_n2273) );
  INV_X1 DP_mult_209_U2774 ( .A(DP_coeffs_ff_int[88]), .ZN(DP_mult_209_n2270)
         );
  INV_X1 DP_mult_209_U2773 ( .A(DP_coeffs_ff_int[88]), .ZN(DP_mult_209_n2269)
         );
  INV_X1 DP_mult_209_U2772 ( .A(DP_coeffs_ff_int[90]), .ZN(DP_mult_209_n2265)
         );
  INV_X1 DP_mult_209_U2771 ( .A(DP_coeffs_ff_int[90]), .ZN(DP_mult_209_n2264)
         );
  INV_X1 DP_mult_209_U2770 ( .A(DP_mult_209_n2264), .ZN(DP_mult_209_n2263) );
  INV_X1 DP_mult_209_U2769 ( .A(DP_coeffs_ff_int[92]), .ZN(DP_mult_209_n2260)
         );
  INV_X1 DP_mult_209_U2768 ( .A(DP_mult_209_n2020), .ZN(DP_mult_209_n2259) );
  INV_X1 DP_mult_209_U2767 ( .A(DP_coeffs_ff_int[94]), .ZN(DP_mult_209_n2255)
         );
  INV_X1 DP_mult_209_U2766 ( .A(DP_coeffs_ff_int[94]), .ZN(DP_mult_209_n2254)
         );
  INV_X1 DP_mult_209_U2765 ( .A(DP_mult_209_n2255), .ZN(DP_mult_209_n2253) );
  INV_X1 DP_mult_209_U2764 ( .A(DP_mult_209_n2244), .ZN(DP_mult_209_n2243) );
  INV_X1 DP_mult_209_U2763 ( .A(DP_mult_209_n2186), .ZN(DP_mult_209_n2228) );
  INV_X1 DP_mult_209_U2762 ( .A(DP_mult_209_n279), .ZN(DP_mult_209_n2221) );
  XNOR2_X1 DP_mult_209_U2761 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2263), .ZN(
        DP_mult_209_n1713) );
  XNOR2_X1 DP_mult_209_U2760 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2263), .ZN(
        DP_mult_209_n1711) );
  XNOR2_X1 DP_mult_209_U2759 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2263), .ZN(
        DP_mult_209_n1719) );
  XNOR2_X1 DP_mult_209_U2758 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2262), .ZN(
        DP_mult_209_n1715) );
  XNOR2_X1 DP_mult_209_U2757 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2262), .ZN(
        DP_mult_209_n1709) );
  OAI22_X1 DP_mult_209_U2756 ( .A1(DP_mult_209_n2220), .A2(DP_mult_209_n1683), 
        .B1(DP_mult_209_n1682), .B2(DP_mult_209_n2246), .ZN(DP_mult_209_n836)
         );
  XNOR2_X1 DP_mult_209_U2755 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2262), .ZN(
        DP_mult_209_n1717) );
  OAI22_X1 DP_mult_209_U2754 ( .A1(DP_mult_209_n2220), .A2(DP_mult_209_n1693), 
        .B1(DP_mult_209_n1692), .B2(DP_mult_209_n2246), .ZN(DP_mult_209_n1396)
         );
  OAI22_X1 DP_mult_209_U2753 ( .A1(DP_mult_209_n2157), .A2(DP_mult_209_n2270), 
        .B1(DP_mult_209_n1706), .B2(DP_mult_209_n2245), .ZN(DP_mult_209_n1190)
         );
  OAI22_X1 DP_mult_209_U2752 ( .A1(DP_mult_209_n2158), .A2(DP_mult_209_n1684), 
        .B1(DP_mult_209_n2245), .B2(DP_mult_209_n1683), .ZN(DP_mult_209_n1387)
         );
  INV_X1 DP_mult_209_U2751 ( .A(DP_mult_209_n2027), .ZN(DP_mult_209_n837) );
  OAI22_X1 DP_mult_209_U2750 ( .A1(DP_mult_209_n2158), .A2(DP_mult_209_n1688), 
        .B1(DP_mult_209_n2245), .B2(DP_mult_209_n1687), .ZN(DP_mult_209_n1391)
         );
  OAI22_X1 DP_mult_209_U2749 ( .A1(DP_mult_209_n2158), .A2(DP_mult_209_n1685), 
        .B1(DP_mult_209_n1684), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1388)
         );
  OAI22_X1 DP_mult_209_U2748 ( .A1(DP_mult_209_n2157), .A2(DP_mult_209_n1692), 
        .B1(DP_mult_209_n2245), .B2(DP_mult_209_n1691), .ZN(DP_mult_209_n1395)
         );
  OAI22_X1 DP_mult_209_U2747 ( .A1(DP_mult_209_n2157), .A2(DP_mult_209_n1687), 
        .B1(DP_mult_209_n1686), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1390)
         );
  OAI22_X1 DP_mult_209_U2746 ( .A1(DP_mult_209_n2157), .A2(DP_mult_209_n1690), 
        .B1(DP_mult_209_n1993), .B2(DP_mult_209_n1689), .ZN(DP_mult_209_n1393)
         );
  OAI22_X1 DP_mult_209_U2745 ( .A1(DP_mult_209_n2158), .A2(DP_mult_209_n1689), 
        .B1(DP_mult_209_n1688), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1392)
         );
  OAI22_X1 DP_mult_209_U2744 ( .A1(DP_mult_209_n2023), .A2(DP_mult_209_n1686), 
        .B1(DP_mult_209_n2245), .B2(DP_mult_209_n1685), .ZN(DP_mult_209_n1389)
         );
  OAI22_X1 DP_mult_209_U2743 ( .A1(DP_mult_209_n2219), .A2(DP_mult_209_n1691), 
        .B1(DP_mult_209_n1690), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1394)
         );
  OAI21_X1 DP_mult_209_U2742 ( .B1(DP_mult_209_n2163), .B2(DP_mult_209_n398), 
        .A(DP_mult_209_n399), .ZN(DP_mult_209_n397) );
  OAI21_X1 DP_mult_209_U2741 ( .B1(DP_mult_209_n2162), .B2(DP_mult_209_n389), 
        .A(DP_mult_209_n390), .ZN(DP_mult_209_n388) );
  OAI21_X1 DP_mult_209_U2740 ( .B1(DP_mult_209_n2163), .B2(DP_mult_209_n431), 
        .A(DP_mult_209_n432), .ZN(DP_mult_209_n430) );
  OAI21_X1 DP_mult_209_U2739 ( .B1(DP_mult_209_n2162), .B2(DP_mult_209_n411), 
        .A(DP_mult_209_n412), .ZN(DP_mult_209_n410) );
  OAI21_X1 DP_mult_209_U2738 ( .B1(DP_mult_209_n301), .B2(DP_mult_209_n420), 
        .A(DP_mult_209_n421), .ZN(DP_mult_209_n419) );
  OAI21_X1 DP_mult_209_U2737 ( .B1(DP_mult_209_n301), .B2(DP_mult_209_n343), 
        .A(DP_mult_209_n344), .ZN(DP_mult_209_n342) );
  OAI21_X1 DP_mult_209_U2736 ( .B1(DP_mult_209_n2162), .B2(DP_mult_209_n380), 
        .A(DP_mult_209_n381), .ZN(DP_mult_209_n379) );
  OAI21_X1 DP_mult_209_U2735 ( .B1(DP_mult_209_n2163), .B2(DP_mult_209_n371), 
        .A(DP_mult_209_n372), .ZN(DP_mult_209_n370) );
  OAI21_X1 DP_mult_209_U2734 ( .B1(DP_mult_209_n301), .B2(DP_mult_209_n354), 
        .A(DP_mult_209_n355), .ZN(DP_mult_209_n353) );
  OAI21_X1 DP_mult_209_U2733 ( .B1(DP_mult_209_n2163), .B2(DP_mult_209_n438), 
        .A(DP_mult_209_n439), .ZN(DP_mult_209_n437) );
  INV_X1 DP_mult_209_U2732 ( .A(DP_mult_209_n2162), .ZN(DP_mult_209_n448) );
  OAI21_X1 DP_mult_209_U2731 ( .B1(DP_mult_209_n326), .B2(DP_mult_209_n301), 
        .A(DP_mult_209_n327), .ZN(DP_mult_209_n325) );
  XNOR2_X1 DP_mult_209_U2730 ( .A(DP_mult_209_n437), .B(DP_mult_209_n311), 
        .ZN(DP_pipe0_coeff_pipe03[13]) );
  XNOR2_X1 DP_mult_209_U2729 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2284), .ZN(
        DP_mult_209_n1584) );
  XNOR2_X1 DP_mult_209_U2728 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2284), .ZN(
        DP_mult_209_n1586) );
  XNOR2_X1 DP_mult_209_U2727 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2284), .ZN(
        DP_mult_209_n1594) );
  OAI22_X1 DP_mult_209_U2726 ( .A1(DP_mult_209_n1962), .A2(DP_mult_209_n1558), 
        .B1(DP_mult_209_n1557), .B2(DP_mult_209_n2230), .ZN(DP_mult_209_n706)
         );
  XNOR2_X1 DP_mult_209_U2725 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2284), .ZN(
        DP_mult_209_n1590) );
  XNOR2_X1 DP_mult_209_U2724 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2284), .ZN(
        DP_mult_209_n1592) );
  XNOR2_X1 DP_mult_209_U2723 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2284), .ZN(
        DP_mult_209_n1588) );
  OAI22_X1 DP_mult_209_U2722 ( .A1(DP_mult_209_n2210), .A2(DP_mult_209_n1562), 
        .B1(DP_mult_209_n1561), .B2(DP_mult_209_n2230), .ZN(DP_mult_209_n1270)
         );
  OAI22_X1 DP_mult_209_U2721 ( .A1(DP_mult_209_n2209), .A2(DP_mult_209_n1568), 
        .B1(DP_mult_209_n1567), .B2(DP_mult_209_n2231), .ZN(DP_mult_209_n1276)
         );
  OAI22_X1 DP_mult_209_U2720 ( .A1(DP_mult_209_n2210), .A2(DP_mult_209_n2292), 
        .B1(DP_mult_209_n1581), .B2(DP_mult_209_n2230), .ZN(DP_mult_209_n1185)
         );
  OAI22_X1 DP_mult_209_U2719 ( .A1(DP_mult_209_n1962), .A2(DP_mult_209_n1559), 
        .B1(DP_mult_209_n2230), .B2(DP_mult_209_n1558), .ZN(DP_mult_209_n1267)
         );
  OAI22_X1 DP_mult_209_U2718 ( .A1(DP_mult_209_n1962), .A2(DP_mult_209_n1560), 
        .B1(DP_mult_209_n1559), .B2(DP_mult_209_n2230), .ZN(DP_mult_209_n1268)
         );
  OAI22_X1 DP_mult_209_U2717 ( .A1(DP_mult_209_n2210), .A2(DP_mult_209_n1565), 
        .B1(DP_mult_209_n2230), .B2(DP_mult_209_n1564), .ZN(DP_mult_209_n1273)
         );
  OAI22_X1 DP_mult_209_U2716 ( .A1(DP_mult_209_n1963), .A2(DP_mult_209_n1561), 
        .B1(DP_mult_209_n2230), .B2(DP_mult_209_n1560), .ZN(DP_mult_209_n1269)
         );
  OAI22_X1 DP_mult_209_U2715 ( .A1(DP_mult_209_n1963), .A2(DP_mult_209_n1564), 
        .B1(DP_mult_209_n1563), .B2(DP_mult_209_n2230), .ZN(DP_mult_209_n1272)
         );
  OAI22_X1 DP_mult_209_U2714 ( .A1(DP_mult_209_n1962), .A2(DP_mult_209_n1566), 
        .B1(DP_mult_209_n1565), .B2(DP_mult_209_n2230), .ZN(DP_mult_209_n1274)
         );
  OAI22_X1 DP_mult_209_U2713 ( .A1(DP_mult_209_n1963), .A2(DP_mult_209_n1567), 
        .B1(DP_mult_209_n2230), .B2(DP_mult_209_n1566), .ZN(DP_mult_209_n1275)
         );
  OAI22_X1 DP_mult_209_U2712 ( .A1(DP_mult_209_n1963), .A2(DP_mult_209_n1563), 
        .B1(DP_mult_209_n2230), .B2(DP_mult_209_n1562), .ZN(DP_mult_209_n1271)
         );
  NAND2_X1 DP_mult_209_U2711 ( .A1(DP_mult_209_n694), .A2(DP_mult_209_n689), 
        .ZN(DP_mult_209_n378) );
  NAND2_X1 DP_mult_209_U2710 ( .A1(DP_mult_209_n2177), .A2(DP_mult_209_n2179), 
        .ZN(DP_mult_209_n364) );
  NAND2_X1 DP_mult_209_U2709 ( .A1(DP_mult_209_n382), .A2(DP_mult_209_n2177), 
        .ZN(DP_mult_209_n371) );
  AOI21_X1 DP_mult_209_U2708 ( .B1(DP_mult_209_n383), .B2(DP_mult_209_n2177), 
        .A(DP_mult_209_n376), .ZN(DP_mult_209_n372) );
  NAND2_X1 DP_mult_209_U2707 ( .A1(DP_mult_209_n2177), .A2(DP_mult_209_n378), 
        .ZN(DP_mult_209_n305) );
  INV_X1 DP_mult_209_U2706 ( .A(DP_mult_209_n325), .ZN(
        DP_pipe0_coeff_pipe03[23]) );
  NAND2_X1 DP_mult_209_U2705 ( .A1(DP_mult_209_n1815), .A2(DP_mult_209_n2067), 
        .ZN(DP_mult_209_n279) );
  XNOR2_X1 DP_mult_209_U2704 ( .A(DP_pipe03[13]), .B(DP_mult_209_n1940), .ZN(
        DP_mult_209_n1742) );
  XNOR2_X1 DP_mult_209_U2703 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2258), .ZN(
        DP_mult_209_n1738) );
  XNOR2_X1 DP_mult_209_U2702 ( .A(DP_pipe03[11]), .B(DP_mult_209_n1941), .ZN(
        DP_mult_209_n1744) );
  XNOR2_X1 DP_mult_209_U2701 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2258), .ZN(
        DP_mult_209_n1736) );
  XNOR2_X1 DP_mult_209_U2700 ( .A(DP_pipe03[15]), .B(DP_mult_209_n1941), .ZN(
        DP_mult_209_n1740) );
  OAI22_X1 DP_mult_209_U2699 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1724), 
        .B1(DP_mult_209_n1723), .B2(DP_mult_209_n2247), .ZN(DP_mult_209_n1426)
         );
  XNOR2_X1 DP_mult_209_U2698 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2258), .ZN(
        DP_mult_209_n1734) );
  OAI22_X1 DP_mult_209_U2697 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1714), 
        .B1(DP_mult_209_n1713), .B2(DP_mult_209_n2247), .ZN(DP_mult_209_n1416)
         );
  OAI22_X1 DP_mult_209_U2696 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1719), 
        .B1(DP_mult_209_n1959), .B2(DP_mult_209_n1718), .ZN(DP_mult_209_n1421)
         );
  OAI22_X1 DP_mult_209_U2695 ( .A1(DP_mult_209_n2193), .A2(DP_mult_209_n1716), 
        .B1(DP_mult_209_n1715), .B2(DP_mult_209_n1958), .ZN(DP_mult_209_n1418)
         );
  OAI22_X1 DP_mult_209_U2694 ( .A1(DP_mult_209_n2089), .A2(DP_mult_209_n1712), 
        .B1(DP_mult_209_n1711), .B2(DP_mult_209_n1959), .ZN(DP_mult_209_n1414)
         );
  OAI22_X1 DP_mult_209_U2693 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1722), 
        .B1(DP_mult_209_n1721), .B2(DP_mult_209_n1958), .ZN(DP_mult_209_n1424)
         );
  OAI22_X1 DP_mult_209_U2692 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1729), 
        .B1(DP_mult_209_n1958), .B2(DP_mult_209_n1728), .ZN(DP_mult_209_n1431)
         );
  OAI22_X1 DP_mult_209_U2691 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1728), 
        .B1(DP_mult_209_n1727), .B2(DP_mult_209_n1959), .ZN(DP_mult_209_n1430)
         );
  OAI22_X1 DP_mult_209_U2690 ( .A1(DP_mult_209_n2193), .A2(DP_mult_209_n1710), 
        .B1(DP_mult_209_n1709), .B2(DP_mult_209_n1958), .ZN(DP_mult_209_n1412)
         );
  OAI22_X1 DP_mult_209_U2689 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1723), 
        .B1(DP_mult_209_n1958), .B2(DP_mult_209_n1722), .ZN(DP_mult_209_n1425)
         );
  OAI22_X1 DP_mult_209_U2688 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1725), 
        .B1(DP_mult_209_n1959), .B2(DP_mult_209_n1724), .ZN(DP_mult_209_n1427)
         );
  OAI22_X1 DP_mult_209_U2687 ( .A1(DP_mult_209_n2089), .A2(DP_mult_209_n1708), 
        .B1(DP_mult_209_n1707), .B2(DP_mult_209_n2247), .ZN(DP_mult_209_n874)
         );
  OAI22_X1 DP_mult_209_U2686 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1730), 
        .B1(DP_mult_209_n1729), .B2(DP_mult_209_n1959), .ZN(DP_mult_209_n1432)
         );
  OAI22_X1 DP_mult_209_U2685 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1726), 
        .B1(DP_mult_209_n1725), .B2(DP_mult_209_n1958), .ZN(DP_mult_209_n1428)
         );
  OAI22_X1 DP_mult_209_U2684 ( .A1(DP_mult_209_n2089), .A2(DP_mult_209_n1718), 
        .B1(DP_mult_209_n1717), .B2(DP_mult_209_n1958), .ZN(DP_mult_209_n1420)
         );
  OAI22_X1 DP_mult_209_U2683 ( .A1(DP_mult_209_n2193), .A2(DP_mult_209_n2264), 
        .B1(DP_mult_209_n1731), .B2(DP_mult_209_n1959), .ZN(DP_mult_209_n1191)
         );
  OAI22_X1 DP_mult_209_U2682 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1721), 
        .B1(DP_mult_209_n1959), .B2(DP_mult_209_n1720), .ZN(DP_mult_209_n1423)
         );
  OAI22_X1 DP_mult_209_U2681 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1720), 
        .B1(DP_mult_209_n1719), .B2(DP_mult_209_n1958), .ZN(DP_mult_209_n1422)
         );
  OAI22_X1 DP_mult_209_U2680 ( .A1(DP_mult_209_n2022), .A2(DP_mult_209_n1727), 
        .B1(DP_mult_209_n1959), .B2(DP_mult_209_n1726), .ZN(DP_mult_209_n1429)
         );
  OAI21_X1 DP_mult_209_U2679 ( .B1(DP_mult_209_n1951), .B2(DP_mult_209_n498), 
        .A(DP_mult_209_n499), .ZN(DP_mult_209_n497) );
  OAI21_X1 DP_mult_209_U2678 ( .B1(DP_mult_209_n1950), .B2(DP_mult_209_n487), 
        .A(DP_mult_209_n488), .ZN(DP_mult_209_n486) );
  OAI21_X1 DP_mult_209_U2677 ( .B1(DP_mult_209_n1949), .B2(DP_mult_209_n476), 
        .A(DP_mult_209_n477), .ZN(DP_mult_209_n475) );
  OAI21_X1 DP_mult_209_U2676 ( .B1(DP_mult_209_n1949), .B2(DP_mult_209_n2150), 
        .A(DP_mult_209_n524), .ZN(DP_mult_209_n522) );
  OAI21_X1 DP_mult_209_U2675 ( .B1(DP_mult_209_n1951), .B2(DP_mult_209_n463), 
        .A(DP_mult_209_n464), .ZN(DP_mult_209_n462) );
  OAI21_X1 DP_mult_209_U2674 ( .B1(DP_mult_209_n1951), .B2(DP_mult_209_n2151), 
        .A(DP_mult_209_n535), .ZN(DP_mult_209_n533) );
  OAI21_X1 DP_mult_209_U2673 ( .B1(DP_mult_209_n1950), .B2(DP_mult_209_n516), 
        .A(DP_mult_209_n517), .ZN(DP_mult_209_n515) );
  OAI21_X1 DP_mult_209_U2672 ( .B1(DP_mult_209_n1949), .B2(DP_mult_209_n2136), 
        .A(DP_mult_209_n2197), .ZN(DP_mult_209_n504) );
  XNOR2_X1 DP_mult_209_U2671 ( .A(DP_mult_209_n533), .B(DP_mult_209_n320), 
        .ZN(DP_pipe0_coeff_pipe03[4]) );
  XNOR2_X1 DP_mult_209_U2670 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1642) );
  XNOR2_X1 DP_mult_209_U2669 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1640) );
  XNOR2_X1 DP_mult_209_U2668 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1638) );
  XNOR2_X1 DP_mult_209_U2667 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1644) );
  OAI22_X1 DP_mult_209_U2666 ( .A1(DP_mult_209_n1991), .A2(DP_mult_209_n1608), 
        .B1(DP_mult_209_n1607), .B2(DP_mult_209_n2238), .ZN(DP_mult_209_n746)
         );
  XNOR2_X1 DP_mult_209_U2665 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1634) );
  XNOR2_X1 DP_mult_209_U2664 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1636) );
  OAI22_X1 DP_mult_209_U2663 ( .A1(DP_mult_209_n2213), .A2(DP_mult_209_n1614), 
        .B1(DP_mult_209_n1613), .B2(DP_mult_209_n2238), .ZN(DP_mult_209_n1320)
         );
  OAI22_X1 DP_mult_209_U2662 ( .A1(DP_mult_209_n1991), .A2(DP_mult_209_n1618), 
        .B1(DP_mult_209_n1617), .B2(DP_mult_209_n2238), .ZN(DP_mult_209_n1324)
         );
  OAI22_X1 DP_mult_209_U2661 ( .A1(DP_mult_209_n2011), .A2(DP_mult_209_n1609), 
        .B1(DP_mult_209_n2238), .B2(DP_mult_209_n1608), .ZN(DP_mult_209_n1315)
         );
  OAI22_X1 DP_mult_209_U2660 ( .A1(DP_mult_209_n1992), .A2(DP_mult_209_n1616), 
        .B1(DP_mult_209_n1615), .B2(DP_mult_209_n2238), .ZN(DP_mult_209_n1322)
         );
  INV_X1 DP_mult_209_U2659 ( .A(DP_mult_209_n746), .ZN(DP_mult_209_n747) );
  OAI22_X1 DP_mult_209_U2658 ( .A1(DP_mult_209_n2213), .A2(DP_mult_209_n1615), 
        .B1(DP_mult_209_n2237), .B2(DP_mult_209_n1614), .ZN(DP_mult_209_n1321)
         );
  OAI22_X1 DP_mult_209_U2657 ( .A1(DP_mult_209_n2213), .A2(DP_mult_209_n1611), 
        .B1(DP_mult_209_n2237), .B2(DP_mult_209_n1610), .ZN(DP_mult_209_n1317)
         );
  OAI22_X1 DP_mult_209_U2656 ( .A1(DP_mult_209_n1992), .A2(DP_mult_209_n2282), 
        .B1(DP_mult_209_n1631), .B2(DP_mult_209_n2237), .ZN(DP_mult_209_n1187)
         );
  OAI22_X1 DP_mult_209_U2655 ( .A1(DP_mult_209_n2213), .A2(DP_mult_209_n1617), 
        .B1(DP_mult_209_n2238), .B2(DP_mult_209_n1616), .ZN(DP_mult_209_n1323)
         );
  OAI22_X1 DP_mult_209_U2654 ( .A1(DP_mult_209_n2011), .A2(DP_mult_209_n1612), 
        .B1(DP_mult_209_n1611), .B2(DP_mult_209_n2238), .ZN(DP_mult_209_n1318)
         );
  OAI22_X1 DP_mult_209_U2653 ( .A1(DP_mult_209_n1991), .A2(DP_mult_209_n1613), 
        .B1(DP_mult_209_n2238), .B2(DP_mult_209_n1612), .ZN(DP_mult_209_n1319)
         );
  OAI22_X1 DP_mult_209_U2652 ( .A1(DP_mult_209_n2011), .A2(DP_mult_209_n1610), 
        .B1(DP_mult_209_n1609), .B2(DP_mult_209_n2237), .ZN(DP_mult_209_n1316)
         );
  NAND2_X1 DP_mult_209_U2651 ( .A1(DP_mult_209_n717), .A2(DP_mult_209_n726), 
        .ZN(DP_mult_209_n418) );
  AOI21_X1 DP_mult_209_U2650 ( .B1(DP_mult_209_n346), .B2(DP_mult_209_n2181), 
        .A(DP_mult_209_n339), .ZN(DP_mult_209_n337) );
  INV_X1 DP_mult_209_U2649 ( .A(DP_mult_209_n346), .ZN(DP_mult_209_n344) );
  OAI21_X1 DP_mult_209_U2648 ( .B1(DP_mult_209_n506), .B2(DP_mult_209_n452), 
        .A(DP_mult_209_n453), .ZN(DP_mult_209_n451) );
  OAI22_X1 DP_mult_209_U2647 ( .A1(DP_mult_209_n2222), .A2(DP_mult_209_n1733), 
        .B1(DP_mult_209_n1732), .B2(DP_mult_209_n2248), .ZN(DP_mult_209_n916)
         );
  XNOR2_X1 DP_mult_209_U2646 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2036), .ZN(
        DP_mult_209_n1613) );
  XNOR2_X1 DP_mult_209_U2645 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2036), .ZN(
        DP_mult_209_n1615) );
  XNOR2_X1 DP_mult_209_U2644 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2036), .ZN(
        DP_mult_209_n1619) );
  OAI22_X1 DP_mult_209_U2643 ( .A1(DP_mult_209_n2155), .A2(DP_mult_209_n1605), 
        .B1(DP_mult_209_n1604), .B2(DP_mult_209_n2235), .ZN(DP_mult_209_n1312)
         );
  XNOR2_X1 DP_mult_209_U2642 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2035), .ZN(
        DP_mult_209_n1617) );
  XNOR2_X1 DP_mult_209_U2641 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2035), .ZN(
        DP_mult_209_n1611) );
  OAI22_X1 DP_mult_209_U2640 ( .A1(DP_mult_209_n2156), .A2(DP_mult_209_n1604), 
        .B1(DP_mult_209_n2234), .B2(DP_mult_209_n1603), .ZN(DP_mult_209_n1311)
         );
  XNOR2_X1 DP_mult_209_U2639 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2036), .ZN(
        DP_mult_209_n1609) );
  OAI22_X1 DP_mult_209_U2638 ( .A1(DP_mult_209_n2155), .A2(DP_mult_209_n1599), 
        .B1(DP_mult_209_n1598), .B2(DP_mult_209_n2234), .ZN(DP_mult_209_n1306)
         );
  OAI22_X1 DP_mult_209_U2637 ( .A1(DP_mult_209_n2212), .A2(DP_mult_209_n1603), 
        .B1(DP_mult_209_n1602), .B2(DP_mult_209_n2234), .ZN(DP_mult_209_n1310)
         );
  OAI22_X1 DP_mult_209_U2636 ( .A1(DP_mult_209_n2211), .A2(DP_mult_209_n1595), 
        .B1(DP_mult_209_n1594), .B2(DP_mult_209_n2234), .ZN(DP_mult_209_n1302)
         );
  OAI22_X1 DP_mult_209_U2635 ( .A1(DP_mult_209_n2212), .A2(DP_mult_209_n1598), 
        .B1(DP_mult_209_n2234), .B2(DP_mult_209_n1597), .ZN(DP_mult_209_n1305)
         );
  OAI22_X1 DP_mult_209_U2634 ( .A1(DP_mult_209_n2212), .A2(DP_mult_209_n1597), 
        .B1(DP_mult_209_n1596), .B2(DP_mult_209_n2235), .ZN(DP_mult_209_n1304)
         );
  OAI22_X1 DP_mult_209_U2633 ( .A1(DP_mult_209_n2156), .A2(DP_mult_209_n1601), 
        .B1(DP_mult_209_n1600), .B2(DP_mult_209_n2234), .ZN(DP_mult_209_n1308)
         );
  OAI22_X1 DP_mult_209_U2632 ( .A1(DP_mult_209_n2211), .A2(DP_mult_209_n1600), 
        .B1(DP_mult_209_n2235), .B2(DP_mult_209_n1599), .ZN(DP_mult_209_n1307)
         );
  OAI22_X1 DP_mult_209_U2631 ( .A1(DP_mult_209_n2211), .A2(DP_mult_209_n1596), 
        .B1(DP_mult_209_n2235), .B2(DP_mult_209_n1595), .ZN(DP_mult_209_n1303)
         );
  OAI22_X1 DP_mult_209_U2630 ( .A1(DP_mult_209_n2155), .A2(DP_mult_209_n1602), 
        .B1(DP_mult_209_n2235), .B2(DP_mult_209_n1601), .ZN(DP_mult_209_n1309)
         );
  OAI22_X1 DP_mult_209_U2629 ( .A1(DP_mult_209_n2156), .A2(DP_mult_209_n1594), 
        .B1(DP_mult_209_n2234), .B2(DP_mult_209_n1593), .ZN(DP_mult_209_n1301)
         );
  OAI21_X1 DP_mult_209_U2628 ( .B1(DP_mult_209_n572), .B2(DP_mult_209_n569), 
        .A(DP_mult_209_n570), .ZN(DP_mult_209_n568) );
  XNOR2_X1 DP_mult_209_U2627 ( .A(DP_mult_209_n430), .B(DP_mult_209_n310), 
        .ZN(DP_pipe0_coeff_pipe03[14]) );
  AOI21_X1 DP_mult_209_U2626 ( .B1(DP_mult_209_n490), .B2(DP_mult_209_n454), 
        .A(DP_mult_209_n455), .ZN(DP_mult_209_n453) );
  NAND2_X1 DP_mult_209_U2625 ( .A1(DP_mult_209_n454), .A2(DP_mult_209_n489), 
        .ZN(DP_mult_209_n452) );
  OAI22_X1 DP_mult_209_U2624 ( .A1(DP_mult_209_n2096), .A2(DP_mult_209_n1553), 
        .B1(DP_mult_209_n1552), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1262)
         );
  OAI22_X1 DP_mult_209_U2623 ( .A1(DP_mult_209_n2097), .A2(DP_mult_209_n1554), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1553), .ZN(DP_mult_209_n1263)
         );
  OAI22_X1 DP_mult_209_U2622 ( .A1(DP_mult_209_n2096), .A2(DP_mult_209_n1551), 
        .B1(DP_mult_209_n1550), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1260)
         );
  OAI22_X1 DP_mult_209_U2621 ( .A1(DP_mult_209_n2208), .A2(DP_mult_209_n1550), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1549), .ZN(DP_mult_209_n1259)
         );
  OAI22_X1 DP_mult_209_U2620 ( .A1(DP_mult_209_n2208), .A2(DP_mult_209_n1555), 
        .B1(DP_mult_209_n1554), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1264)
         );
  OAI22_X1 DP_mult_209_U2619 ( .A1(DP_mult_209_n2096), .A2(DP_mult_209_n1547), 
        .B1(DP_mult_209_n1546), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1256)
         );
  OAI22_X1 DP_mult_209_U2618 ( .A1(DP_mult_209_n2096), .A2(DP_mult_209_n1545), 
        .B1(DP_mult_209_n1544), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1254)
         );
  OAI22_X1 DP_mult_209_U2617 ( .A1(DP_mult_209_n2207), .A2(DP_mult_209_n1549), 
        .B1(DP_mult_209_n1548), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1258)
         );
  OAI22_X1 DP_mult_209_U2616 ( .A1(DP_mult_209_n2097), .A2(DP_mult_209_n1552), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1551), .ZN(DP_mult_209_n1261)
         );
  OAI22_X1 DP_mult_209_U2615 ( .A1(DP_mult_209_n2097), .A2(DP_mult_209_n1548), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1547), .ZN(DP_mult_209_n1257)
         );
  OAI22_X1 DP_mult_209_U2614 ( .A1(DP_mult_209_n2208), .A2(DP_mult_209_n1546), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1545), .ZN(DP_mult_209_n1255)
         );
  OAI22_X1 DP_mult_209_U2613 ( .A1(DP_mult_209_n2207), .A2(DP_mult_209_n1544), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1543), .ZN(DP_mult_209_n1253)
         );
  XNOR2_X1 DP_mult_209_U2612 ( .A(DP_mult_209_n419), .B(DP_mult_209_n309), 
        .ZN(DP_pipe0_coeff_pipe03[15]) );
  OAI22_X1 DP_mult_209_U2611 ( .A1(DP_mult_209_n2215), .A2(DP_mult_209_n1646), 
        .B1(DP_mult_209_n2240), .B2(DP_mult_209_n1645), .ZN(DP_mult_209_n1351)
         );
  OAI22_X1 DP_mult_209_U2610 ( .A1(DP_mult_209_n2160), .A2(DP_mult_209_n1655), 
        .B1(DP_mult_209_n1654), .B2(DP_mult_209_n2240), .ZN(DP_mult_209_n1360)
         );
  OAI22_X1 DP_mult_209_U2609 ( .A1(DP_mult_209_n2024), .A2(DP_mult_209_n1654), 
        .B1(DP_mult_209_n2241), .B2(DP_mult_209_n1653), .ZN(DP_mult_209_n1359)
         );
  OAI22_X1 DP_mult_209_U2608 ( .A1(DP_mult_209_n2025), .A2(DP_mult_209_n1644), 
        .B1(DP_mult_209_n2240), .B2(DP_mult_209_n1643), .ZN(DP_mult_209_n1349)
         );
  OAI22_X1 DP_mult_209_U2607 ( .A1(DP_mult_209_n2215), .A2(DP_mult_209_n1645), 
        .B1(DP_mult_209_n1644), .B2(DP_mult_209_n2240), .ZN(DP_mult_209_n1350)
         );
  OAI22_X1 DP_mult_209_U2606 ( .A1(DP_mult_209_n2216), .A2(DP_mult_209_n1650), 
        .B1(DP_mult_209_n2240), .B2(DP_mult_209_n1649), .ZN(DP_mult_209_n1355)
         );
  OAI22_X1 DP_mult_209_U2605 ( .A1(DP_mult_209_n2160), .A2(DP_mult_209_n1647), 
        .B1(DP_mult_209_n1646), .B2(DP_mult_209_n2240), .ZN(DP_mult_209_n1352)
         );
  OAI22_X1 DP_mult_209_U2604 ( .A1(DP_mult_209_n2025), .A2(DP_mult_209_n1653), 
        .B1(DP_mult_209_n1652), .B2(DP_mult_209_n2240), .ZN(DP_mult_209_n1358)
         );
  OAI22_X1 DP_mult_209_U2603 ( .A1(DP_mult_209_n2216), .A2(DP_mult_209_n1648), 
        .B1(DP_mult_209_n2241), .B2(DP_mult_209_n1647), .ZN(DP_mult_209_n1353)
         );
  OAI22_X1 DP_mult_209_U2602 ( .A1(DP_mult_209_n2160), .A2(DP_mult_209_n1652), 
        .B1(DP_mult_209_n2240), .B2(DP_mult_209_n1651), .ZN(DP_mult_209_n1357)
         );
  OAI22_X1 DP_mult_209_U2601 ( .A1(DP_mult_209_n2216), .A2(DP_mult_209_n1649), 
        .B1(DP_mult_209_n1648), .B2(DP_mult_209_n2241), .ZN(DP_mult_209_n1354)
         );
  NAND2_X1 DP_mult_209_U2600 ( .A1(DP_mult_209_n1071), .A2(DP_mult_209_n1084), 
        .ZN(DP_mult_209_n591) );
  XNOR2_X1 DP_mult_209_U2599 ( .A(DP_mult_209_n410), .B(DP_mult_209_n308), 
        .ZN(DP_pipe0_coeff_pipe03[16]) );
  XNOR2_X1 DP_mult_209_U2598 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2295), .ZN(
        DP_mult_209_n1538) );
  XNOR2_X1 DP_mult_209_U2597 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2295), .ZN(
        DP_mult_209_n1540) );
  XNOR2_X1 DP_mult_209_U2596 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2295), .ZN(
        DP_mult_209_n1544) );
  XNOR2_X1 DP_mult_209_U2595 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2295), .ZN(
        DP_mult_209_n1542) );
  OAI22_X1 DP_mult_209_U2594 ( .A1(DP_mult_209_n2014), .A2(DP_mult_209_n1527), 
        .B1(DP_mult_209_n2227), .B2(DP_mult_209_n1526), .ZN(DP_mult_209_n1237)
         );
  OAI22_X1 DP_mult_209_U2593 ( .A1(DP_mult_209_n1954), .A2(DP_mult_209_n1530), 
        .B1(DP_mult_209_n1529), .B2(DP_mult_209_n2228), .ZN(DP_mult_209_n1240)
         );
  XNOR2_X1 DP_mult_209_U2592 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2295), .ZN(
        DP_mult_209_n1536) );
  OAI22_X1 DP_mult_209_U2591 ( .A1(DP_mult_209_n2014), .A2(DP_mult_209_n1528), 
        .B1(DP_mult_209_n1527), .B2(DP_mult_209_n2228), .ZN(DP_mult_209_n1238)
         );
  OAI22_X1 DP_mult_209_U2590 ( .A1(DP_mult_209_n2102), .A2(DP_mult_209_n1529), 
        .B1(DP_mult_209_n2227), .B2(DP_mult_209_n1528), .ZN(DP_mult_209_n1239)
         );
  OAI22_X1 DP_mult_209_U2589 ( .A1(DP_mult_209_n1524), .A2(DP_mult_209_n2015), 
        .B1(DP_mult_209_n1523), .B2(DP_mult_209_n2228), .ZN(DP_mult_209_n1234)
         );
  OAI22_X1 DP_mult_209_U2588 ( .A1(DP_mult_209_n2206), .A2(DP_mult_209_n1526), 
        .B1(DP_mult_209_n1525), .B2(DP_mult_209_n2227), .ZN(DP_mult_209_n1236)
         );
  XNOR2_X1 DP_mult_209_U2587 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2295), .ZN(
        DP_mult_209_n1534) );
  OAI22_X1 DP_mult_209_U2586 ( .A1(DP_mult_209_n2102), .A2(DP_mult_209_n1523), 
        .B1(DP_mult_209_n2228), .B2(DP_mult_209_n1522), .ZN(DP_mult_209_n1233)
         );
  OAI22_X1 DP_mult_209_U2585 ( .A1(DP_mult_209_n2102), .A2(DP_mult_209_n1525), 
        .B1(DP_mult_209_n2228), .B2(DP_mult_209_n1524), .ZN(DP_mult_209_n1235)
         );
  OAI22_X1 DP_mult_209_U2584 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1519), 
        .B1(DP_mult_209_n2228), .B2(DP_mult_209_n1518), .ZN(DP_mult_209_n1229)
         );
  OAI22_X1 DP_mult_209_U2583 ( .A1(DP_mult_209_n2015), .A2(DP_mult_209_n1520), 
        .B1(DP_mult_209_n1519), .B2(DP_mult_209_n2227), .ZN(DP_mult_209_n1230)
         );
  OAI22_X1 DP_mult_209_U2582 ( .A1(DP_mult_209_n2206), .A2(DP_mult_209_n1521), 
        .B1(DP_mult_209_n2227), .B2(DP_mult_209_n1520), .ZN(DP_mult_209_n1231)
         );
  OAI22_X1 DP_mult_209_U2581 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1522), 
        .B1(DP_mult_209_n1521), .B2(DP_mult_209_n2228), .ZN(DP_mult_209_n1232)
         );
  XNOR2_X1 DP_mult_209_U2580 ( .A(DP_coeffs_ff_int[87]), .B(
        DP_coeffs_ff_int[88]), .ZN(DP_mult_209_n259) );
  XNOR2_X1 DP_mult_209_U2579 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2268), .ZN(
        DP_mult_209_n1692) );
  XNOR2_X1 DP_mult_209_U2578 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2268), .ZN(
        DP_mult_209_n1694) );
  XNOR2_X1 DP_mult_209_U2577 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2268), .ZN(
        DP_mult_209_n1684) );
  XNOR2_X1 DP_mult_209_U2576 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2268), .ZN(
        DP_mult_209_n1690) );
  XNOR2_X1 DP_mult_209_U2575 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2267), .ZN(
        DP_mult_209_n1686) );
  OAI22_X1 DP_mult_209_U2574 ( .A1(DP_mult_209_n1668), .A2(DP_mult_209_n2217), 
        .B1(DP_mult_209_n1667), .B2(DP_mult_209_n2242), .ZN(DP_mult_209_n1372)
         );
  XNOR2_X1 DP_mult_209_U2573 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2268), .ZN(
        DP_mult_209_n1688) );
  OAI22_X1 DP_mult_209_U2572 ( .A1(DP_mult_209_n2217), .A2(DP_mult_209_n1659), 
        .B1(DP_mult_209_n2242), .B2(DP_mult_209_n1658), .ZN(DP_mult_209_n1363)
         );
  OAI22_X1 DP_mult_209_U2571 ( .A1(DP_mult_209_n2217), .A2(DP_mult_209_n1666), 
        .B1(DP_mult_209_n1665), .B2(DP_mult_209_n2243), .ZN(DP_mult_209_n1370)
         );
  OAI22_X1 DP_mult_209_U2570 ( .A1(DP_mult_209_n2192), .A2(DP_mult_209_n1662), 
        .B1(DP_mult_209_n1661), .B2(DP_mult_209_n2242), .ZN(DP_mult_209_n1366)
         );
  OAI22_X1 DP_mult_209_U2569 ( .A1(DP_mult_209_n2192), .A2(DP_mult_209_n1665), 
        .B1(DP_mult_209_n2243), .B2(DP_mult_209_n1664), .ZN(DP_mult_209_n1369)
         );
  OAI22_X1 DP_mult_209_U2568 ( .A1(DP_mult_209_n2217), .A2(DP_mult_209_n1658), 
        .B1(DP_mult_209_n1657), .B2(DP_mult_209_n2243), .ZN(DP_mult_209_n802)
         );
  OAI22_X1 DP_mult_209_U2567 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1667), 
        .B1(DP_mult_209_n2243), .B2(DP_mult_209_n1666), .ZN(DP_mult_209_n1371)
         );
  OAI22_X1 DP_mult_209_U2566 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1664), 
        .B1(DP_mult_209_n1663), .B2(DP_mult_209_n2242), .ZN(DP_mult_209_n1368)
         );
  OAI22_X1 DP_mult_209_U2565 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1988), 
        .B1(DP_mult_209_n1681), .B2(DP_mult_209_n2242), .ZN(DP_mult_209_n1189)
         );
  OAI22_X1 DP_mult_209_U2564 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1663), 
        .B1(DP_mult_209_n2243), .B2(DP_mult_209_n1662), .ZN(DP_mult_209_n1367)
         );
  OAI22_X1 DP_mult_209_U2563 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1660), 
        .B1(DP_mult_209_n1659), .B2(DP_mult_209_n2242), .ZN(DP_mult_209_n1364)
         );
  OAI22_X1 DP_mult_209_U2562 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1661), 
        .B1(DP_mult_209_n2242), .B2(DP_mult_209_n1660), .ZN(DP_mult_209_n1365)
         );
  XNOR2_X1 DP_mult_209_U2561 ( .A(DP_mult_209_n397), .B(DP_mult_209_n307), 
        .ZN(DP_pipe0_coeff_pipe03[17]) );
  NAND2_X1 DP_mult_209_U2560 ( .A1(DP_mult_209_n332), .A2(DP_mult_209_n2182), 
        .ZN(DP_mult_209_n326) );
  OAI22_X1 DP_mult_209_U2559 ( .A1(DP_mult_209_n2194), .A2(DP_mult_209_n1755), 
        .B1(DP_mult_209_n1754), .B2(DP_mult_209_n2248), .ZN(DP_mult_209_n1456)
         );
  OAI22_X1 DP_mult_209_U2558 ( .A1(DP_mult_209_n2222), .A2(DP_mult_209_n1751), 
        .B1(DP_mult_209_n1750), .B2(DP_mult_209_n2248), .ZN(DP_mult_209_n1452)
         );
  OAI22_X1 DP_mult_209_U2557 ( .A1(DP_mult_209_n2222), .A2(DP_mult_209_n1752), 
        .B1(DP_mult_209_n2019), .B2(DP_mult_209_n1751), .ZN(DP_mult_209_n1453)
         );
  OAI22_X1 DP_mult_209_U2556 ( .A1(DP_mult_209_n2195), .A2(DP_mult_209_n1754), 
        .B1(DP_mult_209_n2248), .B2(DP_mult_209_n1753), .ZN(DP_mult_209_n1455)
         );
  OAI22_X1 DP_mult_209_U2555 ( .A1(DP_mult_209_n2222), .A2(DP_mult_209_n1746), 
        .B1(DP_mult_209_n2248), .B2(DP_mult_209_n1745), .ZN(DP_mult_209_n1447)
         );
  OAI22_X1 DP_mult_209_U2554 ( .A1(DP_mult_209_n2196), .A2(DP_mult_209_n1744), 
        .B1(DP_mult_209_n2248), .B2(DP_mult_209_n1743), .ZN(DP_mult_209_n1445)
         );
  OAI22_X1 DP_mult_209_U2553 ( .A1(DP_mult_209_n2195), .A2(DP_mult_209_n1748), 
        .B1(DP_mult_209_n2019), .B2(DP_mult_209_n1747), .ZN(DP_mult_209_n1449)
         );
  OAI22_X1 DP_mult_209_U2552 ( .A1(DP_mult_209_n2196), .A2(DP_mult_209_n1745), 
        .B1(DP_mult_209_n1744), .B2(DP_mult_209_n2019), .ZN(DP_mult_209_n1446)
         );
  OAI22_X1 DP_mult_209_U2551 ( .A1(DP_mult_209_n2194), .A2(DP_mult_209_n1749), 
        .B1(DP_mult_209_n1748), .B2(DP_mult_209_n2019), .ZN(DP_mult_209_n1450)
         );
  OAI22_X1 DP_mult_209_U2550 ( .A1(DP_mult_209_n2194), .A2(DP_mult_209_n1750), 
        .B1(DP_mult_209_n2248), .B2(DP_mult_209_n1749), .ZN(DP_mult_209_n1451)
         );
  OAI22_X1 DP_mult_209_U2549 ( .A1(DP_mult_209_n2195), .A2(DP_mult_209_n1747), 
        .B1(DP_mult_209_n1746), .B2(DP_mult_209_n2019), .ZN(DP_mult_209_n1448)
         );
  OAI22_X1 DP_mult_209_U2548 ( .A1(DP_mult_209_n2195), .A2(DP_mult_209_n1753), 
        .B1(DP_mult_209_n1752), .B2(DP_mult_209_n2019), .ZN(DP_mult_209_n1454)
         );
  OAI21_X1 DP_mult_209_U2547 ( .B1(DP_mult_209_n594), .B2(DP_mult_209_n582), 
        .A(DP_mult_209_n583), .ZN(DP_mult_209_n581) );
  XNOR2_X1 DP_mult_209_U2546 ( .A(DP_mult_209_n388), .B(DP_mult_209_n306), 
        .ZN(DP_pipe0_coeff_pipe03[18]) );
  NAND2_X1 DP_mult_209_U2545 ( .A1(DP_mult_209_n1816), .A2(DP_mult_209_n2072), 
        .ZN(DP_mult_209_n277) );
  XNOR2_X1 DP_mult_209_U2544 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2253), .ZN(
        DP_mult_209_n1761) );
  XNOR2_X1 DP_mult_209_U2543 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2253), .ZN(
        DP_mult_209_n1765) );
  XNOR2_X1 DP_mult_209_U2542 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2253), .ZN(
        DP_mult_209_n1769) );
  XNOR2_X1 DP_mult_209_U2541 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2252), .ZN(
        DP_mult_209_n1759) );
  XNOR2_X1 DP_mult_209_U2540 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2252), .ZN(
        DP_mult_209_n1767) );
  XNOR2_X1 DP_mult_209_U2539 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2252), .ZN(
        DP_mult_209_n1763) );
  OAI22_X1 DP_mult_209_U2538 ( .A1(DP_mult_209_n2194), .A2(DP_mult_209_n1743), 
        .B1(DP_mult_209_n1742), .B2(DP_mult_209_n2019), .ZN(DP_mult_209_n1444)
         );
  OAI22_X1 DP_mult_209_U2537 ( .A1(DP_mult_209_n2222), .A2(DP_mult_209_n1737), 
        .B1(DP_mult_209_n1736), .B2(DP_mult_209_n2019), .ZN(DP_mult_209_n1438)
         );
  OAI22_X1 DP_mult_209_U2536 ( .A1(DP_mult_209_n2195), .A2(DP_mult_209_n1735), 
        .B1(DP_mult_209_n1734), .B2(DP_mult_209_n2248), .ZN(DP_mult_209_n1436)
         );
  OAI22_X1 DP_mult_209_U2535 ( .A1(DP_mult_209_n2196), .A2(DP_mult_209_n1739), 
        .B1(DP_mult_209_n1738), .B2(DP_mult_209_n2248), .ZN(DP_mult_209_n1440)
         );
  INV_X1 DP_mult_209_U2534 ( .A(DP_mult_209_n916), .ZN(DP_mult_209_n917) );
  OAI22_X1 DP_mult_209_U2533 ( .A1(DP_mult_209_n2195), .A2(DP_mult_209_n2259), 
        .B1(DP_mult_209_n1756), .B2(DP_mult_209_n2019), .ZN(DP_mult_209_n1192)
         );
  NAND2_X1 DP_mult_209_U2532 ( .A1(DP_mult_209_n805), .A2(DP_mult_209_n820), 
        .ZN(DP_mult_209_n496) );
  XNOR2_X1 DP_mult_209_U2531 ( .A(DP_mult_209_n379), .B(DP_mult_209_n305), 
        .ZN(DP_pipe0_coeff_pipe03[19]) );
  XNOR2_X1 DP_mult_209_U2530 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1667) );
  XNOR2_X1 DP_mult_209_U2529 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1659) );
  XNOR2_X1 DP_mult_209_U2528 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1665) );
  XNOR2_X1 DP_mult_209_U2527 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1669) );
  XNOR2_X1 DP_mult_209_U2526 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1661) );
  XNOR2_X1 DP_mult_209_U2525 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1663) );
  OAI22_X1 DP_mult_209_U2524 ( .A1(DP_mult_209_n2215), .A2(DP_mult_209_n1643), 
        .B1(DP_mult_209_n1642), .B2(DP_mult_209_n2241), .ZN(DP_mult_209_n1348)
         );
  OAI22_X1 DP_mult_209_U2523 ( .A1(DP_mult_209_n2024), .A2(DP_mult_209_n1641), 
        .B1(DP_mult_209_n1640), .B2(DP_mult_209_n2241), .ZN(DP_mult_209_n1346)
         );
  OAI22_X1 DP_mult_209_U2522 ( .A1(DP_mult_209_n2025), .A2(DP_mult_209_n2278), 
        .B1(DP_mult_209_n1656), .B2(DP_mult_209_n2241), .ZN(DP_mult_209_n1188)
         );
  OAI22_X1 DP_mult_209_U2521 ( .A1(DP_mult_209_n2215), .A2(DP_mult_209_n1642), 
        .B1(DP_mult_209_n2241), .B2(DP_mult_209_n1641), .ZN(DP_mult_209_n1347)
         );
  OAI22_X1 DP_mult_209_U2520 ( .A1(DP_mult_209_n2160), .A2(DP_mult_209_n1633), 
        .B1(DP_mult_209_n1632), .B2(DP_mult_209_n2240), .ZN(DP_mult_209_n772)
         );
  OAI22_X1 DP_mult_209_U2519 ( .A1(DP_mult_209_n2024), .A2(DP_mult_209_n1638), 
        .B1(DP_mult_209_n2240), .B2(DP_mult_209_n1637), .ZN(DP_mult_209_n1343)
         );
  OAI22_X1 DP_mult_209_U2518 ( .A1(DP_mult_209_n2160), .A2(DP_mult_209_n1640), 
        .B1(DP_mult_209_n2240), .B2(DP_mult_209_n1639), .ZN(DP_mult_209_n1345)
         );
  OAI22_X1 DP_mult_209_U2517 ( .A1(DP_mult_209_n2216), .A2(DP_mult_209_n1639), 
        .B1(DP_mult_209_n1638), .B2(DP_mult_209_n2241), .ZN(DP_mult_209_n1344)
         );
  OAI22_X1 DP_mult_209_U2516 ( .A1(DP_mult_209_n2024), .A2(DP_mult_209_n1635), 
        .B1(DP_mult_209_n1634), .B2(DP_mult_209_n2241), .ZN(DP_mult_209_n1340)
         );
  OAI22_X1 DP_mult_209_U2515 ( .A1(DP_mult_209_n2160), .A2(DP_mult_209_n1634), 
        .B1(DP_mult_209_n2241), .B2(DP_mult_209_n1633), .ZN(DP_mult_209_n1339)
         );
  OAI22_X1 DP_mult_209_U2514 ( .A1(DP_mult_209_n2024), .A2(DP_mult_209_n1636), 
        .B1(DP_mult_209_n2241), .B2(DP_mult_209_n1635), .ZN(DP_mult_209_n1341)
         );
  OAI22_X1 DP_mult_209_U2513 ( .A1(DP_mult_209_n2025), .A2(DP_mult_209_n1637), 
        .B1(DP_mult_209_n1636), .B2(DP_mult_209_n2241), .ZN(DP_mult_209_n1342)
         );
  NAND2_X1 DP_mult_209_U2512 ( .A1(DP_mult_209_n1806), .A2(DP_mult_209_n2116), 
        .ZN(DP_mult_209_n297) );
  OAI22_X1 DP_mult_209_U2511 ( .A1(DP_mult_209_n2204), .A2(DP_mult_209_n1504), 
        .B1(DP_mult_209_n2045), .B2(DP_mult_209_n1503), .ZN(DP_mult_209_n1215)
         );
  OAI22_X1 DP_mult_209_U2510 ( .A1(DP_mult_209_n2204), .A2(DP_mult_209_n1498), 
        .B1(DP_mult_209_n2045), .B2(DP_mult_209_n1497), .ZN(DP_mult_209_n1209)
         );
  OAI22_X1 DP_mult_209_U2509 ( .A1(DP_mult_209_n2204), .A2(DP_mult_209_n1505), 
        .B1(DP_mult_209_n1504), .B2(DP_mult_209_n2064), .ZN(DP_mult_209_n1216)
         );
  OAI22_X1 DP_mult_209_U2508 ( .A1(DP_mult_209_n1968), .A2(DP_mult_209_n1499), 
        .B1(DP_mult_209_n1498), .B2(DP_mult_209_n2045), .ZN(DP_mult_209_n1210)
         );
  OAI22_X1 DP_mult_209_U2507 ( .A1(DP_mult_209_n2204), .A2(DP_mult_209_n2305), 
        .B1(DP_mult_209_n1506), .B2(DP_mult_209_n2045), .ZN(DP_mult_209_n1182)
         );
  OAI22_X1 DP_mult_209_U2506 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1493), 
        .B1(DP_mult_209_n1492), .B2(DP_mult_209_n2064), .ZN(DP_mult_209_n1204)
         );
  OAI22_X1 DP_mult_209_U2505 ( .A1(DP_mult_209_n1968), .A2(DP_mult_209_n1503), 
        .B1(DP_mult_209_n1502), .B2(DP_mult_209_n2064), .ZN(DP_mult_209_n1214)
         );
  OAI22_X1 DP_mult_209_U2504 ( .A1(DP_mult_209_n1968), .A2(DP_mult_209_n1500), 
        .B1(DP_mult_209_n2045), .B2(DP_mult_209_n1499), .ZN(DP_mult_209_n1211)
         );
  OAI22_X1 DP_mult_209_U2503 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1501), 
        .B1(DP_mult_209_n1500), .B2(DP_mult_209_n2045), .ZN(DP_mult_209_n1212)
         );
  OAI22_X1 DP_mult_209_U2502 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1502), 
        .B1(DP_mult_209_n2045), .B2(DP_mult_209_n1501), .ZN(DP_mult_209_n1213)
         );
  OAI22_X1 DP_mult_209_U2501 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1489), 
        .B1(DP_mult_209_n1488), .B2(DP_mult_209_n2064), .ZN(DP_mult_209_n1200)
         );
  OAI22_X1 DP_mult_209_U2500 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1494), 
        .B1(DP_mult_209_n2064), .B2(DP_mult_209_n1493), .ZN(DP_mult_209_n1205)
         );
  OAI22_X1 DP_mult_209_U2499 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1495), 
        .B1(DP_mult_209_n1494), .B2(DP_mult_209_n2064), .ZN(DP_mult_209_n1206)
         );
  OAI22_X1 DP_mult_209_U2498 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1496), 
        .B1(DP_mult_209_n2064), .B2(DP_mult_209_n1495), .ZN(DP_mult_209_n1207)
         );
  OAI22_X1 DP_mult_209_U2497 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1497), 
        .B1(DP_mult_209_n1496), .B2(DP_mult_209_n2045), .ZN(DP_mult_209_n1208)
         );
  OAI22_X1 DP_mult_209_U2496 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1487), 
        .B1(DP_mult_209_n1486), .B2(DP_mult_209_n2064), .ZN(DP_mult_209_n1198)
         );
  OAI22_X1 DP_mult_209_U2495 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1491), 
        .B1(DP_mult_209_n1490), .B2(DP_mult_209_n2064), .ZN(DP_mult_209_n1202)
         );
  OAI22_X1 DP_mult_209_U2494 ( .A1(DP_mult_209_n1938), .A2(DP_mult_209_n1485), 
        .B1(DP_mult_209_n1484), .B2(DP_mult_209_n2045), .ZN(DP_mult_209_n1196)
         );
  OAI22_X1 DP_mult_209_U2493 ( .A1(DP_mult_209_n1938), .A2(DP_mult_209_n1483), 
        .B1(DP_mult_209_n1482), .B2(DP_mult_209_n2064), .ZN(DP_mult_209_n676)
         );
  XNOR2_X1 DP_mult_209_U2492 ( .A(DP_mult_209_n370), .B(DP_mult_209_n304), 
        .ZN(DP_pipe0_coeff_pipe03[20]) );
  OAI21_X1 DP_mult_209_U2491 ( .B1(DP_mult_209_n542), .B2(DP_mult_209_n550), 
        .A(DP_mult_209_n543), .ZN(DP_mult_209_n541) );
  INV_X1 DP_mult_209_U2490 ( .A(DP_mult_209_n2145), .ZN(DP_mult_209_n673) );
  XNOR2_X1 DP_mult_209_U2489 ( .A(DP_mult_209_n353), .B(DP_mult_209_n303), 
        .ZN(DP_pipe0_coeff_pipe03[21]) );
  OAI22_X1 DP_mult_209_U2488 ( .A1(DP_mult_209_n2158), .A2(DP_mult_209_n1703), 
        .B1(DP_mult_209_n1702), .B2(DP_mult_209_n2245), .ZN(DP_mult_209_n1406)
         );
  OAI22_X1 DP_mult_209_U2487 ( .A1(DP_mult_209_n2157), .A2(DP_mult_209_n1705), 
        .B1(DP_mult_209_n1704), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1408)
         );
  NAND2_X1 DP_mult_209_U2486 ( .A1(DP_mult_209_n761), .A2(DP_mult_209_n774), 
        .ZN(DP_mult_209_n461) );
  OAI22_X1 DP_mult_209_U2485 ( .A1(DP_mult_209_n2214), .A2(DP_mult_209_n1628), 
        .B1(DP_mult_209_n1627), .B2(DP_mult_209_n2237), .ZN(DP_mult_209_n1334)
         );
  OAI22_X1 DP_mult_209_U2484 ( .A1(DP_mult_209_n1992), .A2(DP_mult_209_n1630), 
        .B1(DP_mult_209_n1629), .B2(DP_mult_209_n2238), .ZN(DP_mult_209_n1336)
         );
  NAND2_X1 DP_mult_209_U2483 ( .A1(DP_mult_209_n709), .A2(DP_mult_209_n716), 
        .ZN(DP_mult_209_n409) );
  OAI22_X1 DP_mult_209_U2482 ( .A1(DP_mult_209_n2209), .A2(DP_mult_209_n1576), 
        .B1(DP_mult_209_n1575), .B2(DP_mult_209_n2231), .ZN(DP_mult_209_n1284)
         );
  OAI22_X1 DP_mult_209_U2481 ( .A1(DP_mult_209_n2209), .A2(DP_mult_209_n1574), 
        .B1(DP_mult_209_n1573), .B2(DP_mult_209_n2231), .ZN(DP_mult_209_n1282)
         );
  OAI22_X1 DP_mult_209_U2480 ( .A1(DP_mult_209_n2209), .A2(DP_mult_209_n1572), 
        .B1(DP_mult_209_n1571), .B2(DP_mult_209_n2231), .ZN(DP_mult_209_n1280)
         );
  OAI22_X1 DP_mult_209_U2479 ( .A1(DP_mult_209_n2209), .A2(DP_mult_209_n1577), 
        .B1(DP_mult_209_n2231), .B2(DP_mult_209_n1576), .ZN(DP_mult_209_n1285)
         );
  OAI22_X1 DP_mult_209_U2478 ( .A1(DP_mult_209_n1962), .A2(DP_mult_209_n1573), 
        .B1(DP_mult_209_n2230), .B2(DP_mult_209_n1572), .ZN(DP_mult_209_n1281)
         );
  OAI22_X1 DP_mult_209_U2477 ( .A1(DP_mult_209_n2209), .A2(DP_mult_209_n1578), 
        .B1(DP_mult_209_n1577), .B2(DP_mult_209_n2231), .ZN(DP_mult_209_n1286)
         );
  OAI22_X1 DP_mult_209_U2476 ( .A1(DP_mult_209_n2209), .A2(DP_mult_209_n1569), 
        .B1(DP_mult_209_n2231), .B2(DP_mult_209_n1568), .ZN(DP_mult_209_n1277)
         );
  OAI22_X1 DP_mult_209_U2475 ( .A1(DP_mult_209_n2209), .A2(DP_mult_209_n1579), 
        .B1(DP_mult_209_n2231), .B2(DP_mult_209_n1578), .ZN(DP_mult_209_n1287)
         );
  OAI22_X1 DP_mult_209_U2474 ( .A1(DP_mult_209_n1963), .A2(DP_mult_209_n1580), 
        .B1(DP_mult_209_n1579), .B2(DP_mult_209_n2230), .ZN(DP_mult_209_n1288)
         );
  OAI22_X1 DP_mult_209_U2473 ( .A1(DP_mult_209_n1962), .A2(DP_mult_209_n1571), 
        .B1(DP_mult_209_n2230), .B2(DP_mult_209_n1570), .ZN(DP_mult_209_n1279)
         );
  OAI22_X1 DP_mult_209_U2472 ( .A1(DP_mult_209_n1962), .A2(DP_mult_209_n1575), 
        .B1(DP_mult_209_n2230), .B2(DP_mult_209_n1574), .ZN(DP_mult_209_n1283)
         );
  OAI22_X1 DP_mult_209_U2471 ( .A1(DP_mult_209_n1963), .A2(DP_mult_209_n1570), 
        .B1(DP_mult_209_n1569), .B2(DP_mult_209_n2230), .ZN(DP_mult_209_n1278)
         );
  XNOR2_X1 DP_mult_209_U2470 ( .A(DP_mult_209_n342), .B(DP_mult_209_n302), 
        .ZN(DP_pipe0_coeff_pipe03[22]) );
  OAI22_X1 DP_mult_209_U2469 ( .A1(DP_mult_209_n2208), .A2(DP_mult_209_n1538), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1537), .ZN(DP_mult_209_n1247)
         );
  OAI22_X1 DP_mult_209_U2468 ( .A1(DP_mult_209_n2207), .A2(DP_mult_209_n1533), 
        .B1(DP_mult_209_n1532), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n692)
         );
  OAI22_X1 DP_mult_209_U2467 ( .A1(DP_mult_209_n2097), .A2(DP_mult_209_n1539), 
        .B1(DP_mult_209_n1538), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1248)
         );
  OAI22_X1 DP_mult_209_U2466 ( .A1(DP_mult_209_n2207), .A2(DP_mult_209_n1540), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1539), .ZN(DP_mult_209_n1249)
         );
  OAI22_X1 DP_mult_209_U2465 ( .A1(DP_mult_209_n2097), .A2(DP_mult_209_n2297), 
        .B1(DP_mult_209_n1556), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1184)
         );
  OAI22_X1 DP_mult_209_U2464 ( .A1(DP_mult_209_n2208), .A2(DP_mult_209_n1541), 
        .B1(DP_mult_209_n1540), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1250)
         );
  OAI22_X1 DP_mult_209_U2463 ( .A1(DP_mult_209_n2207), .A2(DP_mult_209_n1542), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1541), .ZN(DP_mult_209_n1251)
         );
  OAI22_X1 DP_mult_209_U2462 ( .A1(DP_mult_209_n2208), .A2(DP_mult_209_n1543), 
        .B1(DP_mult_209_n1542), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1252)
         );
  INV_X1 DP_mult_209_U2461 ( .A(DP_mult_209_n692), .ZN(DP_mult_209_n693) );
  OAI22_X1 DP_mult_209_U2460 ( .A1(DP_mult_209_n2097), .A2(DP_mult_209_n1537), 
        .B1(DP_mult_209_n1536), .B2(DP_mult_209_n2229), .ZN(DP_mult_209_n1246)
         );
  OAI22_X1 DP_mult_209_U2459 ( .A1(DP_mult_209_n2208), .A2(DP_mult_209_n1534), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1533), .ZN(DP_mult_209_n1243)
         );
  OAI22_X1 DP_mult_209_U2458 ( .A1(DP_mult_209_n2207), .A2(DP_mult_209_n1535), 
        .B1(DP_mult_209_n1534), .B2(DP_mult_209_n2063), .ZN(DP_mult_209_n1244)
         );
  OAI22_X1 DP_mult_209_U2457 ( .A1(DP_mult_209_n2207), .A2(DP_mult_209_n1536), 
        .B1(DP_mult_209_n2229), .B2(DP_mult_209_n1535), .ZN(DP_mult_209_n1245)
         );
  OAI21_X1 DP_mult_209_U2456 ( .B1(DP_mult_209_n364), .B2(DP_mult_209_n387), 
        .A(DP_mult_209_n365), .ZN(DP_mult_209_n363) );
  NAND2_X1 DP_mult_209_U2455 ( .A1(DP_mult_209_n345), .A2(DP_mult_209_n2181), 
        .ZN(DP_mult_209_n336) );
  INV_X1 DP_mult_209_U2454 ( .A(DP_mult_209_n345), .ZN(DP_mult_209_n343) );
  OAI22_X1 DP_mult_209_U2453 ( .A1(DP_mult_209_n1954), .A2(DP_mult_209_n1516), 
        .B1(DP_mult_209_n1515), .B2(DP_mult_209_n2227), .ZN(DP_mult_209_n1226)
         );
  OAI22_X1 DP_mult_209_U2452 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n2301), 
        .B1(DP_mult_209_n1531), .B2(DP_mult_209_n2228), .ZN(DP_mult_209_n1183)
         );
  OR2_X1 DP_mult_209_U2451 ( .A1(DP_mult_209_n1215), .A2(DP_mult_209_n1237), 
        .ZN(DP_mult_209_n938) );
  OAI22_X1 DP_mult_209_U2450 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1512), 
        .B1(DP_mult_209_n1511), .B2(DP_mult_209_n2227), .ZN(DP_mult_209_n1222)
         );
  XNOR2_X1 DP_mult_209_U2449 ( .A(DP_mult_209_n1945), .B(DP_mult_209_n1215), 
        .ZN(DP_mult_209_n939) );
  OAI22_X1 DP_mult_209_U2448 ( .A1(DP_mult_209_n1954), .A2(DP_mult_209_n1514), 
        .B1(DP_mult_209_n1513), .B2(DP_mult_209_n2228), .ZN(DP_mult_209_n1224)
         );
  OAI22_X1 DP_mult_209_U2447 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1510), 
        .B1(DP_mult_209_n1509), .B2(DP_mult_209_n2227), .ZN(DP_mult_209_n1220)
         );
  OAI22_X1 DP_mult_209_U2446 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1518), 
        .B1(DP_mult_209_n1517), .B2(DP_mult_209_n2227), .ZN(DP_mult_209_n1228)
         );
  OAI22_X1 DP_mult_209_U2445 ( .A1(DP_mult_209_n2206), .A2(DP_mult_209_n1508), 
        .B1(DP_mult_209_n1507), .B2(DP_mult_209_n2227), .ZN(DP_mult_209_n682)
         );
  INV_X1 DP_mult_209_U2444 ( .A(DP_mult_209_n2202), .ZN(DP_mult_209_n508) );
  AOI21_X1 DP_mult_209_U2443 ( .B1(DP_mult_209_n508), .B2(DP_mult_209_n2118), 
        .A(DP_mult_209_n2108), .ZN(DP_mult_209_n488) );
  AOI21_X1 DP_mult_209_U2442 ( .B1(DP_mult_209_n508), .B2(DP_mult_209_n478), 
        .A(DP_mult_209_n479), .ZN(DP_mult_209_n477) );
  AOI21_X1 DP_mult_209_U2441 ( .B1(DP_mult_209_n508), .B2(DP_mult_209_n465), 
        .A(DP_mult_209_n466), .ZN(DP_mult_209_n464) );
  AOI21_X1 DP_mult_209_U2440 ( .B1(DP_mult_209_n508), .B2(DP_mult_209_n668), 
        .A(DP_mult_209_n501), .ZN(DP_mult_209_n499) );
  OAI22_X1 DP_mult_209_U2439 ( .A1(DP_mult_209_n2211), .A2(DP_mult_209_n2288), 
        .B1(DP_mult_209_n1606), .B2(DP_mult_209_n2234), .ZN(DP_mult_209_n1186)
         );
  OAI22_X1 DP_mult_209_U2438 ( .A1(DP_mult_209_n2211), .A2(DP_mult_209_n1586), 
        .B1(DP_mult_209_n2235), .B2(DP_mult_209_n1585), .ZN(DP_mult_209_n1293)
         );
  OAI22_X1 DP_mult_209_U2437 ( .A1(DP_mult_209_n2155), .A2(DP_mult_209_n1585), 
        .B1(DP_mult_209_n1584), .B2(DP_mult_209_n2234), .ZN(DP_mult_209_n1292)
         );
  OAI22_X1 DP_mult_209_U2436 ( .A1(DP_mult_209_n2212), .A2(DP_mult_209_n1591), 
        .B1(DP_mult_209_n1590), .B2(DP_mult_209_n2234), .ZN(DP_mult_209_n1298)
         );
  OAI22_X1 DP_mult_209_U2435 ( .A1(DP_mult_209_n2155), .A2(DP_mult_209_n1587), 
        .B1(DP_mult_209_n1586), .B2(DP_mult_209_n2234), .ZN(DP_mult_209_n1294)
         );
  OAI22_X1 DP_mult_209_U2434 ( .A1(DP_mult_209_n2212), .A2(DP_mult_209_n1583), 
        .B1(DP_mult_209_n1582), .B2(DP_mult_209_n2235), .ZN(DP_mult_209_n724)
         );
  OAI22_X1 DP_mult_209_U2433 ( .A1(DP_mult_209_n2156), .A2(DP_mult_209_n1592), 
        .B1(DP_mult_209_n2235), .B2(DP_mult_209_n1591), .ZN(DP_mult_209_n1299)
         );
  OAI22_X1 DP_mult_209_U2432 ( .A1(DP_mult_209_n2156), .A2(DP_mult_209_n1588), 
        .B1(DP_mult_209_n2235), .B2(DP_mult_209_n1587), .ZN(DP_mult_209_n1295)
         );
  OAI22_X1 DP_mult_209_U2431 ( .A1(DP_mult_209_n2156), .A2(DP_mult_209_n1589), 
        .B1(DP_mult_209_n1588), .B2(DP_mult_209_n2235), .ZN(DP_mult_209_n1296)
         );
  OAI22_X1 DP_mult_209_U2430 ( .A1(DP_mult_209_n2156), .A2(DP_mult_209_n1584), 
        .B1(DP_mult_209_n2235), .B2(DP_mult_209_n1583), .ZN(DP_mult_209_n1291)
         );
  OAI22_X1 DP_mult_209_U2429 ( .A1(DP_mult_209_n2211), .A2(DP_mult_209_n1590), 
        .B1(DP_mult_209_n2234), .B2(DP_mult_209_n1589), .ZN(DP_mult_209_n1297)
         );
  OAI22_X1 DP_mult_209_U2428 ( .A1(DP_mult_209_n2211), .A2(DP_mult_209_n1593), 
        .B1(DP_mult_209_n1592), .B2(DP_mult_209_n2235), .ZN(DP_mult_209_n1300)
         );
  OAI21_X1 DP_mult_209_U2427 ( .B1(DP_mult_209_n421), .B2(DP_mult_209_n347), 
        .A(DP_mult_209_n348), .ZN(DP_mult_209_n346) );
  INV_X1 DP_mult_209_U2426 ( .A(DP_mult_209_n421), .ZN(DP_mult_209_n423) );
  OAI21_X1 DP_mult_209_U2425 ( .B1(DP_mult_209_n390), .B2(DP_mult_209_n384), 
        .A(DP_mult_209_n387), .ZN(DP_mult_209_n383) );
  NAND2_X1 DP_mult_209_U2424 ( .A1(DP_mult_209_n525), .A2(DP_mult_209_n511), 
        .ZN(DP_mult_209_n505) );
  NAND2_X1 DP_mult_209_U2423 ( .A1(DP_mult_209_n478), .A2(DP_mult_209_n2004), 
        .ZN(DP_mult_209_n476) );
  OAI21_X1 DP_mult_209_U2422 ( .B1(DP_mult_209_n566), .B2(DP_mult_209_n538), 
        .A(DP_mult_209_n539), .ZN(DP_mult_209_n537) );
  NAND2_X1 DP_mult_209_U2421 ( .A1(DP_mult_209_n983), .A2(DP_mult_209_n1002), 
        .ZN(DP_mult_209_n564) );
  INV_X1 DP_mult_209_U2420 ( .A(DP_mult_209_n2068), .ZN(DP_mult_209_n671) );
  OAI22_X1 DP_mult_209_U2419 ( .A1(DP_mult_209_n2192), .A2(DP_mult_209_n1674), 
        .B1(DP_mult_209_n1673), .B2(DP_mult_209_n2243), .ZN(DP_mult_209_n1378)
         );
  OAI22_X1 DP_mult_209_U2418 ( .A1(DP_mult_209_n2217), .A2(DP_mult_209_n1678), 
        .B1(DP_mult_209_n1677), .B2(DP_mult_209_n2242), .ZN(DP_mult_209_n1382)
         );
  OAI22_X1 DP_mult_209_U2417 ( .A1(DP_mult_209_n2217), .A2(DP_mult_209_n1680), 
        .B1(DP_mult_209_n1679), .B2(DP_mult_209_n2243), .ZN(DP_mult_209_n1384)
         );
  OAI22_X1 DP_mult_209_U2416 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1669), 
        .B1(DP_mult_209_n2242), .B2(DP_mult_209_n1668), .ZN(DP_mult_209_n1373)
         );
  OAI22_X1 DP_mult_209_U2415 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1670), 
        .B1(DP_mult_209_n1669), .B2(DP_mult_209_n2242), .ZN(DP_mult_209_n1374)
         );
  OAI22_X1 DP_mult_209_U2414 ( .A1(DP_mult_209_n2217), .A2(DP_mult_209_n1676), 
        .B1(DP_mult_209_n1675), .B2(DP_mult_209_n2242), .ZN(DP_mult_209_n1380)
         );
  OAI22_X1 DP_mult_209_U2413 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1673), 
        .B1(DP_mult_209_n2243), .B2(DP_mult_209_n1672), .ZN(DP_mult_209_n1377)
         );
  OAI22_X1 DP_mult_209_U2412 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1671), 
        .B1(DP_mult_209_n2242), .B2(DP_mult_209_n1670), .ZN(DP_mult_209_n1375)
         );
  OAI22_X1 DP_mult_209_U2411 ( .A1(DP_mult_209_n2192), .A2(DP_mult_209_n1672), 
        .B1(DP_mult_209_n1671), .B2(DP_mult_209_n2243), .ZN(DP_mult_209_n1376)
         );
  OAI22_X1 DP_mult_209_U2410 ( .A1(DP_mult_209_n2192), .A2(DP_mult_209_n1677), 
        .B1(DP_mult_209_n2243), .B2(DP_mult_209_n1676), .ZN(DP_mult_209_n1381)
         );
  OAI22_X1 DP_mult_209_U2409 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1675), 
        .B1(DP_mult_209_n2243), .B2(DP_mult_209_n1674), .ZN(DP_mult_209_n1379)
         );
  OAI22_X1 DP_mult_209_U2408 ( .A1(DP_mult_209_n2191), .A2(DP_mult_209_n1679), 
        .B1(DP_mult_209_n2242), .B2(DP_mult_209_n1678), .ZN(DP_mult_209_n1383)
         );
  NAND2_X1 DP_mult_209_U2407 ( .A1(DP_mult_209_n941), .A2(DP_mult_209_n962), 
        .ZN(DP_mult_209_n550) );
  NAND2_X1 DP_mult_209_U2406 ( .A1(DP_mult_209_n2005), .A2(DP_mult_209_n474), 
        .ZN(DP_mult_209_n314) );
  NAND2_X1 DP_mult_209_U2405 ( .A1(DP_mult_209_n839), .A2(DP_mult_209_n856), 
        .ZN(DP_mult_209_n514) );
  OAI21_X1 DP_mult_209_U2404 ( .B1(DP_mult_209_n2059), .B2(DP_mult_209_n521), 
        .A(DP_mult_209_n514), .ZN(DP_mult_209_n512) );
  NAND2_X1 DP_mult_209_U2403 ( .A1(DP_mult_209_n749), .A2(DP_mult_209_n760), 
        .ZN(DP_mult_209_n439) );
  NOR2_X1 DP_mult_209_U2402 ( .A1(DP_mult_209_n749), .A2(DP_mult_209_n760), 
        .ZN(DP_mult_209_n438) );
  INV_X1 DP_mult_209_U2401 ( .A(DP_mult_209_n772), .ZN(DP_mult_209_n773) );
  INV_X1 DP_mult_209_U2400 ( .A(DP_mult_209_n706), .ZN(DP_mult_209_n707) );
  OAI21_X1 DP_mult_209_U2399 ( .B1(DP_mult_209_n2066), .B2(DP_mult_209_n2232), 
        .A(DP_mult_209_n2314), .ZN(DP_mult_209_n1266) );
  NAND2_X1 DP_mult_209_U2398 ( .A1(DP_mult_209_n701), .A2(DP_mult_209_n708), 
        .ZN(DP_mult_209_n396) );
  NOR2_X1 DP_mult_209_U2397 ( .A1(DP_mult_209_n336), .A2(DP_mult_209_n334), 
        .ZN(DP_mult_209_n332) );
  AOI21_X1 DP_mult_209_U2396 ( .B1(DP_mult_209_n2047), .B2(DP_mult_209_n2137), 
        .A(DP_mult_209_n519), .ZN(DP_mult_209_n517) );
  INV_X1 DP_mult_209_U2395 ( .A(DP_mult_209_n2131), .ZN(DP_mult_209_n524) );
  OAI21_X1 DP_mult_209_U2394 ( .B1(DP_mult_209_n1975), .B2(DP_mult_209_n2187), 
        .A(DP_mult_209_n2309), .ZN(DP_mult_209_n1386) );
  NAND2_X1 DP_mult_209_U2393 ( .A1(DP_mult_209_n2005), .A2(DP_mult_209_n666), 
        .ZN(DP_mult_209_n467) );
  AOI21_X1 DP_mult_209_U2392 ( .B1(DP_mult_209_n2166), .B2(DP_mult_209_n483), 
        .A(DP_mult_209_n1956), .ZN(DP_mult_209_n468) );
  NAND2_X1 DP_mult_209_U2391 ( .A1(DP_mult_209_n727), .A2(DP_mult_209_n736), 
        .ZN(DP_mult_209_n429) );
  NOR2_X1 DP_mult_209_U2390 ( .A1(DP_mult_209_n897), .A2(DP_mult_209_n918), 
        .ZN(DP_mult_209_n534) );
  NAND2_X1 DP_mult_209_U2389 ( .A1(DP_mult_209_n2114), .A2(DP_mult_209_n2137), 
        .ZN(DP_mult_209_n516) );
  XNOR2_X1 DP_mult_209_U2388 ( .A(DP_mult_209_n462), .B(DP_mult_209_n313), 
        .ZN(DP_pipe0_coeff_pipe03[11]) );
  OAI21_X1 DP_mult_209_U2387 ( .B1(DP_mult_209_n2078), .B2(DP_mult_209_n2012), 
        .A(DP_mult_209_n2311), .ZN(DP_mult_209_n1338) );
  NOR2_X1 DP_mult_209_U2386 ( .A1(DP_mult_209_n737), .A2(DP_mult_209_n748), 
        .ZN(DP_mult_209_n435) );
  OAI21_X1 DP_mult_209_U2385 ( .B1(DP_mult_209_n503), .B2(DP_mult_209_n2154), 
        .A(DP_mult_209_n496), .ZN(DP_mult_209_n490) );
  INV_X1 DP_mult_209_U2384 ( .A(DP_mult_209_n2154), .ZN(DP_mult_209_n667) );
  NAND2_X1 DP_mult_209_U2383 ( .A1(DP_mult_209_n540), .A2(DP_mult_209_n552), 
        .ZN(DP_mult_209_n538) );
  AOI21_X1 DP_mult_209_U2382 ( .B1(DP_mult_209_n540), .B2(DP_mult_209_n553), 
        .A(DP_mult_209_n541), .ZN(DP_mult_209_n539) );
  NAND2_X1 DP_mult_209_U2381 ( .A1(DP_mult_209_n877), .A2(DP_mult_209_n896), 
        .ZN(DP_mult_209_n532) );
  OAI22_X1 DP_mult_209_U2380 ( .A1(DP_mult_209_n2194), .A2(DP_mult_209_n1742), 
        .B1(DP_mult_209_n2019), .B2(DP_mult_209_n1741), .ZN(DP_mult_209_n1443)
         );
  OAI22_X1 DP_mult_209_U2379 ( .A1(DP_mult_209_n2195), .A2(DP_mult_209_n1734), 
        .B1(DP_mult_209_n2248), .B2(DP_mult_209_n1733), .ZN(DP_mult_209_n1435)
         );
  OAI22_X1 DP_mult_209_U2378 ( .A1(DP_mult_209_n2196), .A2(DP_mult_209_n1740), 
        .B1(DP_mult_209_n2248), .B2(DP_mult_209_n1739), .ZN(DP_mult_209_n1441)
         );
  OAI22_X1 DP_mult_209_U2377 ( .A1(DP_mult_209_n2196), .A2(DP_mult_209_n1736), 
        .B1(DP_mult_209_n2019), .B2(DP_mult_209_n1735), .ZN(DP_mult_209_n1437)
         );
  OAI22_X1 DP_mult_209_U2376 ( .A1(DP_mult_209_n2196), .A2(DP_mult_209_n1738), 
        .B1(DP_mult_209_n2248), .B2(DP_mult_209_n1737), .ZN(DP_mult_209_n1439)
         );
  NOR2_X1 DP_mult_209_U2375 ( .A1(DP_mult_209_n456), .A2(DP_mult_209_n480), 
        .ZN(DP_mult_209_n454) );
  INV_X1 DP_mult_209_U2374 ( .A(DP_mult_209_n480), .ZN(DP_mult_209_n666) );
  OAI21_X1 DP_mult_209_U2373 ( .B1(DP_mult_209_n492), .B2(DP_mult_209_n480), 
        .A(DP_mult_209_n481), .ZN(DP_mult_209_n479) );
  NOR2_X1 DP_mult_209_U2372 ( .A1(DP_mult_209_n2119), .A2(DP_mult_209_n480), 
        .ZN(DP_mult_209_n478) );
  AOI21_X1 DP_mult_209_U2371 ( .B1(DP_mult_209_n2169), .B2(DP_mult_209_n2165), 
        .A(DP_mult_209_n1981), .ZN(DP_mult_209_n572) );
  NAND2_X1 DP_mult_209_U2370 ( .A1(DP_mult_209_n2169), .A2(DP_mult_209_n2170), 
        .ZN(DP_mult_209_n571) );
  XNOR2_X1 DP_mult_209_U2369 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2251), .ZN(
        DP_mult_209_n1757) );
  XNOR2_X1 DP_mult_209_U2368 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2251), .ZN(
        DP_mult_209_n1775) );
  XNOR2_X1 DP_mult_209_U2367 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2251), .ZN(
        DP_mult_209_n1777) );
  XNOR2_X1 DP_mult_209_U2366 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2251), .ZN(
        DP_mult_209_n1773) );
  XOR2_X1 DP_mult_209_U2365 ( .A(DP_coeffs_ff_int[95]), .B(
        DP_coeffs_ff_int[94]), .Z(DP_mult_209_n1817) );
  NOR2_X1 DP_mult_209_U2364 ( .A1(DP_mult_209_n531), .A2(DP_mult_209_n534), 
        .ZN(DP_mult_209_n525) );
  OAI22_X1 DP_mult_209_U2363 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n2254), 
        .B1(DP_mult_209_n1781), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1193)
         );
  NOR2_X1 DP_mult_209_U2362 ( .A1(DP_mult_209_n789), .A2(DP_mult_209_n804), 
        .ZN(DP_mult_209_n480) );
  AOI21_X1 DP_mult_209_U2361 ( .B1(DP_mult_209_n359), .B2(DP_mult_209_n2180), 
        .A(DP_mult_209_n350), .ZN(DP_mult_209_n348) );
  NAND2_X1 DP_mult_209_U2360 ( .A1(DP_mult_209_n356), .A2(DP_mult_209_n2180), 
        .ZN(DP_mult_209_n347) );
  XNOR2_X1 DP_mult_209_U2359 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2300), .ZN(
        DP_mult_209_n1515) );
  XNOR2_X1 DP_mult_209_U2358 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2300), .ZN(
        DP_mult_209_n1511) );
  XNOR2_X1 DP_mult_209_U2357 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2300), .ZN(
        DP_mult_209_n1517) );
  XNOR2_X1 DP_mult_209_U2356 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2299), .ZN(
        DP_mult_209_n1519) );
  XNOR2_X1 DP_mult_209_U2355 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2299), .ZN(
        DP_mult_209_n1509) );
  XNOR2_X1 DP_mult_209_U2354 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2300), .ZN(
        DP_mult_209_n1513) );
  OAI21_X1 DP_mult_209_U2353 ( .B1(DP_mult_209_n590), .B2(DP_mult_209_n593), 
        .A(DP_mult_209_n591), .ZN(DP_mult_209_n589) );
  NOR2_X1 DP_mult_209_U2352 ( .A1(DP_mult_209_n590), .A2(DP_mult_209_n592), 
        .ZN(DP_mult_209_n588) );
  OAI21_X1 DP_mult_209_U2351 ( .B1(DP_mult_209_n428), .B2(DP_mult_209_n436), 
        .A(DP_mult_209_n429), .ZN(DP_mult_209_n427) );
  INV_X1 DP_mult_209_U2350 ( .A(DP_mult_209_n428), .ZN(DP_mult_209_n661) );
  AOI21_X1 DP_mult_209_U2349 ( .B1(DP_mult_209_n2167), .B2(DP_mult_209_n1956), 
        .A(DP_mult_209_n459), .ZN(DP_mult_209_n457) );
  INV_X1 DP_mult_209_U2348 ( .A(DP_mult_209_n283), .ZN(DP_mult_209_n2218) );
  INV_X1 DP_mult_209_U2347 ( .A(DP_mult_209_n382), .ZN(DP_mult_209_n380) );
  AOI21_X1 DP_mult_209_U2346 ( .B1(DP_mult_209_n526), .B2(DP_mult_209_n2057), 
        .A(DP_mult_209_n512), .ZN(DP_mult_209_n506) );
  NOR2_X1 DP_mult_209_U2345 ( .A1(DP_mult_209_n727), .A2(DP_mult_209_n736), 
        .ZN(DP_mult_209_n428) );
  AOI21_X1 DP_mult_209_U2344 ( .B1(DP_mult_209_n581), .B2(DP_mult_209_n567), 
        .A(DP_mult_209_n568), .ZN(DP_mult_209_n566) );
  NAND2_X1 DP_mult_209_U2343 ( .A1(DP_mult_209_n1165), .A2(DP_mult_209_n1170), 
        .ZN(DP_mult_209_n632) );
  OAI21_X1 DP_mult_209_U2342 ( .B1(DP_mult_209_n337), .B2(DP_mult_209_n334), 
        .A(DP_mult_209_n335), .ZN(DP_mult_209_n333) );
  AOI21_X1 DP_mult_209_U2341 ( .B1(DP_mult_209_n423), .B2(DP_mult_209_n2172), 
        .A(DP_mult_209_n416), .ZN(DP_mult_209_n412) );
  NAND2_X1 DP_mult_209_U2340 ( .A1(DP_mult_209_n422), .A2(DP_mult_209_n2172), 
        .ZN(DP_mult_209_n411) );
  AOI21_X1 DP_mult_209_U2339 ( .B1(DP_mult_209_n333), .B2(DP_mult_209_n2182), 
        .A(DP_mult_209_n2178), .ZN(DP_mult_209_n327) );
  NAND2_X1 DP_mult_209_U2338 ( .A1(DP_mult_209_n2172), .A2(DP_mult_209_n418), 
        .ZN(DP_mult_209_n309) );
  OAI21_X1 DP_mult_209_U2337 ( .B1(DP_mult_209_n2223), .B2(DP_mult_209_n2188), 
        .A(DP_mult_209_n2307), .ZN(DP_mult_209_n1434) );
  NAND2_X1 DP_mult_209_U2336 ( .A1(DP_mult_209_n2004), .A2(DP_mult_209_n2118), 
        .ZN(DP_mult_209_n487) );
  NOR2_X1 DP_mult_209_U2335 ( .A1(DP_mult_209_n857), .A2(DP_mult_209_n876), 
        .ZN(DP_mult_209_n520) );
  NAND2_X1 DP_mult_209_U2334 ( .A1(DP_mult_209_n857), .A2(DP_mult_209_n876), 
        .ZN(DP_mult_209_n521) );
  NAND2_X1 DP_mult_209_U2333 ( .A1(DP_mult_209_n1171), .A2(DP_mult_209_n1174), 
        .ZN(DP_mult_209_n634) );
  OAI22_X1 DP_mult_209_U2332 ( .A1(DP_mult_209_n2219), .A2(DP_mult_209_n1699), 
        .B1(DP_mult_209_n1698), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1402)
         );
  OAI22_X1 DP_mult_209_U2331 ( .A1(DP_mult_209_n2023), .A2(DP_mult_209_n1700), 
        .B1(DP_mult_209_n2245), .B2(DP_mult_209_n1699), .ZN(DP_mult_209_n1403)
         );
  OAI22_X1 DP_mult_209_U2330 ( .A1(DP_mult_209_n2158), .A2(DP_mult_209_n1697), 
        .B1(DP_mult_209_n1696), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1400)
         );
  OAI22_X1 DP_mult_209_U2329 ( .A1(DP_mult_209_n2157), .A2(DP_mult_209_n1702), 
        .B1(DP_mult_209_n2245), .B2(DP_mult_209_n1701), .ZN(DP_mult_209_n1405)
         );
  OAI22_X1 DP_mult_209_U2328 ( .A1(DP_mult_209_n2219), .A2(DP_mult_209_n1698), 
        .B1(DP_mult_209_n1993), .B2(DP_mult_209_n1697), .ZN(DP_mult_209_n1401)
         );
  OAI22_X1 DP_mult_209_U2327 ( .A1(DP_mult_209_n2023), .A2(DP_mult_209_n1696), 
        .B1(DP_mult_209_n2245), .B2(DP_mult_209_n1695), .ZN(DP_mult_209_n1399)
         );
  OAI22_X1 DP_mult_209_U2326 ( .A1(DP_mult_209_n2219), .A2(DP_mult_209_n1701), 
        .B1(DP_mult_209_n1700), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1404)
         );
  OAI22_X1 DP_mult_209_U2325 ( .A1(DP_mult_209_n2023), .A2(DP_mult_209_n1704), 
        .B1(DP_mult_209_n2245), .B2(DP_mult_209_n1703), .ZN(DP_mult_209_n1407)
         );
  OAI22_X1 DP_mult_209_U2324 ( .A1(DP_mult_209_n2023), .A2(DP_mult_209_n1694), 
        .B1(DP_mult_209_n1993), .B2(DP_mult_209_n1693), .ZN(DP_mult_209_n1397)
         );
  OAI22_X1 DP_mult_209_U2323 ( .A1(DP_mult_209_n2219), .A2(DP_mult_209_n1695), 
        .B1(DP_mult_209_n1694), .B2(DP_mult_209_n1993), .ZN(DP_mult_209_n1398)
         );
  OAI21_X1 DP_mult_209_U2322 ( .B1(DP_mult_209_n2153), .B2(DP_mult_209_n1955), 
        .A(DP_mult_209_n2313), .ZN(DP_mult_209_n1290) );
  NOR2_X1 DP_mult_209_U2321 ( .A1(DP_mult_209_n2145), .A2(DP_mult_209_n547), 
        .ZN(DP_mult_209_n540) );
  OAI21_X1 DP_mult_209_U2320 ( .B1(DP_mult_209_n2221), .B2(DP_mult_209_n2189), 
        .A(DP_mult_209_n2308), .ZN(DP_mult_209_n1410) );
  OAI21_X1 DP_mult_209_U2319 ( .B1(DP_mult_209_n2081), .B2(DP_mult_209_n564), 
        .A(DP_mult_209_n559), .ZN(DP_mult_209_n553) );
  INV_X1 DP_mult_209_U2318 ( .A(DP_mult_209_n558), .ZN(DP_mult_209_n675) );
  AOI21_X1 DP_mult_209_U2317 ( .B1(DP_mult_209_n565), .B2(DP_mult_209_n552), 
        .A(DP_mult_209_n2124), .ZN(DP_mult_209_n551) );
  XNOR2_X1 DP_mult_209_U2316 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2291), .ZN(
        DP_mult_209_n1567) );
  XNOR2_X1 DP_mult_209_U2315 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2291), .ZN(
        DP_mult_209_n1569) );
  XNOR2_X1 DP_mult_209_U2314 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2291), .ZN(
        DP_mult_209_n1565) );
  XNOR2_X1 DP_mult_209_U2313 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2291), .ZN(
        DP_mult_209_n1563) );
  XNOR2_X1 DP_mult_209_U2312 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2291), .ZN(
        DP_mult_209_n1561) );
  XNOR2_X1 DP_mult_209_U2311 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2291), .ZN(
        DP_mult_209_n1559) );
  INV_X1 DP_mult_209_U2310 ( .A(DP_mult_209_n2108), .ZN(DP_mult_209_n492) );
  OAI21_X1 DP_mult_209_U2309 ( .B1(DP_mult_209_n456), .B2(DP_mult_209_n481), 
        .A(DP_mult_209_n457), .ZN(DP_mult_209_n455) );
  INV_X1 DP_mult_209_U2308 ( .A(DP_mult_209_n2149), .ZN(DP_mult_209_n565) );
  NAND2_X1 DP_mult_209_U2307 ( .A1(DP_mult_209_n897), .A2(DP_mult_209_n918), 
        .ZN(DP_mult_209_n535) );
  AOI21_X1 DP_mult_209_U2306 ( .B1(DP_mult_209_n2131), .B2(DP_mult_209_n2057), 
        .A(DP_mult_209_n512), .ZN(DP_mult_209_n2202) );
  INV_X1 DP_mult_209_U2305 ( .A(DP_mult_209_n2223), .ZN(DP_mult_209_n2222) );
  NAND2_X1 DP_mult_209_U2304 ( .A1(DP_mult_209_n588), .A2(DP_mult_209_n2168), 
        .ZN(DP_mult_209_n582) );
  AOI21_X1 DP_mult_209_U2303 ( .B1(DP_mult_209_n589), .B2(DP_mult_209_n2168), 
        .A(DP_mult_209_n1978), .ZN(DP_mult_209_n583) );
  NAND2_X1 DP_mult_209_U2302 ( .A1(DP_mult_209_n1003), .A2(DP_mult_209_n1020), 
        .ZN(DP_mult_209_n570) );
  NAND2_X1 DP_mult_209_U2301 ( .A1(DP_mult_209_n2176), .A2(DP_mult_209_n2174), 
        .ZN(DP_mult_209_n599) );
  INV_X1 DP_mult_209_U2300 ( .A(DP_mult_209_n277), .ZN(DP_mult_209_n2223) );
  OAI22_X1 DP_mult_209_U2299 ( .A1(DP_mult_209_n2214), .A2(DP_mult_209_n1624), 
        .B1(DP_mult_209_n1623), .B2(DP_mult_209_n2238), .ZN(DP_mult_209_n1330)
         );
  OAI22_X1 DP_mult_209_U2298 ( .A1(DP_mult_209_n2052), .A2(DP_mult_209_n1622), 
        .B1(DP_mult_209_n1621), .B2(DP_mult_209_n2237), .ZN(DP_mult_209_n1328)
         );
  OAI22_X1 DP_mult_209_U2297 ( .A1(DP_mult_209_n2052), .A2(DP_mult_209_n1619), 
        .B1(DP_mult_209_n2237), .B2(DP_mult_209_n1618), .ZN(DP_mult_209_n1325)
         );
  OAI22_X1 DP_mult_209_U2296 ( .A1(DP_mult_209_n2213), .A2(DP_mult_209_n1625), 
        .B1(DP_mult_209_n2237), .B2(DP_mult_209_n1624), .ZN(DP_mult_209_n1331)
         );
  OAI22_X1 DP_mult_209_U2295 ( .A1(DP_mult_209_n2213), .A2(DP_mult_209_n1626), 
        .B1(DP_mult_209_n1625), .B2(DP_mult_209_n2237), .ZN(DP_mult_209_n1332)
         );
  OAI22_X1 DP_mult_209_U2294 ( .A1(DP_mult_209_n2011), .A2(DP_mult_209_n1627), 
        .B1(DP_mult_209_n2238), .B2(DP_mult_209_n1626), .ZN(DP_mult_209_n1333)
         );
  OAI22_X1 DP_mult_209_U2293 ( .A1(DP_mult_209_n2011), .A2(DP_mult_209_n1621), 
        .B1(DP_mult_209_n2238), .B2(DP_mult_209_n1620), .ZN(DP_mult_209_n1327)
         );
  OAI22_X1 DP_mult_209_U2292 ( .A1(DP_mult_209_n2213), .A2(DP_mult_209_n1623), 
        .B1(DP_mult_209_n2238), .B2(DP_mult_209_n1622), .ZN(DP_mult_209_n1329)
         );
  OAI22_X1 DP_mult_209_U2291 ( .A1(DP_mult_209_n1991), .A2(DP_mult_209_n1629), 
        .B1(DP_mult_209_n2237), .B2(DP_mult_209_n1628), .ZN(DP_mult_209_n1335)
         );
  OAI22_X1 DP_mult_209_U2290 ( .A1(DP_mult_209_n1992), .A2(DP_mult_209_n1620), 
        .B1(DP_mult_209_n1619), .B2(DP_mult_209_n2237), .ZN(DP_mult_209_n1326)
         );
  NOR2_X1 DP_mult_209_U2289 ( .A1(DP_mult_209_n2010), .A2(DP_mult_209_n2098), 
        .ZN(DP_mult_209_n545) );
  OAI21_X1 DP_mult_209_U2288 ( .B1(DP_mult_209_n1984), .B2(DP_mult_209_n2098), 
        .A(DP_mult_209_n550), .ZN(DP_mult_209_n546) );
  INV_X1 DP_mult_209_U2287 ( .A(DP_mult_209_n537), .ZN(DP_mult_209_n536) );
  NAND2_X1 DP_mult_209_U2286 ( .A1(DP_mult_209_n821), .A2(DP_mult_209_n838), 
        .ZN(DP_mult_209_n503) );
  NAND3_X1 DP_mult_209_U2285 ( .A1(DP_mult_209_n2199), .A2(DP_mult_209_n2200), 
        .A3(DP_mult_209_n2201), .ZN(DP_mult_209_n822) );
  NAND2_X1 DP_mult_209_U2284 ( .A1(DP_mult_209_n844), .A2(DP_mult_209_n827), 
        .ZN(DP_mult_209_n2201) );
  NAND2_X1 DP_mult_209_U2283 ( .A1(DP_mult_209_n2032), .A2(DP_mult_209_n827), 
        .ZN(DP_mult_209_n2200) );
  NAND2_X1 DP_mult_209_U2282 ( .A1(DP_mult_209_n2032), .A2(DP_mult_209_n844), 
        .ZN(DP_mult_209_n2199) );
  XOR2_X1 DP_mult_209_U2281 ( .A(DP_mult_209_n2033), .B(DP_mult_209_n2198), 
        .Z(DP_mult_209_n823) );
  XOR2_X1 DP_mult_209_U2280 ( .A(DP_mult_209_n844), .B(DP_mult_209_n827), .Z(
        DP_mult_209_n2198) );
  OAI21_X1 DP_mult_209_U2279 ( .B1(DP_mult_209_n631), .B2(DP_mult_209_n634), 
        .A(DP_mult_209_n632), .ZN(DP_mult_209_n630) );
  NOR2_X1 DP_mult_209_U2278 ( .A1(DP_mult_209_n633), .A2(DP_mult_209_n631), 
        .ZN(DP_mult_209_n629) );
  XNOR2_X1 DP_mult_209_U2277 ( .A(DP_mult_209_n522), .B(DP_mult_209_n319), 
        .ZN(DP_pipe0_coeff_pipe03[5]) );
  AOI21_X1 DP_mult_209_U2276 ( .B1(DP_mult_209_n401), .B2(DP_mult_209_n2171), 
        .A(DP_mult_209_n394), .ZN(DP_mult_209_n390) );
  INV_X1 DP_mult_209_U2275 ( .A(DP_mult_209_n383), .ZN(DP_mult_209_n381) );
  INV_X1 DP_mult_209_U2274 ( .A(DP_mult_209_n401), .ZN(DP_mult_209_n399) );
  OAI22_X1 DP_mult_209_U2273 ( .A1(DP_mult_209_n2193), .A2(DP_mult_209_n1711), 
        .B1(DP_mult_209_n1958), .B2(DP_mult_209_n1710), .ZN(DP_mult_209_n1413)
         );
  OAI22_X1 DP_mult_209_U2272 ( .A1(DP_mult_209_n2089), .A2(DP_mult_209_n1709), 
        .B1(DP_mult_209_n1959), .B2(DP_mult_209_n1708), .ZN(DP_mult_209_n1411)
         );
  OAI22_X1 DP_mult_209_U2271 ( .A1(DP_mult_209_n2193), .A2(DP_mult_209_n1713), 
        .B1(DP_mult_209_n1958), .B2(DP_mult_209_n1712), .ZN(DP_mult_209_n1415)
         );
  OAI22_X1 DP_mult_209_U2270 ( .A1(DP_mult_209_n2089), .A2(DP_mult_209_n1717), 
        .B1(DP_mult_209_n1959), .B2(DP_mult_209_n1716), .ZN(DP_mult_209_n1419)
         );
  XNOR2_X1 DP_mult_209_U2269 ( .A(DP_mult_209_n515), .B(DP_mult_209_n318), 
        .ZN(DP_pipe0_coeff_pipe03[6]) );
  NAND2_X1 DP_mult_209_U2268 ( .A1(DP_mult_209_n919), .A2(DP_mult_209_n940), 
        .ZN(DP_mult_209_n543) );
  XNOR2_X1 DP_mult_209_U2267 ( .A(DP_mult_209_n504), .B(DP_mult_209_n317), 
        .ZN(DP_pipe0_coeff_pipe03[7]) );
  CLKBUF_X1 DP_mult_209_U2266 ( .A(DP_mult_209_n2202), .Z(DP_mult_209_n2197)
         );
  XNOR2_X1 DP_mult_209_U2265 ( .A(DP_mult_209_n497), .B(DP_mult_209_n316), 
        .ZN(DP_pipe0_coeff_pipe03[8]) );
  XNOR2_X1 DP_mult_209_U2264 ( .A(DP_mult_209_n486), .B(DP_mult_209_n315), 
        .ZN(DP_pipe0_coeff_pipe03[9]) );
  XNOR2_X1 DP_mult_209_U2263 ( .A(DP_mult_209_n475), .B(DP_mult_209_n314), 
        .ZN(DP_pipe0_coeff_pipe03[10]) );
  NOR2_X1 DP_mult_209_U2262 ( .A1(DP_mult_209_n571), .A2(DP_mult_209_n2041), 
        .ZN(DP_mult_209_n567) );
  INV_X1 DP_mult_209_U2261 ( .A(DP_mult_209_n2086), .ZN(DP_mult_209_n2206) );
  OAI21_X1 DP_mult_209_U2260 ( .B1(DP_mult_209_n600), .B2(DP_mult_209_n597), 
        .A(DP_mult_209_n598), .ZN(DP_mult_209_n596) );
  INV_X1 DP_mult_209_U2259 ( .A(DP_mult_209_n1975), .ZN(DP_mult_209_n2220) );
  OAI21_X1 DP_mult_209_U2258 ( .B1(DP_mult_209_n1989), .B2(DP_mult_209_n2017), 
        .A(DP_mult_209_n2315), .ZN(DP_mult_209_n1242) );
  OAI22_X1 DP_mult_209_U2257 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1492), 
        .B1(DP_mult_209_n2045), .B2(DP_mult_209_n1491), .ZN(DP_mult_209_n1203)
         );
  OAI22_X1 DP_mult_209_U2256 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1490), 
        .B1(DP_mult_209_n2045), .B2(DP_mult_209_n1489), .ZN(DP_mult_209_n1201)
         );
  OAI22_X1 DP_mult_209_U2255 ( .A1(DP_mult_209_n2044), .A2(DP_mult_209_n1486), 
        .B1(DP_mult_209_n2064), .B2(DP_mult_209_n1485), .ZN(DP_mult_209_n1197)
         );
  OAI22_X1 DP_mult_209_U2254 ( .A1(DP_mult_209_n1938), .A2(DP_mult_209_n1488), 
        .B1(DP_mult_209_n2064), .B2(DP_mult_209_n1487), .ZN(DP_mult_209_n1199)
         );
  OAI22_X1 DP_mult_209_U2253 ( .A1(DP_mult_209_n1938), .A2(DP_mult_209_n1484), 
        .B1(DP_mult_209_n2064), .B2(DP_mult_209_n1483), .ZN(DP_mult_209_n1195)
         );
  NOR2_X1 DP_mult_209_U2252 ( .A1(DP_mult_209_n420), .A2(DP_mult_209_n347), 
        .ZN(DP_mult_209_n345) );
  AOI21_X1 DP_mult_209_U2251 ( .B1(DP_mult_209_n629), .B2(DP_mult_209_n635), 
        .A(DP_mult_209_n630), .ZN(DP_mult_209_n628) );
  OAI22_X1 DP_mult_209_U2250 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1517), 
        .B1(DP_mult_209_n2227), .B2(DP_mult_209_n1516), .ZN(DP_mult_209_n1227)
         );
  OAI22_X1 DP_mult_209_U2249 ( .A1(DP_mult_209_n2015), .A2(DP_mult_209_n1509), 
        .B1(DP_mult_209_n2228), .B2(DP_mult_209_n1508), .ZN(DP_mult_209_n1219)
         );
  OAI22_X1 DP_mult_209_U2248 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1515), 
        .B1(DP_mult_209_n2228), .B2(DP_mult_209_n1514), .ZN(DP_mult_209_n1225)
         );
  OAI22_X1 DP_mult_209_U2247 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1511), 
        .B1(DP_mult_209_n2227), .B2(DP_mult_209_n1510), .ZN(DP_mult_209_n1221)
         );
  OAI22_X1 DP_mult_209_U2246 ( .A1(DP_mult_209_n2101), .A2(DP_mult_209_n1513), 
        .B1(DP_mult_209_n2228), .B2(DP_mult_209_n1512), .ZN(DP_mult_209_n1223)
         );
  INV_X1 DP_mult_209_U2245 ( .A(DP_mult_209_n521), .ZN(DP_mult_209_n519) );
  NAND2_X1 DP_mult_209_U2244 ( .A1(DP_mult_209_n2137), .A2(DP_mult_209_n521), 
        .ZN(DP_mult_209_n319) );
  NOR2_X1 DP_mult_209_U2243 ( .A1(DP_mult_209_n839), .A2(DP_mult_209_n856), 
        .ZN(DP_mult_209_n513) );
  INV_X1 DP_mult_209_U2242 ( .A(DP_mult_209_n874), .ZN(DP_mult_209_n875) );
  NAND2_X1 DP_mult_209_U2241 ( .A1(DP_mult_209_n963), .A2(DP_mult_209_n982), 
        .ZN(DP_mult_209_n559) );
  INV_X1 DP_mult_209_U2240 ( .A(DP_mult_209_n267), .ZN(DP_mult_209_n2232) );
  INV_X1 DP_mult_209_U2239 ( .A(DP_mult_209_n2260), .ZN(DP_mult_209_n2257) );
  BUF_X1 DP_mult_209_U2238 ( .A(DP_mult_209_n283), .Z(DP_mult_209_n2203) );
  XNOR2_X1 DP_mult_209_U2237 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1482) );
  XNOR2_X1 DP_mult_209_U2236 ( .A(DP_mult_209_n448), .B(DP_mult_209_n312), 
        .ZN(DP_pipe0_coeff_pipe03[12]) );
  NAND2_X1 DP_mult_209_U2235 ( .A1(DP_mult_209_n2167), .A2(DP_mult_209_n461), 
        .ZN(DP_mult_209_n313) );
  NAND2_X1 DP_mult_209_U2234 ( .A1(DP_mult_209_n667), .A2(DP_mult_209_n496), 
        .ZN(DP_mult_209_n316) );
  NAND2_X1 DP_mult_209_U2233 ( .A1(DP_mult_209_n668), .A2(DP_mult_209_n503), 
        .ZN(DP_mult_209_n317) );
  NAND2_X1 DP_mult_209_U2232 ( .A1(DP_mult_209_n2090), .A2(DP_mult_209_n514), 
        .ZN(DP_mult_209_n318) );
  NAND2_X1 DP_mult_209_U2231 ( .A1(DP_mult_209_n671), .A2(DP_mult_209_n532), 
        .ZN(DP_mult_209_n320) );
  INV_X1 DP_mult_209_U2230 ( .A(DP_coeffs_ff_int[95]), .ZN(DP_mult_209_n251)
         );
  XNOR2_X1 DP_mult_209_U2229 ( .A(DP_mult_209_n2300), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1530) );
  XNOR2_X1 DP_mult_209_U2228 ( .A(DP_mult_209_n2287), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1605) );
  XNOR2_X1 DP_mult_209_U2227 ( .A(DP_mult_209_n2272), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1680) );
  XNOR2_X1 DP_mult_209_U2226 ( .A(DP_mult_209_n2258), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1755) );
  OAI22_X1 DP_mult_209_U2225 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1778), 
        .B1(DP_mult_209_n1777), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1479)
         );
  XNOR2_X1 DP_mult_209_U2224 ( .A(DP_mult_209_n2253), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1780) );
  OAI22_X1 DP_mult_209_U2223 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1780), 
        .B1(DP_mult_209_n1779), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1481)
         );
  INV_X1 DP_mult_209_U2222 ( .A(DP_mult_209_n297), .ZN(DP_mult_209_n2205) );
  XNOR2_X1 DP_mult_209_U2221 ( .A(DP_mult_209_n2281), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1630) );
  INV_X1 DP_mult_209_U2220 ( .A(DP_mult_209_n1757), .ZN(DP_mult_209_n2306) );
  OAI21_X1 DP_mult_209_U2219 ( .B1(DP_coeffs_ff_int[95]), .B2(
        DP_mult_209_n2184), .A(DP_mult_209_n2306), .ZN(DP_mult_209_n1458) );
  NAND2_X1 DP_mult_209_U2218 ( .A1(DP_mult_209_n666), .A2(DP_mult_209_n481), 
        .ZN(DP_mult_209_n315) );
  AOI21_X1 DP_mult_209_U2217 ( .B1(DP_mult_209_n565), .B2(DP_mult_209_n545), 
        .A(DP_mult_209_n546), .ZN(DP_mult_209_n544) );
  AOI21_X1 DP_mult_209_U2216 ( .B1(DP_mult_209_n565), .B2(DP_mult_209_n561), 
        .A(DP_mult_209_n562), .ZN(DP_mult_209_n560) );
  INV_X1 DP_mult_209_U2215 ( .A(DP_mult_209_n259), .ZN(DP_mult_209_n2244) );
  INV_X1 DP_mult_209_U2214 ( .A(DP_coeffs_ff_int[72]), .ZN(DP_mult_209_n2305)
         );
  XNOR2_X1 DP_mult_209_U2213 ( .A(DP_pipe03[21]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1484) );
  XNOR2_X1 DP_mult_209_U2212 ( .A(DP_pipe03[19]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1486) );
  XNOR2_X1 DP_mult_209_U2211 ( .A(DP_pipe03[15]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1490) );
  XNOR2_X1 DP_mult_209_U2210 ( .A(DP_pipe03[17]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1488) );
  XNOR2_X1 DP_mult_209_U2209 ( .A(DP_pipe03[13]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1492) );
  XNOR2_X1 DP_mult_209_U2208 ( .A(DP_pipe03[11]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1494) );
  AND2_X1 DP_mult_209_U2207 ( .A1(DP_mult_209_n1817), .A2(DP_mult_209_n2249), 
        .ZN(DP_mult_209_n2184) );
  XNOR2_X1 DP_mult_209_U2206 ( .A(DP_mult_209_n2277), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1655) );
  XNOR2_X1 DP_mult_209_U2205 ( .A(DP_mult_209_n2263), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1730) );
  OAI22_X1 DP_mult_209_U2204 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1776), 
        .B1(DP_mult_209_n1775), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1477)
         );
  XNOR2_X1 DP_mult_209_U2203 ( .A(DP_mult_209_n2291), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1580) );
  XNOR2_X1 DP_mult_209_U2202 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2035), .ZN(
        DP_mult_209_n1625) );
  XNOR2_X1 DP_mult_209_U2201 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2285), .ZN(
        DP_mult_209_n1600) );
  XNOR2_X1 DP_mult_209_U2200 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1500) );
  XNOR2_X1 DP_mult_209_U2199 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1673) );
  XNOR2_X1 DP_mult_209_U2198 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2281), .ZN(
        DP_mult_209_n1623) );
  XNOR2_X1 DP_mult_209_U2197 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2261), .ZN(
        DP_mult_209_n1727) );
  XNOR2_X1 DP_mult_209_U2196 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2095), .ZN(
        DP_mult_209_n1548) );
  XNOR2_X1 DP_mult_209_U2195 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2285), .ZN(
        DP_mult_209_n1602) );
  XNOR2_X1 DP_mult_209_U2194 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1648) );
  XNOR2_X1 DP_mult_209_U2193 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2298), .ZN(
        DP_mult_209_n1523) );
  XNOR2_X1 DP_mult_209_U2192 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1502) );
  XNOR2_X1 DP_mult_209_U2191 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2298), .ZN(
        DP_mult_209_n1525) );
  XNOR2_X1 DP_mult_209_U2190 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1652) );
  XNOR2_X1 DP_mult_209_U2189 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1498) );
  XNOR2_X1 DP_mult_209_U2188 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1677) );
  XNOR2_X1 DP_mult_209_U2187 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2058), .ZN(
        DP_mult_209_n1577) );
  XNOR2_X1 DP_mult_209_U2186 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2281), .ZN(
        DP_mult_209_n1627) );
  XNOR2_X1 DP_mult_209_U2185 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2267), .ZN(
        DP_mult_209_n1700) );
  XNOR2_X1 DP_mult_209_U2184 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2261), .ZN(
        DP_mult_209_n1725) );
  XNOR2_X1 DP_mult_209_U2183 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2256), .ZN(
        DP_mult_209_n1752) );
  XNOR2_X1 DP_mult_209_U2182 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2256), .ZN(
        DP_mult_209_n1748) );
  XNOR2_X1 DP_mult_209_U2181 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2298), .ZN(
        DP_mult_209_n1527) );
  XNOR2_X1 DP_mult_209_U2180 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2290), .ZN(
        DP_mult_209_n1573) );
  XNOR2_X1 DP_mult_209_U2179 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2261), .ZN(
        DP_mult_209_n1723) );
  XNOR2_X1 DP_mult_209_U2178 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2256), .ZN(
        DP_mult_209_n1750) );
  XNOR2_X1 DP_mult_209_U2177 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2095), .ZN(
        DP_mult_209_n1550) );
  XNOR2_X1 DP_mult_209_U2176 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2094), .ZN(
        DP_mult_209_n1552) );
  XNOR2_X1 DP_mult_209_U2175 ( .A(DP_pipe03[3]), .B(DP_mult_209_n2267), .ZN(
        DP_mult_209_n1702) );
  XNOR2_X1 DP_mult_209_U2174 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1675) );
  XNOR2_X1 DP_mult_209_U2173 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2267), .ZN(
        DP_mult_209_n1698) );
  XNOR2_X1 DP_mult_209_U2172 ( .A(DP_pipe03[7]), .B(DP_mult_209_n2285), .ZN(
        DP_mult_209_n1598) );
  XNOR2_X1 DP_mult_209_U2171 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2058), .ZN(
        DP_mult_209_n1575) );
  XNOR2_X1 DP_mult_209_U2170 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2035), .ZN(
        DP_mult_209_n1629) );
  XNOR2_X1 DP_mult_209_U2169 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2267), .ZN(
        DP_mult_209_n1704) );
  XNOR2_X1 DP_mult_209_U2168 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2261), .ZN(
        DP_mult_209_n1729) );
  XNOR2_X1 DP_mult_209_U2167 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2290), .ZN(
        DP_mult_209_n1579) );
  XNOR2_X1 DP_mult_209_U2166 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1504) );
  XNOR2_X1 DP_mult_209_U2165 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2256), .ZN(
        DP_mult_209_n1754) );
  XNOR2_X1 DP_mult_209_U2164 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2285), .ZN(
        DP_mult_209_n1604) );
  XNOR2_X1 DP_mult_209_U2163 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1654) );
  XNOR2_X1 DP_mult_209_U2162 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2094), .ZN(
        DP_mult_209_n1554) );
  XNOR2_X1 DP_mult_209_U2161 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2298), .ZN(
        DP_mult_209_n1529) );
  XNOR2_X1 DP_mult_209_U2160 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1679) );
  XNOR2_X1 DP_mult_209_U2159 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2298), .ZN(
        DP_mult_209_n1521) );
  XNOR2_X1 DP_mult_209_U2158 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2303), .ZN(
        DP_mult_209_n1496) );
  XNOR2_X1 DP_mult_209_U2157 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2261), .ZN(
        DP_mult_209_n1721) );
  XNOR2_X1 DP_mult_209_U2156 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1671) );
  XNOR2_X1 DP_mult_209_U2155 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2095), .ZN(
        DP_mult_209_n1546) );
  XNOR2_X1 DP_mult_209_U2154 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2266), .ZN(
        DP_mult_209_n1696) );
  XNOR2_X1 DP_mult_209_U2153 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2285), .ZN(
        DP_mult_209_n1596) );
  XNOR2_X1 DP_mult_209_U2152 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2035), .ZN(
        DP_mult_209_n1621) );
  XNOR2_X1 DP_mult_209_U2151 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2256), .ZN(
        DP_mult_209_n1746) );
  XNOR2_X1 DP_mult_209_U2150 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2058), .ZN(
        DP_mult_209_n1571) );
  XNOR2_X1 DP_mult_209_U2149 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1646) );
  XNOR2_X1 DP_mult_209_U2148 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2299), .ZN(
        DP_mult_209_n1507) );
  XNOR2_X1 DP_mult_209_U2147 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2285), .ZN(
        DP_mult_209_n1582) );
  XNOR2_X1 DP_mult_209_U2146 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2036), .ZN(
        DP_mult_209_n1607) );
  XNOR2_X1 DP_mult_209_U2145 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2094), .ZN(
        DP_mult_209_n1532) );
  XNOR2_X1 DP_mult_209_U2144 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2261), .ZN(
        DP_mult_209_n1707) );
  XNOR2_X1 DP_mult_209_U2143 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2291), .ZN(
        DP_mult_209_n1557) );
  XNOR2_X1 DP_mult_209_U2142 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2271), .ZN(
        DP_mult_209_n1657) );
  XNOR2_X1 DP_mult_209_U2141 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2275), .ZN(
        DP_mult_209_n1632) );
  XNOR2_X1 DP_mult_209_U2140 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2266), .ZN(
        DP_mult_209_n1682) );
  XNOR2_X1 DP_mult_209_U2139 ( .A(DP_mult_209_n2295), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1555) );
  XNOR2_X1 DP_mult_209_U2138 ( .A(DP_mult_209_n2268), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1705) );
  XNOR2_X1 DP_mult_209_U2137 ( .A(DP_pipe03[1]), .B(DP_mult_209_n2251), .ZN(
        DP_mult_209_n1779) );
  XNOR2_X1 DP_mult_209_U2136 ( .A(DP_mult_209_n2304), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1483) );
  XNOR2_X1 DP_mult_209_U2135 ( .A(DP_mult_209_n2295), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1535) );
  XNOR2_X1 DP_mult_209_U2134 ( .A(DP_mult_209_n2291), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1560) );
  XNOR2_X1 DP_mult_209_U2133 ( .A(DP_mult_209_n2300), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1514) );
  XNOR2_X1 DP_mult_209_U2132 ( .A(DP_mult_209_n2287), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1589) );
  XNOR2_X1 DP_mult_209_U2131 ( .A(DP_mult_209_n2304), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1487) );
  XNOR2_X1 DP_mult_209_U2130 ( .A(DP_mult_209_n2300), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1510) );
  XNOR2_X1 DP_mult_209_U2129 ( .A(DP_mult_209_n2304), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1485) );
  XNOR2_X1 DP_mult_209_U2128 ( .A(DP_mult_209_n2294), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1537) );
  XNOR2_X1 DP_mult_209_U2127 ( .A(DP_mult_209_n2262), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1720) );
  XNOR2_X1 DP_mult_209_U2126 ( .A(DP_mult_209_n2277), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1635) );
  XNOR2_X1 DP_mult_209_U2125 ( .A(DP_mult_209_n2294), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1543) );
  XNOR2_X1 DP_mult_209_U2124 ( .A(DP_mult_209_n2268), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1685) );
  XNOR2_X1 DP_mult_209_U2123 ( .A(DP_mult_209_n2300), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1508) );
  XNOR2_X1 DP_mult_209_U2122 ( .A(DP_mult_209_n2299), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1518) );
  XNOR2_X1 DP_mult_209_U2121 ( .A(DP_mult_209_n2287), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1583) );
  XNOR2_X1 DP_mult_209_U2120 ( .A(DP_mult_209_n2290), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1562) );
  XNOR2_X1 DP_mult_209_U2119 ( .A(DP_mult_209_n1952), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1660) );
  XNOR2_X1 DP_mult_209_U2118 ( .A(DP_mult_209_n2280), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1612) );
  XNOR2_X1 DP_mult_209_U2117 ( .A(DP_mult_209_n2295), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1533) );
  XNOR2_X1 DP_mult_209_U2116 ( .A(DP_mult_209_n2299), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1520) );
  XNOR2_X1 DP_mult_209_U2115 ( .A(DP_mult_209_n2304), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1489) );
  XNOR2_X1 DP_mult_209_U2114 ( .A(DP_mult_209_n2058), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1570) );
  XNOR2_X1 DP_mult_209_U2113 ( .A(DP_mult_209_n2291), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1564) );
  XNOR2_X1 DP_mult_209_U2112 ( .A(DP_mult_209_n2304), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1493) );
  XNOR2_X1 DP_mult_209_U2111 ( .A(DP_mult_209_n2281), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1610) );
  XNOR2_X1 DP_mult_209_U2110 ( .A(DP_mult_209_n2286), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1587) );
  XNOR2_X1 DP_mult_209_U2109 ( .A(DP_mult_209_n2304), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1495) );
  XNOR2_X1 DP_mult_209_U2108 ( .A(DP_mult_209_n2281), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1608) );
  XNOR2_X1 DP_mult_209_U2107 ( .A(DP_mult_209_n2272), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1670) );
  XNOR2_X1 DP_mult_209_U2106 ( .A(DP_mult_209_n2267), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1687) );
  XNOR2_X1 DP_mult_209_U2105 ( .A(DP_mult_209_n2268), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1689) );
  XNOR2_X1 DP_mult_209_U2104 ( .A(DP_mult_209_n2277), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1639) );
  XNOR2_X1 DP_mult_209_U2103 ( .A(DP_mult_209_n2299), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1512) );
  XNOR2_X1 DP_mult_209_U2102 ( .A(DP_mult_209_n2287), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1585) );
  XNOR2_X1 DP_mult_209_U2101 ( .A(DP_mult_209_n2295), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1539) );
  XNOR2_X1 DP_mult_209_U2100 ( .A(DP_mult_209_n2291), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1558) );
  XNOR2_X1 DP_mult_209_U2099 ( .A(DP_mult_209_n1953), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1674) );
  XNOR2_X1 DP_mult_209_U2098 ( .A(DP_mult_209_n2280), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1620) );
  XNOR2_X1 DP_mult_209_U2097 ( .A(DP_mult_209_n2286), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1593) );
  XNOR2_X1 DP_mult_209_U2096 ( .A(DP_mult_209_n2262), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1718) );
  XNOR2_X1 DP_mult_209_U2095 ( .A(DP_mult_209_n2280), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1626) );
  XNOR2_X1 DP_mult_209_U2094 ( .A(DP_mult_209_n2281), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1614) );
  XNOR2_X1 DP_mult_209_U2093 ( .A(DP_mult_209_n2258), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1739) );
  XNOR2_X1 DP_mult_209_U2092 ( .A(DP_mult_209_n2267), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1695) );
  XNOR2_X1 DP_mult_209_U2091 ( .A(DP_mult_209_n2294), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1545) );
  XNOR2_X1 DP_mult_209_U2090 ( .A(DP_mult_209_n2263), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1708) );
  XNOR2_X1 DP_mult_209_U2089 ( .A(DP_mult_209_n2286), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1601) );
  XNOR2_X1 DP_mult_209_U2088 ( .A(DP_mult_209_n2273), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1662) );
  XNOR2_X1 DP_mult_209_U2087 ( .A(DP_mult_209_n1953), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1664) );
  XNOR2_X1 DP_mult_209_U2086 ( .A(DP_mult_209_n2304), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1501) );
  XNOR2_X1 DP_mult_209_U2085 ( .A(DP_mult_209_n2277), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1633) );
  XNOR2_X1 DP_mult_209_U2084 ( .A(DP_mult_209_n2276), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1637) );
  XNOR2_X1 DP_mult_209_U2083 ( .A(DP_mult_209_n2276), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1651) );
  XNOR2_X1 DP_mult_209_U2082 ( .A(DP_mult_209_n2258), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1735) );
  XNOR2_X1 DP_mult_209_U2081 ( .A(DP_mult_209_n2263), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1710) );
  XNOR2_X1 DP_mult_209_U2080 ( .A(DP_mult_209_n2276), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1649) );
  XNOR2_X1 DP_mult_209_U2079 ( .A(DP_mult_209_n2280), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1624) );
  XNOR2_X1 DP_mult_209_U2078 ( .A(DP_mult_209_n2280), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1618) );
  XNOR2_X1 DP_mult_209_U2077 ( .A(DP_mult_209_n2304), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1499) );
  XNOR2_X1 DP_mult_209_U2076 ( .A(DP_mult_209_n2294), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1549) );
  XNOR2_X1 DP_mult_209_U2075 ( .A(DP_mult_209_n2058), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1568) );
  XNOR2_X1 DP_mult_209_U2074 ( .A(DP_mult_209_n2299), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1524) );
  XNOR2_X1 DP_mult_209_U2073 ( .A(DP_mult_209_n2262), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1726) );
  XNOR2_X1 DP_mult_209_U2072 ( .A(DP_mult_209_n2286), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1595) );
  XNOR2_X1 DP_mult_209_U2071 ( .A(DP_mult_209_n2267), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1701) );
  XNOR2_X1 DP_mult_209_U2070 ( .A(DP_mult_209_n2266), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1693) );
  XNOR2_X1 DP_mult_209_U2069 ( .A(DP_mult_209_n2273), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1658) );
  XNOR2_X1 DP_mult_209_U2068 ( .A(DP_mult_209_n2058), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1574) );
  XNOR2_X1 DP_mult_209_U2067 ( .A(DP_mult_209_n2262), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1712) );
  XNOR2_X1 DP_mult_209_U2066 ( .A(DP_mult_209_n2258), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1733) );
  XNOR2_X1 DP_mult_209_U2065 ( .A(DP_mult_209_n2276), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1643) );
  XNOR2_X1 DP_mult_209_U2064 ( .A(DP_mult_209_n2294), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1551) );
  XNOR2_X1 DP_mult_209_U2063 ( .A(DP_mult_209_n2276), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1645) );
  XNOR2_X1 DP_mult_209_U2062 ( .A(DP_mult_209_n2262), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1724) );
  XNOR2_X1 DP_mult_209_U2061 ( .A(DP_mult_209_n2299), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1526) );
  XNOR2_X1 DP_mult_209_U2060 ( .A(DP_mult_209_n1942), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1743) );
  XNOR2_X1 DP_mult_209_U2059 ( .A(DP_mult_209_n1952), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1676) );
  XNOR2_X1 DP_mult_209_U2058 ( .A(DP_mult_209_n2267), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1699) );
  XNOR2_X1 DP_mult_209_U2057 ( .A(DP_mult_209_n1942), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1745) );
  XNOR2_X1 DP_mult_209_U2056 ( .A(DP_mult_209_n1941), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1749) );
  XNOR2_X1 DP_mult_209_U2055 ( .A(DP_mult_209_n2286), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1599) );
  XNOR2_X1 DP_mult_209_U2054 ( .A(DP_mult_209_n2263), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1714) );
  XNOR2_X1 DP_mult_209_U2053 ( .A(DP_mult_209_n2290), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1576) );
  XNOR2_X1 DP_mult_209_U2052 ( .A(DP_mult_209_n2272), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1668) );
  XNOR2_X1 DP_mult_209_U2051 ( .A(DP_mult_209_n1942), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1751) );
  XNOR2_X1 DP_mult_209_U2050 ( .A(DP_mult_209_n1940), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1737) );
  XNOR2_X1 DP_mult_209_U2049 ( .A(DP_pipe03[9]), .B(DP_mult_209_n2251), .ZN(
        DP_mult_209_n1771) );
  XNOR2_X1 DP_mult_209_U2048 ( .A(DP_mult_209_n2291), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1566) );
  XNOR2_X1 DP_mult_209_U2047 ( .A(DP_mult_209_n2304), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1491) );
  XNOR2_X1 DP_mult_209_U2046 ( .A(DP_mult_209_n2294), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1541) );
  XNOR2_X1 DP_mult_209_U2045 ( .A(DP_mult_209_n2299), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1516) );
  XNOR2_X1 DP_mult_209_U2044 ( .A(DP_mult_209_n2262), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1716) );
  XNOR2_X1 DP_mult_209_U2043 ( .A(DP_mult_209_n2286), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1591) );
  XNOR2_X1 DP_mult_209_U2042 ( .A(DP_mult_209_n2294), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1547) );
  XNOR2_X1 DP_mult_209_U2041 ( .A(DP_mult_209_n1952), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1672) );
  XNOR2_X1 DP_mult_209_U2040 ( .A(DP_mult_209_n1942), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1753) );
  XNOR2_X1 DP_mult_209_U2039 ( .A(DP_mult_209_n2266), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1691) );
  XNOR2_X1 DP_mult_209_U2038 ( .A(DP_mult_209_n2299), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1522) );
  XNOR2_X1 DP_mult_209_U2037 ( .A(DP_mult_209_n2276), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1647) );
  XNOR2_X1 DP_mult_209_U2036 ( .A(DP_mult_209_n2280), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1616) );
  XNOR2_X1 DP_mult_209_U2035 ( .A(DP_mult_209_n2262), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1722) );
  XNOR2_X1 DP_mult_209_U2034 ( .A(DP_mult_209_n2262), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1728) );
  XNOR2_X1 DP_mult_209_U2033 ( .A(DP_mult_209_n2267), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1697) );
  XNOR2_X1 DP_mult_209_U2032 ( .A(DP_mult_209_n2286), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1603) );
  XNOR2_X1 DP_mult_209_U2031 ( .A(DP_mult_209_n2290), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1578) );
  XNOR2_X1 DP_mult_209_U2030 ( .A(DP_mult_209_n2286), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1597) );
  XNOR2_X1 DP_mult_209_U2029 ( .A(DP_mult_209_n1941), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1747) );
  XNOR2_X1 DP_mult_209_U2028 ( .A(DP_mult_209_n2291), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1572) );
  XNOR2_X1 DP_mult_209_U2027 ( .A(DP_mult_209_n2276), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1641) );
  XNOR2_X1 DP_mult_209_U2026 ( .A(DP_mult_209_n2304), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1503) );
  XNOR2_X1 DP_mult_209_U2025 ( .A(DP_mult_209_n2304), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1497) );
  XNOR2_X1 DP_mult_209_U2024 ( .A(DP_mult_209_n2299), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1528) );
  XNOR2_X1 DP_mult_209_U2023 ( .A(DP_mult_209_n1942), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1741) );
  XNOR2_X1 DP_mult_209_U2022 ( .A(DP_mult_209_n2294), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1553) );
  XNOR2_X1 DP_mult_209_U2021 ( .A(DP_mult_209_n2276), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1653) );
  XNOR2_X1 DP_mult_209_U2020 ( .A(DP_mult_209_n2280), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1622) );
  XNOR2_X1 DP_mult_209_U2019 ( .A(DP_mult_209_n1953), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1678) );
  XNOR2_X1 DP_mult_209_U2018 ( .A(DP_mult_209_n2280), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1628) );
  XNOR2_X1 DP_mult_209_U2017 ( .A(DP_mult_209_n2267), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1703) );
  XNOR2_X1 DP_mult_209_U2016 ( .A(DP_mult_209_n2253), .B(DP_pipe03[20]), .ZN(
        DP_mult_209_n1760) );
  XNOR2_X1 DP_mult_209_U2015 ( .A(DP_mult_209_n2253), .B(DP_pipe03[16]), .ZN(
        DP_mult_209_n1764) );
  XNOR2_X1 DP_mult_209_U2014 ( .A(DP_mult_209_n2253), .B(DP_pipe03[22]), .ZN(
        DP_mult_209_n1758) );
  XNOR2_X1 DP_mult_209_U2013 ( .A(DP_mult_209_n2252), .B(DP_pipe03[4]), .ZN(
        DP_mult_209_n1776) );
  XNOR2_X1 DP_mult_209_U2012 ( .A(DP_mult_209_n2252), .B(DP_pipe03[6]), .ZN(
        DP_mult_209_n1774) );
  XNOR2_X1 DP_mult_209_U2011 ( .A(DP_mult_209_n2252), .B(DP_pipe03[18]), .ZN(
        DP_mult_209_n1762) );
  XNOR2_X1 DP_mult_209_U2010 ( .A(DP_mult_209_n2252), .B(DP_pipe03[12]), .ZN(
        DP_mult_209_n1768) );
  XNOR2_X1 DP_mult_209_U2009 ( .A(DP_mult_209_n2252), .B(DP_pipe03[10]), .ZN(
        DP_mult_209_n1770) );
  XNOR2_X1 DP_mult_209_U2008 ( .A(DP_mult_209_n2252), .B(DP_pipe03[14]), .ZN(
        DP_mult_209_n1766) );
  XNOR2_X1 DP_mult_209_U2007 ( .A(DP_mult_209_n2252), .B(DP_pipe03[8]), .ZN(
        DP_mult_209_n1772) );
  XNOR2_X1 DP_mult_209_U2006 ( .A(DP_mult_209_n2252), .B(DP_pipe03[2]), .ZN(
        DP_mult_209_n1778) );
  XNOR2_X1 DP_mult_209_U2005 ( .A(DP_mult_209_n2304), .B(DP_pipe03[0]), .ZN(
        DP_mult_209_n1505) );
  INV_X1 DP_mult_209_U2004 ( .A(DP_mult_209_n1482), .ZN(DP_mult_209_n2317) );
  OAI21_X1 DP_mult_209_U2003 ( .B1(DP_mult_209_n2205), .B2(DP_mult_209_n2185), 
        .A(DP_mult_209_n2317), .ZN(DP_mult_209_n1194) );
  INV_X1 DP_mult_209_U2002 ( .A(DP_mult_209_n1582), .ZN(DP_mult_209_n2313) );
  INV_X1 DP_mult_209_U2001 ( .A(DP_mult_209_n1732), .ZN(DP_mult_209_n2307) );
  INV_X1 DP_mult_209_U2000 ( .A(DP_mult_209_n1657), .ZN(DP_mult_209_n2310) );
  OAI22_X1 DP_mult_209_U1999 ( .A1(DP_mult_209_n2225), .A2(DP_mult_209_n1758), 
        .B1(DP_mult_209_n1757), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1459)
         );
  INV_X1 DP_mult_209_U1998 ( .A(DP_mult_209_n1607), .ZN(DP_mult_209_n2312) );
  OAI21_X1 DP_mult_209_U1997 ( .B1(DP_mult_209_n1961), .B2(DP_mult_209_n2061), 
        .A(DP_mult_209_n2312), .ZN(DP_mult_209_n1314) );
  INV_X1 DP_mult_209_U1996 ( .A(DP_mult_209_n1557), .ZN(DP_mult_209_n2314) );
  NOR2_X1 DP_mult_209_U1995 ( .A1(DP_mult_209_n2230), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1289) );
  NOR2_X1 DP_mult_209_U1994 ( .A1(DP_mult_209_n2237), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1337) );
  OAI22_X1 DP_mult_209_U1993 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1765), 
        .B1(DP_mult_209_n1764), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1466)
         );
  NOR2_X1 DP_mult_209_U1992 ( .A1(DP_mult_209_n2229), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1265) );
  INV_X1 DP_mult_209_U1991 ( .A(DP_mult_209_n802), .ZN(DP_mult_209_n803) );
  INV_X1 DP_mult_209_U1990 ( .A(DP_mult_209_n1707), .ZN(DP_mult_209_n2308) );
  OAI22_X1 DP_mult_209_U1989 ( .A1(DP_mult_209_n2225), .A2(DP_mult_209_n1766), 
        .B1(DP_mult_209_n1765), .B2(DP_mult_209_n2249), .ZN(DP_mult_209_n1467)
         );
  NOR2_X1 DP_mult_209_U1988 ( .A1(DP_mult_209_n2228), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1241) );
  NOR2_X1 DP_mult_209_U1987 ( .A1(DP_mult_209_n2240), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1361) );
  OAI22_X1 DP_mult_209_U1986 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1771), 
        .B1(DP_mult_209_n1770), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1472)
         );
  OAI22_X1 DP_mult_209_U1985 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1759), 
        .B1(DP_mult_209_n1758), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1460)
         );
  INV_X1 DP_mult_209_U1984 ( .A(DP_mult_209_n1682), .ZN(DP_mult_209_n2309) );
  OAI22_X1 DP_mult_209_U1983 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1772), 
        .B1(DP_mult_209_n1771), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1473)
         );
  OAI22_X1 DP_mult_209_U1982 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1774), 
        .B1(DP_mult_209_n1773), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1475)
         );
  OAI21_X1 DP_mult_209_U1981 ( .B1(DP_mult_209_n2244), .B2(DP_mult_209_n2218), 
        .A(DP_mult_209_n2310), .ZN(DP_mult_209_n1362) );
  OAI22_X1 DP_mult_209_U1980 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1775), 
        .B1(DP_mult_209_n1774), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1476)
         );
  OAI22_X1 DP_mult_209_U1979 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1769), 
        .B1(DP_mult_209_n1768), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1470)
         );
  NOR2_X1 DP_mult_209_U1978 ( .A1(DP_mult_209_n2234), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1313) );
  NOR2_X1 DP_mult_209_U1977 ( .A1(DP_mult_209_n2045), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1217) );
  OAI22_X1 DP_mult_209_U1976 ( .A1(DP_mult_209_n2225), .A2(DP_mult_209_n1761), 
        .B1(DP_mult_209_n1760), .B2(DP_mult_209_n2249), .ZN(DP_mult_209_n1462)
         );
  OAI22_X1 DP_mult_209_U1975 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1767), 
        .B1(DP_mult_209_n1766), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1468)
         );
  OAI22_X1 DP_mult_209_U1974 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1777), 
        .B1(DP_mult_209_n1776), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1478)
         );
  INV_X1 DP_mult_209_U1973 ( .A(DP_mult_209_n1632), .ZN(DP_mult_209_n2311) );
  INV_X1 DP_mult_209_U1972 ( .A(DP_mult_209_n724), .ZN(DP_mult_209_n725) );
  NOR2_X1 DP_mult_209_U1971 ( .A1(DP_mult_209_n1181), .A2(DP_mult_209_n1192), 
        .ZN(DP_mult_209_n644) );
  NAND2_X1 DP_mult_209_U1970 ( .A1(DP_mult_209_n1181), .A2(DP_mult_209_n1192), 
        .ZN(DP_mult_209_n645) );
  NAND2_X1 DP_mult_209_U1969 ( .A1(DP_mult_209_n2294), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1556) );
  NAND2_X1 DP_mult_209_U1968 ( .A1(DP_mult_209_n2291), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1581) );
  NAND2_X1 DP_mult_209_U1967 ( .A1(DP_mult_209_n2286), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1606) );
  NAND2_X1 DP_mult_209_U1966 ( .A1(DP_mult_209_n2272), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1681) );
  NAND2_X1 DP_mult_209_U1965 ( .A1(DP_mult_209_n2267), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1706) );
  NAND2_X1 DP_mult_209_U1964 ( .A1(DP_mult_209_n2304), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1506) );
  NAND2_X1 DP_mult_209_U1963 ( .A1(DP_mult_209_n2276), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1656) );
  NAND2_X1 DP_mult_209_U1962 ( .A1(DP_mult_209_n2280), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1631) );
  AOI21_X1 DP_mult_209_U1961 ( .B1(DP_mult_209_n1970), .B2(DP_mult_209_n1969), 
        .A(DP_mult_209_n1976), .ZN(DP_mult_209_n646) );
  NAND2_X1 DP_mult_209_U1960 ( .A1(DP_mult_209_n2299), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1531) );
  NAND2_X1 DP_mult_209_U1959 ( .A1(DP_mult_209_n2252), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1781) );
  NOR2_X1 DP_mult_209_U1958 ( .A1(DP_mult_209_n1958), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1433) );
  NOR2_X1 DP_mult_209_U1957 ( .A1(DP_mult_209_n2245), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1409) );
  INV_X1 DP_mult_209_U1956 ( .A(DP_mult_209_n2186), .ZN(DP_mult_209_n2227) );
  INV_X1 DP_mult_209_U1955 ( .A(DP_mult_209_n1994), .ZN(DP_mult_209_n2240) );
  INV_X1 DP_mult_209_U1954 ( .A(DP_mult_209_n1961), .ZN(DP_mult_209_n2237) );
  INV_X1 DP_mult_209_U1953 ( .A(DP_mult_209_n2077), .ZN(DP_mult_209_n2215) );
  INV_X1 DP_mult_209_U1952 ( .A(DP_mult_209_n2061), .ZN(DP_mult_209_n2214) );
  NOR2_X1 DP_mult_209_U1951 ( .A1(DP_mult_209_n2243), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1385) );
  INV_X1 DP_mult_209_U1950 ( .A(DP_mult_209_n1532), .ZN(DP_mult_209_n2315) );
  INV_X1 DP_mult_209_U1949 ( .A(DP_mult_209_n682), .ZN(DP_mult_209_n683) );
  NAND2_X1 DP_mult_209_U1948 ( .A1(DP_mult_209_n2262), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1731) );
  INV_X1 DP_mult_209_U1947 ( .A(DP_mult_209_n1507), .ZN(DP_mult_209_n2316) );
  OAI21_X1 DP_mult_209_U1946 ( .B1(DP_mult_209_n2087), .B2(DP_mult_209_n2016), 
        .A(DP_mult_209_n2316), .ZN(DP_mult_209_n1218) );
  OAI22_X1 DP_mult_209_U1945 ( .A1(DP_mult_209_n2225), .A2(DP_mult_209_n1770), 
        .B1(DP_mult_209_n1769), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1471)
         );
  OAI22_X1 DP_mult_209_U1944 ( .A1(DP_mult_209_n2225), .A2(DP_mult_209_n1763), 
        .B1(DP_mult_209_n1762), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1464)
         );
  OAI22_X1 DP_mult_209_U1943 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1773), 
        .B1(DP_mult_209_n1772), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1474)
         );
  OAI22_X1 DP_mult_209_U1942 ( .A1(DP_mult_209_n2225), .A2(DP_mult_209_n1762), 
        .B1(DP_mult_209_n1761), .B2(DP_mult_209_n2249), .ZN(DP_mult_209_n1463)
         );
  OAI22_X1 DP_mult_209_U1941 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1768), 
        .B1(DP_mult_209_n1767), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1469)
         );
  OAI22_X1 DP_mult_209_U1940 ( .A1(DP_mult_209_n2225), .A2(DP_mult_209_n1760), 
        .B1(DP_mult_209_n1759), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1461)
         );
  OAI22_X1 DP_mult_209_U1939 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1764), 
        .B1(DP_mult_209_n1763), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1465)
         );
  NOR2_X1 DP_mult_209_U1938 ( .A1(DP_mult_209_n2248), .A2(DP_mult_209_n1997), 
        .ZN(DP_mult_209_n1457) );
  INV_X1 DP_mult_209_U1937 ( .A(DP_mult_209_n2296), .ZN(DP_mult_209_n2294) );
  INV_X1 DP_mult_209_U1936 ( .A(DP_mult_209_n2289), .ZN(DP_mult_209_n2286) );
  OAI22_X1 DP_mult_209_U1935 ( .A1(DP_mult_209_n2224), .A2(DP_mult_209_n1779), 
        .B1(DP_mult_209_n1778), .B2(DP_mult_209_n2250), .ZN(DP_mult_209_n1480)
         );
  NAND2_X1 DP_mult_209_U1934 ( .A1(DP_mult_209_n1941), .A2(DP_mult_209_n1996), 
        .ZN(DP_mult_209_n1756) );
  OR2_X1 DP_mult_209_U1933 ( .A1(DP_mult_209_n1194), .A2(DP_mult_209_n676), 
        .ZN(DP_mult_209_n2182) );
  NAND2_X1 DP_mult_209_U1932 ( .A1(DP_mult_209_n678), .A2(DP_mult_209_n677), 
        .ZN(DP_mult_209_n335) );
  NAND2_X1 DP_mult_209_U1931 ( .A1(DP_mult_209_n1159), .A2(DP_mult_209_n1161), 
        .ZN(DP_mult_209_n627) );
  NOR2_X1 DP_mult_209_U1930 ( .A1(DP_mult_209_n1171), .A2(DP_mult_209_n1174), 
        .ZN(DP_mult_209_n633) );
  NAND2_X1 DP_mult_209_U1929 ( .A1(DP_mult_209_n1175), .A2(DP_mult_209_n1178), 
        .ZN(DP_mult_209_n637) );
  NAND2_X1 DP_mult_209_U1928 ( .A1(DP_mult_209_n679), .A2(DP_mult_209_n680), 
        .ZN(DP_mult_209_n341) );
  NAND2_X1 DP_mult_209_U1927 ( .A1(DP_mult_209_n681), .A2(DP_mult_209_n684), 
        .ZN(DP_mult_209_n352) );
  NAND2_X1 DP_mult_209_U1926 ( .A1(DP_mult_209_n685), .A2(DP_mult_209_n688), 
        .ZN(DP_mult_209_n369) );
  NOR2_X1 DP_mult_209_U1925 ( .A1(DP_mult_209_n1159), .A2(DP_mult_209_n1161), 
        .ZN(DP_mult_209_n626) );
  OR2_X1 DP_mult_209_U1924 ( .A1(DP_mult_209_n679), .A2(DP_mult_209_n680), 
        .ZN(DP_mult_209_n2181) );
  OR2_X1 DP_mult_209_U1923 ( .A1(DP_mult_209_n681), .A2(DP_mult_209_n684), 
        .ZN(DP_mult_209_n2180) );
  NOR2_X1 DP_mult_209_U1922 ( .A1(DP_mult_209_n678), .A2(DP_mult_209_n677), 
        .ZN(DP_mult_209_n334) );
  NOR2_X1 DP_mult_209_U1921 ( .A1(DP_mult_209_n1165), .A2(DP_mult_209_n1170), 
        .ZN(DP_mult_209_n631) );
  NOR2_X1 DP_mult_209_U1920 ( .A1(DP_mult_209_n1175), .A2(DP_mult_209_n1178), 
        .ZN(DP_mult_209_n636) );
  OR2_X1 DP_mult_209_U1919 ( .A1(DP_mult_209_n685), .A2(DP_mult_209_n688), 
        .ZN(DP_mult_209_n2179) );
  OAI21_X1 DP_mult_209_U1918 ( .B1(DP_mult_209_n646), .B2(DP_mult_209_n644), 
        .A(DP_mult_209_n645), .ZN(DP_mult_209_n643) );
  AOI21_X1 DP_mult_209_U1917 ( .B1(DP_mult_209_n643), .B2(DP_mult_209_n1971), 
        .A(DP_mult_209_n1977), .ZN(DP_mult_209_n638) );
  AND2_X1 DP_mult_209_U1916 ( .A1(DP_mult_209_n1194), .A2(DP_mult_209_n676), 
        .ZN(DP_mult_209_n2178) );
  INV_X1 DP_mult_209_U1915 ( .A(DP_mult_209_n676), .ZN(DP_mult_209_n677) );
  NAND2_X1 DP_mult_209_U1914 ( .A1(DP_mult_209_n2179), .A2(DP_mult_209_n369), 
        .ZN(DP_mult_209_n304) );
  NAND2_X1 DP_mult_209_U1913 ( .A1(DP_mult_209_n2180), .A2(DP_mult_209_n352), 
        .ZN(DP_mult_209_n303) );
  NAND2_X1 DP_mult_209_U1912 ( .A1(DP_mult_209_n2181), .A2(DP_mult_209_n341), 
        .ZN(DP_mult_209_n302) );
  NAND2_X1 DP_mult_209_U1911 ( .A1(DP_mult_209_n2159), .A2(DP_mult_209_n2175), 
        .ZN(DP_mult_209_n610) );
  NOR2_X1 DP_mult_209_U1910 ( .A1(DP_mult_209_n1085), .A2(DP_mult_209_n1098), 
        .ZN(DP_mult_209_n592) );
  NAND2_X1 DP_mult_209_U1909 ( .A1(DP_mult_209_n1085), .A2(DP_mult_209_n1098), 
        .ZN(DP_mult_209_n593) );
  NAND2_X1 DP_mult_209_U1908 ( .A1(DP_mult_209_n1099), .A2(DP_mult_209_n1110), 
        .ZN(DP_mult_209_n598) );
  INV_X1 DP_mult_209_U1907 ( .A(DP_mult_209_n369), .ZN(DP_mult_209_n367) );
  OR2_X1 DP_mult_209_U1906 ( .A1(DP_mult_209_n694), .A2(DP_mult_209_n689), 
        .ZN(DP_mult_209_n2177) );
  NAND2_X1 DP_mult_209_U1905 ( .A1(DP_mult_209_n695), .A2(DP_mult_209_n700), 
        .ZN(DP_mult_209_n387) );
  OR2_X1 DP_mult_209_U1904 ( .A1(DP_mult_209_n1111), .A2(DP_mult_209_n1122), 
        .ZN(DP_mult_209_n2176) );
  OR2_X1 DP_mult_209_U1903 ( .A1(DP_mult_209_n1133), .A2(DP_mult_209_n1142), 
        .ZN(DP_mult_209_n2175) );
  AOI21_X1 DP_mult_209_U1902 ( .B1(DP_mult_209_n2176), .B2(DP_mult_209_n1973), 
        .A(DP_mult_209_n1980), .ZN(DP_mult_209_n600) );
  NOR2_X1 DP_mult_209_U1901 ( .A1(DP_mult_209_n1099), .A2(DP_mult_209_n1110), 
        .ZN(DP_mult_209_n597) );
  AOI21_X1 DP_mult_209_U1900 ( .B1(DP_mult_209_n376), .B2(DP_mult_209_n2179), 
        .A(DP_mult_209_n367), .ZN(DP_mult_209_n365) );
  AOI21_X1 DP_mult_209_U1899 ( .B1(DP_mult_209_n362), .B2(DP_mult_209_n394), 
        .A(DP_mult_209_n363), .ZN(DP_mult_209_n361) );
  OAI21_X1 DP_mult_209_U1898 ( .B1(DP_mult_209_n405), .B2(DP_mult_209_n360), 
        .A(DP_mult_209_n361), .ZN(DP_mult_209_n359) );
  AOI21_X1 DP_mult_209_U1897 ( .B1(DP_mult_209_n2175), .B2(DP_mult_209_n1972), 
        .A(DP_mult_209_n1979), .ZN(DP_mult_209_n611) );
  OR2_X1 DP_mult_209_U1896 ( .A1(DP_mult_209_n1123), .A2(DP_mult_209_n1132), 
        .ZN(DP_mult_209_n2174) );
  OAI21_X1 DP_mult_209_U1895 ( .B1(DP_mult_209_n628), .B2(DP_mult_209_n626), 
        .A(DP_mult_209_n627), .ZN(DP_mult_209_n625) );
  AOI21_X1 DP_mult_209_U1894 ( .B1(DP_mult_209_n625), .B2(DP_mult_209_n1982), 
        .A(DP_mult_209_n1974), .ZN(DP_mult_209_n620) );
  OR2_X1 DP_mult_209_U1893 ( .A1(DP_mult_209_n709), .A2(DP_mult_209_n716), 
        .ZN(DP_mult_209_n2173) );
  INV_X1 DP_mult_209_U1892 ( .A(DP_mult_209_n341), .ZN(DP_mult_209_n339) );
  OR2_X1 DP_mult_209_U1891 ( .A1(DP_mult_209_n717), .A2(DP_mult_209_n726), 
        .ZN(DP_mult_209_n2172) );
  OR2_X1 DP_mult_209_U1890 ( .A1(DP_mult_209_n701), .A2(DP_mult_209_n708), 
        .ZN(DP_mult_209_n2171) );
  NOR2_X1 DP_mult_209_U1889 ( .A1(DP_mult_209_n695), .A2(DP_mult_209_n700), 
        .ZN(DP_mult_209_n384) );
  INV_X1 DP_mult_209_U1888 ( .A(DP_mult_209_n352), .ZN(DP_mult_209_n350) );
  OAI21_X1 DP_mult_209_U1887 ( .B1(DP_mult_209_n638), .B2(DP_mult_209_n636), 
        .A(DP_mult_209_n637), .ZN(DP_mult_209_n635) );
  INV_X1 DP_mult_209_U1886 ( .A(DP_mult_209_n384), .ZN(DP_mult_209_n657) );
  NAND2_X1 DP_mult_209_U1885 ( .A1(DP_mult_209_n657), .A2(DP_mult_209_n387), 
        .ZN(DP_mult_209_n306) );
  NAND2_X1 DP_mult_209_U1884 ( .A1(DP_mult_209_n661), .A2(DP_mult_209_n429), 
        .ZN(DP_mult_209_n310) );
  NAND2_X1 DP_mult_209_U1883 ( .A1(DP_mult_209_n2171), .A2(DP_mult_209_n396), 
        .ZN(DP_mult_209_n307) );
  NAND2_X1 DP_mult_209_U1882 ( .A1(DP_mult_209_n2173), .A2(DP_mult_209_n409), 
        .ZN(DP_mult_209_n308) );
  OR2_X1 DP_mult_209_U1881 ( .A1(DP_mult_209_n1039), .A2(DP_mult_209_n1054), 
        .ZN(DP_mult_209_n2170) );
  OR2_X1 DP_mult_209_U1880 ( .A1(DP_mult_209_n1021), .A2(DP_mult_209_n1038), 
        .ZN(DP_mult_209_n2169) );
  NAND2_X1 DP_mult_209_U1879 ( .A1(DP_mult_209_n400), .A2(DP_mult_209_n2171), 
        .ZN(DP_mult_209_n389) );
  NOR2_X1 DP_mult_209_U1878 ( .A1(DP_mult_209_n389), .A2(DP_mult_209_n384), 
        .ZN(DP_mult_209_n382) );
  INV_X1 DP_mult_209_U1877 ( .A(DP_mult_209_n378), .ZN(DP_mult_209_n376) );
  INV_X1 DP_mult_209_U1876 ( .A(DP_mult_209_n418), .ZN(DP_mult_209_n416) );
  NOR2_X1 DP_mult_209_U1875 ( .A1(DP_mult_209_n1003), .A2(DP_mult_209_n1020), 
        .ZN(DP_mult_209_n569) );
  INV_X1 DP_mult_209_U1874 ( .A(DP_mult_209_n396), .ZN(DP_mult_209_n394) );
  NOR2_X1 DP_mult_209_U1873 ( .A1(DP_mult_209_n597), .A2(DP_mult_209_n599), 
        .ZN(DP_mult_209_n595) );
  OAI21_X1 DP_mult_209_U1872 ( .B1(DP_mult_209_n620), .B2(DP_mult_209_n610), 
        .A(DP_mult_209_n611), .ZN(DP_mult_209_n609) );
  NAND2_X1 DP_mult_209_U1871 ( .A1(DP_mult_209_n362), .A2(DP_mult_209_n2171), 
        .ZN(DP_mult_209_n360) );
  OR2_X1 DP_mult_209_U1870 ( .A1(DP_mult_209_n761), .A2(DP_mult_209_n774), 
        .ZN(DP_mult_209_n2167) );
  NOR2_X1 DP_mult_209_U1869 ( .A1(DP_mult_209_n983), .A2(DP_mult_209_n1002), 
        .ZN(DP_mult_209_n563) );
  NOR2_X1 DP_mult_209_U1868 ( .A1(DP_mult_209_n1071), .A2(DP_mult_209_n1084), 
        .ZN(DP_mult_209_n590) );
  NAND2_X1 DP_mult_209_U1867 ( .A1(DP_mult_209_n737), .A2(DP_mult_209_n748), 
        .ZN(DP_mult_209_n436) );
  NAND2_X1 DP_mult_209_U1866 ( .A1(DP_mult_209_n789), .A2(DP_mult_209_n804), 
        .ZN(DP_mult_209_n481) );
  NAND2_X1 DP_mult_209_U1865 ( .A1(DP_mult_209_n2172), .A2(DP_mult_209_n2173), 
        .ZN(DP_mult_209_n402) );
  AOI21_X1 DP_mult_209_U1864 ( .B1(DP_mult_209_n423), .B2(DP_mult_209_n356), 
        .A(DP_mult_209_n359), .ZN(DP_mult_209_n355) );
  NAND2_X1 DP_mult_209_U1863 ( .A1(DP_mult_209_n422), .A2(DP_mult_209_n356), 
        .ZN(DP_mult_209_n354) );
  AND2_X1 DP_mult_209_U1862 ( .A1(DP_mult_209_n1039), .A2(DP_mult_209_n1054), 
        .ZN(DP_mult_209_n2165) );
  NOR2_X1 DP_mult_209_U1861 ( .A1(DP_mult_209_n821), .A2(DP_mult_209_n838), 
        .ZN(DP_mult_209_n502) );
  AOI21_X1 DP_mult_209_U1860 ( .B1(DP_mult_209_n426), .B2(DP_mult_209_n445), 
        .A(DP_mult_209_n427), .ZN(DP_mult_209_n421) );
  INV_X1 DP_mult_209_U1859 ( .A(DP_mult_209_n409), .ZN(DP_mult_209_n407) );
  AOI21_X1 DP_mult_209_U1858 ( .B1(DP_mult_209_n2173), .B2(DP_mult_209_n416), 
        .A(DP_mult_209_n407), .ZN(DP_mult_209_n405) );
  NOR2_X1 DP_mult_209_U1857 ( .A1(DP_mult_209_n805), .A2(DP_mult_209_n820), 
        .ZN(DP_mult_209_n495) );
  NOR2_X1 DP_mult_209_U1856 ( .A1(DP_mult_209_n435), .A2(DP_mult_209_n428), 
        .ZN(DP_mult_209_n426) );
  NOR2_X1 DP_mult_209_U1855 ( .A1(DP_mult_209_n384), .A2(DP_mult_209_n364), 
        .ZN(DP_mult_209_n362) );
  NAND2_X1 DP_mult_209_U1854 ( .A1(DP_mult_209_n662), .A2(DP_mult_209_n436), 
        .ZN(DP_mult_209_n311) );
  NAND2_X1 DP_mult_209_U1853 ( .A1(DP_mult_209_n2166), .A2(DP_mult_209_n2167), 
        .ZN(DP_mult_209_n456) );
  INV_X1 DP_mult_209_U1852 ( .A(DP_mult_209_n563), .ZN(DP_mult_209_n561) );
  INV_X1 DP_mult_209_U1851 ( .A(DP_mult_209_n564), .ZN(DP_mult_209_n562) );
  NAND2_X1 DP_mult_209_U1850 ( .A1(DP_mult_209_n663), .A2(DP_mult_209_n439), 
        .ZN(DP_mult_209_n312) );
  NAND2_X1 DP_mult_209_U1849 ( .A1(DP_mult_209_n426), .A2(DP_mult_209_n663), 
        .ZN(DP_mult_209_n420) );
  INV_X1 DP_mult_209_U1848 ( .A(DP_mult_209_n502), .ZN(DP_mult_209_n668) );
  OAI21_X1 DP_mult_209_U1847 ( .B1(DP_mult_209_n421), .B2(DP_mult_209_n402), 
        .A(DP_mult_209_n405), .ZN(DP_mult_209_n401) );
  INV_X1 DP_mult_209_U1846 ( .A(DP_mult_209_n439), .ZN(DP_mult_209_n445) );
  INV_X1 DP_mult_209_U1845 ( .A(DP_mult_209_n438), .ZN(DP_mult_209_n663) );
  INV_X1 DP_mult_209_U1844 ( .A(DP_mult_209_n436), .ZN(DP_mult_209_n434) );
  AOI21_X1 DP_mult_209_U1843 ( .B1(DP_mult_209_n662), .B2(DP_mult_209_n445), 
        .A(DP_mult_209_n434), .ZN(DP_mult_209_n432) );
  NAND2_X1 DP_mult_209_U1842 ( .A1(DP_mult_209_n663), .A2(DP_mult_209_n662), 
        .ZN(DP_mult_209_n431) );
  INV_X1 DP_mult_209_U1841 ( .A(DP_mult_209_n503), .ZN(DP_mult_209_n501) );
  INV_X1 DP_mult_209_U1840 ( .A(DP_mult_209_n481), .ZN(DP_mult_209_n483) );
  OAI21_X1 DP_mult_209_U1839 ( .B1(DP_mult_209_n492), .B2(DP_mult_209_n467), 
        .A(DP_mult_209_n468), .ZN(DP_mult_209_n466) );
  INV_X1 DP_mult_209_U1838 ( .A(DP_mult_209_n461), .ZN(DP_mult_209_n459) );
  INV_X1 DP_mult_209_U1837 ( .A(DP_mult_209_n435), .ZN(DP_mult_209_n662) );
  NOR2_X1 DP_mult_209_U1836 ( .A1(DP_mult_209_n402), .A2(DP_mult_209_n360), 
        .ZN(DP_mult_209_n356) );
  OAI21_X1 DP_mult_209_U1835 ( .B1(DP_mult_209_n531), .B2(DP_mult_209_n535), 
        .A(DP_mult_209_n532), .ZN(DP_mult_209_n526) );
  NOR2_X1 DP_mult_209_U1834 ( .A1(DP_mult_209_n420), .A2(DP_mult_209_n402), 
        .ZN(DP_mult_209_n400) );
  NAND2_X1 DP_mult_209_U1833 ( .A1(DP_mult_209_n2004), .A2(DP_mult_209_n668), 
        .ZN(DP_mult_209_n498) );
  INV_X1 DP_mult_209_U1832 ( .A(DP_mult_209_n420), .ZN(DP_mult_209_n422) );
  NOR2_X1 DP_mult_209_U1831 ( .A1(DP_mult_209_n2119), .A2(DP_mult_209_n467), 
        .ZN(DP_mult_209_n465) );
  INV_X1 DP_mult_209_U1830 ( .A(DP_mult_209_n400), .ZN(DP_mult_209_n398) );
  NOR2_X1 DP_mult_209_U1829 ( .A1(DP_mult_209_n2123), .A2(DP_mult_209_n451), 
        .ZN(DP_mult_209_n301) );
  NAND2_X1 DP_mult_209_U1828 ( .A1(DP_mult_209_n465), .A2(DP_mult_209_n2004), 
        .ZN(DP_mult_209_n463) );
  NOR2_X1 DP_mult_209_U1827 ( .A1(DP_mult_209_n451), .A2(DP_mult_209_n2164), 
        .ZN(DP_mult_209_n2162) );
  NOR2_X1 DP_mult_209_U1826 ( .A1(DP_mult_209_n2123), .A2(DP_mult_209_n451), 
        .ZN(DP_mult_209_n2163) );
  INV_X1 DP_mult_209_U1825 ( .A(DP_mult_209_n2077), .ZN(DP_mult_209_n2160) );
  INV_X2 DP_mult_209_U1824 ( .A(DP_mult_209_n2062), .ZN(DP_mult_209_n2213) );
  INV_X2 DP_mult_209_U1823 ( .A(DP_mult_209_n2305), .ZN(DP_mult_209_n2304) );
  OR2_X1 DP_mult_209_U1822 ( .A1(DP_mult_209_n1143), .A2(DP_mult_209_n1150), 
        .ZN(DP_mult_209_n2159) );
  INV_X2 DP_mult_209_U1821 ( .A(DP_mult_209_n2274), .ZN(DP_mult_209_n2271) );
  INV_X1 DP_mult_209_U1820 ( .A(DP_mult_209_n1975), .ZN(DP_mult_209_n2157) );
  INV_X2 DP_mult_209_U1819 ( .A(DP_mult_209_n2270), .ZN(DP_mult_209_n2267) );
  INV_X2 DP_mult_209_U1818 ( .A(DP_mult_209_n2265), .ZN(DP_mult_209_n2262) );
  INV_X1 DP_mult_209_U1817 ( .A(DP_mult_209_n2153), .ZN(DP_mult_209_n2212) );
  NOR2_X1 DP_mult_209_U1816 ( .A1(DP_mult_209_n805), .A2(DP_mult_209_n820), 
        .ZN(DP_mult_209_n2154) );
  BUF_X2 DP_mult_209_U1815 ( .A(DP_mult_209_n279), .Z(DP_mult_209_n2193) );
  INV_X2 DP_mult_209_U1814 ( .A(DP_mult_209_n2232), .ZN(DP_mult_209_n2230) );
  BUF_X2 DP_mult_209_U1813 ( .A(DP_mult_209_n2003), .Z(DP_mult_209_n2196) );
  INV_X1 DP_mult_209_U1812 ( .A(DP_mult_209_n2122), .ZN(DP_mult_209_n2151) );
  OR2_X1 DP_mult_209_U1811 ( .A1(DP_mult_209_n2068), .A2(DP_mult_209_n534), 
        .ZN(DP_mult_209_n2150) );
  INV_X2 DP_mult_209_U1810 ( .A(DP_mult_209_n2152), .ZN(DP_mult_209_n2156) );
  AOI21_X1 DP_mult_209_U1809 ( .B1(DP_mult_209_n1957), .B2(DP_mult_209_n567), 
        .A(DP_mult_209_n1948), .ZN(DP_mult_209_n2149) );
  NAND3_X1 DP_mult_209_U1808 ( .A1(DP_mult_209_n2146), .A2(DP_mult_209_n2147), 
        .A3(DP_mult_209_n2148), .ZN(DP_mult_209_n1022) );
  NAND2_X1 DP_mult_209_U1807 ( .A1(DP_mult_209_n1027), .A2(DP_mult_209_n1044), 
        .ZN(DP_mult_209_n2148) );
  NAND2_X1 DP_mult_209_U1806 ( .A1(DP_mult_209_n1042), .A2(DP_mult_209_n1044), 
        .ZN(DP_mult_209_n2147) );
  NAND2_X1 DP_mult_209_U1805 ( .A1(DP_mult_209_n1042), .A2(DP_mult_209_n2026), 
        .ZN(DP_mult_209_n2146) );
  INV_X2 DP_mult_209_U1804 ( .A(DP_mult_209_n2232), .ZN(DP_mult_209_n2231) );
  NOR2_X1 DP_mult_209_U1803 ( .A1(DP_mult_209_n919), .A2(DP_mult_209_n940), 
        .ZN(DP_mult_209_n542) );
  NOR2_X1 DP_mult_209_U1802 ( .A1(DP_mult_209_n919), .A2(DP_mult_209_n940), 
        .ZN(DP_mult_209_n2145) );
  NAND3_X1 DP_mult_209_U1801 ( .A1(DP_mult_209_n2142), .A2(DP_mult_209_n2143), 
        .A3(DP_mult_209_n2144), .ZN(DP_mult_209_n992) );
  NAND2_X1 DP_mult_209_U1800 ( .A1(DP_mult_209_n1394), .A2(DP_mult_209_n1018), 
        .ZN(DP_mult_209_n2144) );
  NAND2_X1 DP_mult_209_U1799 ( .A1(DP_mult_209_n1001), .A2(DP_mult_209_n1018), 
        .ZN(DP_mult_209_n2143) );
  NAND2_X1 DP_mult_209_U1798 ( .A1(DP_mult_209_n1001), .A2(DP_mult_209_n1394), 
        .ZN(DP_mult_209_n2142) );
  XOR2_X1 DP_mult_209_U1797 ( .A(DP_mult_209_n2141), .B(DP_mult_209_n1018), 
        .Z(DP_mult_209_n993) );
  XOR2_X1 DP_mult_209_U1796 ( .A(DP_mult_209_n1001), .B(DP_mult_209_n1394), 
        .Z(DP_mult_209_n2141) );
  NAND3_X1 DP_mult_209_U1795 ( .A1(DP_mult_209_n2138), .A2(DP_mult_209_n2139), 
        .A3(DP_mult_209_n2140), .ZN(DP_mult_209_n1018) );
  NAND2_X1 DP_mult_209_U1794 ( .A1(DP_mult_209_n1351), .A2(DP_mult_209_n1285), 
        .ZN(DP_mult_209_n2140) );
  NAND2_X1 DP_mult_209_U1793 ( .A1(DP_mult_209_n1263), .A2(DP_mult_209_n1285), 
        .ZN(DP_mult_209_n2139) );
  NAND2_X1 DP_mult_209_U1792 ( .A1(DP_mult_209_n1263), .A2(DP_mult_209_n1351), 
        .ZN(DP_mult_209_n2138) );
  OR2_X1 DP_mult_209_U1791 ( .A1(DP_mult_209_n857), .A2(DP_mult_209_n876), 
        .ZN(DP_mult_209_n2137) );
  INV_X1 DP_mult_209_U1790 ( .A(DP_mult_209_n2004), .ZN(DP_mult_209_n2136) );
  NAND3_X1 DP_mult_209_U1789 ( .A1(DP_mult_209_n2133), .A2(DP_mult_209_n2134), 
        .A3(DP_mult_209_n2135), .ZN(DP_mult_209_n954) );
  NAND2_X1 DP_mult_209_U1788 ( .A1(DP_mult_209_n1414), .A2(DP_mult_209_n1282), 
        .ZN(DP_mult_209_n2135) );
  NAND2_X1 DP_mult_209_U1787 ( .A1(DP_mult_209_n1304), .A2(DP_mult_209_n1282), 
        .ZN(DP_mult_209_n2134) );
  NAND2_X1 DP_mult_209_U1786 ( .A1(DP_mult_209_n1414), .A2(DP_mult_209_n1304), 
        .ZN(DP_mult_209_n2133) );
  XOR2_X1 DP_mult_209_U1785 ( .A(DP_mult_209_n2132), .B(DP_mult_209_n2120), 
        .Z(DP_mult_209_n955) );
  XOR2_X1 DP_mult_209_U1784 ( .A(DP_mult_209_n1414), .B(DP_mult_209_n1282), 
        .Z(DP_mult_209_n2132) );
  OAI21_X1 DP_mult_209_U1783 ( .B1(DP_mult_209_n2068), .B2(DP_mult_209_n535), 
        .A(DP_mult_209_n532), .ZN(DP_mult_209_n2131) );
  INV_X2 DP_mult_209_U1782 ( .A(DP_mult_209_n2152), .ZN(DP_mult_209_n2211) );
  INV_X2 DP_mult_209_U1781 ( .A(DP_mult_209_n2265), .ZN(DP_mult_209_n2261) );
  NAND3_X1 DP_mult_209_U1780 ( .A1(DP_mult_209_n2128), .A2(DP_mult_209_n2129), 
        .A3(DP_mult_209_n2130), .ZN(DP_mult_209_n1026) );
  NAND2_X1 DP_mult_209_U1779 ( .A1(DP_mult_209_n1048), .A2(DP_mult_209_n1033), 
        .ZN(DP_mult_209_n2130) );
  NAND2_X1 DP_mult_209_U1778 ( .A1(DP_mult_209_n1031), .A2(DP_mult_209_n1033), 
        .ZN(DP_mult_209_n2129) );
  NAND2_X1 DP_mult_209_U1777 ( .A1(DP_mult_209_n1031), .A2(DP_mult_209_n1048), 
        .ZN(DP_mult_209_n2128) );
  INV_X2 DP_mult_209_U1776 ( .A(DP_mult_209_n2254), .ZN(DP_mult_209_n2251) );
  BUF_X2 DP_mult_209_U1775 ( .A(DP_mult_209_n2003), .Z(DP_mult_209_n2195) );
  NAND3_X1 DP_mult_209_U1774 ( .A1(DP_mult_209_n2125), .A2(DP_mult_209_n2126), 
        .A3(DP_mult_209_n2127), .ZN(DP_mult_209_n918) );
  NAND2_X1 DP_mult_209_U1773 ( .A1(DP_mult_209_n942), .A2(DP_mult_209_n923), 
        .ZN(DP_mult_209_n2127) );
  NAND2_X1 DP_mult_209_U1772 ( .A1(DP_mult_209_n921), .A2(DP_mult_209_n923), 
        .ZN(DP_mult_209_n2126) );
  NAND2_X1 DP_mult_209_U1771 ( .A1(DP_mult_209_n921), .A2(DP_mult_209_n942), 
        .ZN(DP_mult_209_n2125) );
  AND2_X1 DP_mult_209_U1770 ( .A1(DP_mult_209_n537), .A2(DP_mult_209_n2013), 
        .ZN(DP_mult_209_n2164) );
  INV_X1 DP_mult_209_U1769 ( .A(DP_mult_209_n1984), .ZN(DP_mult_209_n2124) );
  AND2_X1 DP_mult_209_U1768 ( .A1(DP_mult_209_n537), .A2(DP_mult_209_n2013), 
        .ZN(DP_mult_209_n2123) );
  BUF_X2 DP_mult_209_U1767 ( .A(DP_mult_209_n2003), .Z(DP_mult_209_n2194) );
  XNOR2_X1 DP_mult_209_U1766 ( .A(DP_coeffs_ff_int[89]), .B(DP_mult_209_n2269), 
        .ZN(DP_mult_209_n1814) );
  OR2_X1 DP_mult_209_U1765 ( .A1(DP_mult_209_n897), .A2(DP_mult_209_n918), 
        .ZN(DP_mult_209_n2122) );
  XNOR2_X1 DP_mult_209_U1764 ( .A(DP_mult_209_n1048), .B(DP_mult_209_n1033), 
        .ZN(DP_mult_209_n2121) );
  XNOR2_X1 DP_mult_209_U1763 ( .A(DP_mult_209_n2121), .B(DP_mult_209_n1031), 
        .ZN(DP_mult_209_n1027) );
  BUF_X1 DP_mult_209_U1762 ( .A(DP_mult_209_n1304), .Z(DP_mult_209_n2120) );
  OR2_X1 DP_mult_209_U1761 ( .A1(DP_mult_209_n495), .A2(DP_mult_209_n502), 
        .ZN(DP_mult_209_n2119) );
  AND2_X1 DP_mult_209_U1760 ( .A1(DP_mult_209_n1810), .A2(DP_mult_209_n2233), 
        .ZN(DP_mult_209_n2152) );
  INV_X2 DP_mult_209_U1759 ( .A(DP_mult_209_n2301), .ZN(DP_mult_209_n2298) );
  NOR2_X1 DP_mult_209_U1758 ( .A1(DP_mult_209_n495), .A2(DP_mult_209_n502), 
        .ZN(DP_mult_209_n489) );
  CLKBUF_X1 DP_mult_209_U1757 ( .A(DP_mult_209_n489), .Z(DP_mult_209_n2118) );
  INV_X1 DP_mult_209_U1756 ( .A(DP_mult_209_n2190), .ZN(DP_mult_209_n2233) );
  INV_X2 DP_mult_209_U1755 ( .A(DP_mult_209_n2187), .ZN(DP_mult_209_n2245) );
  XNOR2_X1 DP_mult_209_U1754 ( .A(DP_coeffs_ff_int[89]), .B(
        DP_coeffs_ff_int[90]), .ZN(DP_mult_209_n2117) );
  INV_X2 DP_mult_209_U1753 ( .A(DP_mult_209_n2082), .ZN(DP_mult_209_n2224) );
  XNOR2_X1 DP_mult_209_U1752 ( .A(DP_mult_209_n1027), .B(DP_mult_209_n1044), 
        .ZN(DP_mult_209_n2115) );
  XNOR2_X1 DP_mult_209_U1751 ( .A(DP_mult_209_n1042), .B(DP_mult_209_n2115), 
        .ZN(DP_mult_209_n1023) );
  INV_X1 DP_mult_209_U1750 ( .A(DP_mult_209_n2150), .ZN(DP_mult_209_n2114) );
  NAND2_X1 DP_mult_209_U1749 ( .A1(DP_mult_209_n2112), .A2(DP_mult_209_n2113), 
        .ZN(DP_mult_209_n1417) );
  OR2_X1 DP_mult_209_U1748 ( .A1(DP_mult_209_n1959), .A2(DP_mult_209_n1714), 
        .ZN(DP_mult_209_n2113) );
  OR2_X1 DP_mult_209_U1747 ( .A1(DP_mult_209_n2193), .A2(DP_mult_209_n1715), 
        .ZN(DP_mult_209_n2112) );
  NAND3_X1 DP_mult_209_U1746 ( .A1(DP_mult_209_n2109), .A2(DP_mult_209_n2110), 
        .A3(DP_mult_209_n2111), .ZN(DP_mult_209_n1014) );
  NAND2_X1 DP_mult_209_U1745 ( .A1(DP_mult_209_n1462), .A2(DP_mult_209_n1395), 
        .ZN(DP_mult_209_n2111) );
  NAND2_X1 DP_mult_209_U1744 ( .A1(DP_mult_209_n1417), .A2(DP_mult_209_n1395), 
        .ZN(DP_mult_209_n2110) );
  NAND2_X1 DP_mult_209_U1743 ( .A1(DP_mult_209_n1417), .A2(DP_mult_209_n1462), 
        .ZN(DP_mult_209_n2109) );
  NAND2_X1 DP_mult_209_U1742 ( .A1(DP_mult_209_n849), .A2(DP_mult_209_n864), 
        .ZN(DP_mult_209_n2107) );
  NAND2_X1 DP_mult_209_U1741 ( .A1(DP_mult_209_n862), .A2(DP_mult_209_n864), 
        .ZN(DP_mult_209_n2106) );
  NAND2_X1 DP_mult_209_U1740 ( .A1(DP_mult_209_n862), .A2(DP_mult_209_n849), 
        .ZN(DP_mult_209_n2105) );
  XOR2_X1 DP_mult_209_U1739 ( .A(DP_mult_209_n862), .B(DP_mult_209_n2104), .Z(
        DP_mult_209_n843) );
  XOR2_X1 DP_mult_209_U1738 ( .A(DP_mult_209_n849), .B(DP_mult_209_n864), .Z(
        DP_mult_209_n2104) );
  INV_X2 DP_mult_209_U1737 ( .A(DP_mult_209_n2184), .ZN(DP_mult_209_n2225) );
  XNOR2_X1 DP_mult_209_U1736 ( .A(DP_mult_209_n942), .B(DP_mult_209_n923), 
        .ZN(DP_mult_209_n2103) );
  XNOR2_X1 DP_mult_209_U1735 ( .A(DP_coeffs_ff_int[73]), .B(DP_mult_209_n1937), 
        .ZN(DP_mult_209_n1806) );
  INV_X1 DP_mult_209_U1734 ( .A(DP_mult_209_n2087), .ZN(DP_mult_209_n2102) );
  OR2_X1 DP_mult_209_U1733 ( .A1(DP_mult_209_n941), .A2(DP_mult_209_n962), 
        .ZN(DP_mult_209_n2100) );
  XNOR2_X1 DP_mult_209_U1732 ( .A(DP_mult_209_n1263), .B(DP_mult_209_n1351), 
        .ZN(DP_mult_209_n2099) );
  XNOR2_X1 DP_mult_209_U1731 ( .A(DP_mult_209_n2099), .B(DP_mult_209_n1285), 
        .ZN(DP_mult_209_n1019) );
  BUF_X2 DP_mult_209_U1730 ( .A(DP_mult_209_n2203), .Z(DP_mult_209_n2191) );
  INV_X2 DP_mult_209_U1729 ( .A(DP_mult_209_n2278), .ZN(DP_mult_209_n2275) );
  XNOR2_X1 DP_mult_209_U1728 ( .A(DP_coeffs_ff_int[93]), .B(DP_mult_209_n2260), 
        .ZN(DP_mult_209_n1816) );
  INV_X2 DP_mult_209_U1727 ( .A(DP_mult_209_n2218), .ZN(DP_mult_209_n2217) );
  INV_X1 DP_mult_209_U1726 ( .A(DP_mult_209_n1960), .ZN(DP_mult_209_n2236) );
  NOR2_X1 DP_mult_209_U1725 ( .A1(DP_mult_209_n941), .A2(DP_mult_209_n962), 
        .ZN(DP_mult_209_n547) );
  INV_X1 DP_mult_209_U1724 ( .A(DP_mult_209_n1989), .ZN(DP_mult_209_n2207) );
  INV_X1 DP_mult_209_U1723 ( .A(DP_mult_209_n1989), .ZN(DP_mult_209_n2096) );
  INV_X1 DP_mult_209_U1722 ( .A(DP_mult_209_n2297), .ZN(DP_mult_209_n2094) );
  INV_X1 DP_mult_209_U1721 ( .A(DP_mult_209_n2297), .ZN(DP_mult_209_n2095) );
  BUF_X1 DP_mult_209_U1720 ( .A(DP_mult_209_n547), .Z(DP_mult_209_n2098) );
  NAND3_X1 DP_mult_209_U1719 ( .A1(DP_mult_209_n2091), .A2(DP_mult_209_n2092), 
        .A3(DP_mult_209_n2093), .ZN(DP_mult_209_n896) );
  NAND2_X1 DP_mult_209_U1718 ( .A1(DP_mult_209_n920), .A2(DP_mult_209_n901), 
        .ZN(DP_mult_209_n2093) );
  NAND2_X1 DP_mult_209_U1717 ( .A1(DP_mult_209_n899), .A2(DP_mult_209_n901), 
        .ZN(DP_mult_209_n2092) );
  NAND2_X1 DP_mult_209_U1716 ( .A1(DP_mult_209_n899), .A2(DP_mult_209_n920), 
        .ZN(DP_mult_209_n2091) );
  OR2_X1 DP_mult_209_U1715 ( .A1(DP_mult_209_n856), .A2(DP_mult_209_n839), 
        .ZN(DP_mult_209_n2090) );
  XNOR2_X1 DP_mult_209_U1714 ( .A(DP_mult_209_n1462), .B(DP_mult_209_n1395), 
        .ZN(DP_mult_209_n2088) );
  XNOR2_X1 DP_mult_209_U1713 ( .A(DP_mult_209_n1417), .B(DP_mult_209_n2088), 
        .ZN(DP_mult_209_n1015) );
  INV_X2 DP_mult_209_U1712 ( .A(DP_mult_209_n2302), .ZN(DP_mult_209_n2299) );
  AND2_X1 DP_mult_209_U1711 ( .A1(DP_mult_209_n1807), .A2(DP_mult_209_n2226), 
        .ZN(DP_mult_209_n2087) );
  NAND3_X1 DP_mult_209_U1710 ( .A1(DP_mult_209_n2083), .A2(DP_mult_209_n2084), 
        .A3(DP_mult_209_n2085), .ZN(DP_mult_209_n946) );
  NAND2_X1 DP_mult_209_U1709 ( .A1(DP_mult_209_n953), .A2(DP_mult_209_n959), 
        .ZN(DP_mult_209_n2085) );
  NAND2_X1 DP_mult_209_U1708 ( .A1(DP_mult_209_n972), .A2(DP_mult_209_n959), 
        .ZN(DP_mult_209_n2084) );
  NAND2_X1 DP_mult_209_U1707 ( .A1(DP_mult_209_n972), .A2(DP_mult_209_n953), 
        .ZN(DP_mult_209_n2083) );
  AND2_X1 DP_mult_209_U1706 ( .A1(DP_mult_209_n1817), .A2(DP_mult_209_n2249), 
        .ZN(DP_mult_209_n2082) );
  NOR2_X1 DP_mult_209_U1705 ( .A1(DP_mult_209_n963), .A2(DP_mult_209_n982), 
        .ZN(DP_mult_209_n558) );
  NOR2_X1 DP_mult_209_U1704 ( .A1(DP_mult_209_n963), .A2(DP_mult_209_n982), 
        .ZN(DP_mult_209_n2081) );
  INV_X1 DP_mult_209_U1703 ( .A(DP_mult_209_n2190), .ZN(DP_mult_209_n2234) );
  NAND2_X1 DP_mult_209_U1702 ( .A1(DP_mult_209_n2079), .A2(DP_mult_209_n2080), 
        .ZN(DP_mult_209_n1356) );
  OR2_X1 DP_mult_209_U1701 ( .A1(DP_mult_209_n1650), .A2(DP_mult_209_n2241), 
        .ZN(DP_mult_209_n2080) );
  OR2_X1 DP_mult_209_U1700 ( .A1(DP_mult_209_n2161), .A2(DP_mult_209_n1651), 
        .ZN(DP_mult_209_n2079) );
  AND2_X2 DP_mult_209_U1699 ( .A1(DP_mult_209_n1812), .A2(DP_mult_209_n2239), 
        .ZN(DP_mult_209_n2078) );
  AND2_X1 DP_mult_209_U1698 ( .A1(DP_mult_209_n1812), .A2(DP_mult_209_n2239), 
        .ZN(DP_mult_209_n2077) );
  INV_X2 DP_mult_209_U1697 ( .A(DP_mult_209_n2065), .ZN(DP_mult_209_n2209) );
  XNOR2_X1 DP_mult_209_U1696 ( .A(DP_mult_209_n953), .B(DP_mult_209_n959), 
        .ZN(DP_mult_209_n2076) );
  XNOR2_X1 DP_mult_209_U1695 ( .A(DP_mult_209_n972), .B(DP_mult_209_n2076), 
        .ZN(DP_mult_209_n947) );
  INV_X2 DP_mult_209_U1694 ( .A(DP_mult_209_n2293), .ZN(DP_mult_209_n2291) );
  NAND3_X1 DP_mult_209_U1693 ( .A1(DP_mult_209_n2073), .A2(DP_mult_209_n2074), 
        .A3(DP_mult_209_n2075), .ZN(DP_mult_209_n1094) );
  NAND2_X1 DP_mult_209_U1692 ( .A1(DP_mult_209_n1400), .A2(DP_mult_209_n1467), 
        .ZN(DP_mult_209_n2075) );
  NAND2_X1 DP_mult_209_U1691 ( .A1(DP_mult_209_n1186), .A2(DP_mult_209_n1467), 
        .ZN(DP_mult_209_n2074) );
  NAND2_X1 DP_mult_209_U1690 ( .A1(DP_mult_209_n1186), .A2(DP_mult_209_n1400), 
        .ZN(DP_mult_209_n2073) );
  INV_X1 DP_mult_209_U1689 ( .A(DP_mult_209_n2288), .ZN(DP_mult_209_n2284) );
  INV_X1 DP_mult_209_U1688 ( .A(DP_mult_209_n2078), .ZN(DP_mult_209_n2161) );
  INV_X1 DP_mult_209_U1687 ( .A(DP_mult_209_n2183), .ZN(DP_mult_209_n2239) );
  INV_X2 DP_mult_209_U1686 ( .A(DP_mult_209_n2244), .ZN(DP_mult_209_n2242) );
  XNOR2_X1 DP_mult_209_U1685 ( .A(DP_coeffs_ff_int[93]), .B(
        DP_coeffs_ff_int[94]), .ZN(DP_mult_209_n2072) );
  NAND3_X1 DP_mult_209_U1684 ( .A1(DP_mult_209_n2069), .A2(DP_mult_209_n2070), 
        .A3(DP_mult_209_n2071), .ZN(DP_mult_209_n940) );
  NAND2_X1 DP_mult_209_U1683 ( .A1(DP_mult_209_n964), .A2(DP_mult_209_n945), 
        .ZN(DP_mult_209_n2071) );
  NAND2_X1 DP_mult_209_U1682 ( .A1(DP_mult_209_n943), .A2(DP_mult_209_n945), 
        .ZN(DP_mult_209_n2070) );
  NAND2_X1 DP_mult_209_U1681 ( .A1(DP_mult_209_n943), .A2(DP_mult_209_n964), 
        .ZN(DP_mult_209_n2069) );
  NOR2_X1 DP_mult_209_U1680 ( .A1(DP_mult_209_n877), .A2(DP_mult_209_n896), 
        .ZN(DP_mult_209_n531) );
  NOR2_X1 DP_mult_209_U1679 ( .A1(DP_mult_209_n877), .A2(DP_mult_209_n896), 
        .ZN(DP_mult_209_n2068) );
  INV_X1 DP_mult_209_U1678 ( .A(DP_mult_209_n2288), .ZN(DP_mult_209_n2285) );
  XNOR2_X1 DP_mult_209_U1677 ( .A(DP_coeffs_ff_int[81]), .B(DP_mult_209_n2288), 
        .ZN(DP_mult_209_n1810) );
  INV_X1 DP_mult_209_U1676 ( .A(DP_mult_209_n2116), .ZN(DP_mult_209_n2185) );
  XNOR2_X1 DP_mult_209_U1675 ( .A(DP_coeffs_ff_int[91]), .B(
        DP_coeffs_ff_int[92]), .ZN(DP_mult_209_n2067) );
  AND2_X1 DP_mult_209_U1674 ( .A1(DP_mult_209_n1809), .A2(DP_mult_209_n267), 
        .ZN(DP_mult_209_n2065) );
  INV_X2 DP_mult_209_U1673 ( .A(DP_mult_209_n2185), .ZN(DP_mult_209_n2064) );
  INV_X1 DP_mult_209_U1672 ( .A(DP_mult_209_n1961), .ZN(DP_mult_209_n2238) );
  INV_X1 DP_mult_209_U1671 ( .A(DP_mult_209_n2186), .ZN(DP_mult_209_n2226) );
  XNOR2_X1 DP_mult_209_U1670 ( .A(DP_coeffs_ff_int[77]), .B(
        DP_coeffs_ff_int[78]), .ZN(DP_mult_209_n2063) );
  XNOR2_X1 DP_mult_209_U1669 ( .A(DP_mult_209_n920), .B(DP_mult_209_n901), 
        .ZN(DP_mult_209_n2060) );
  XNOR2_X1 DP_mult_209_U1668 ( .A(DP_mult_209_n899), .B(DP_mult_209_n2060), 
        .ZN(DP_mult_209_n897) );
  INV_X1 DP_mult_209_U1667 ( .A(DP_mult_209_n1975), .ZN(DP_mult_209_n2219) );
  NOR2_X1 DP_mult_209_U1666 ( .A1(DP_mult_209_n839), .A2(DP_mult_209_n856), 
        .ZN(DP_mult_209_n2059) );
  XNOR2_X1 DP_mult_209_U1665 ( .A(DP_coeffs_ff_int[75]), .B(DP_mult_209_n2301), 
        .ZN(DP_mult_209_n1807) );
  XOR2_X1 DP_mult_209_U1664 ( .A(DP_coeffs_ff_int[76]), .B(
        DP_coeffs_ff_int[75]), .Z(DP_mult_209_n2186) );
  INV_X1 DP_mult_209_U1663 ( .A(DP_mult_209_n2293), .ZN(DP_mult_209_n2290) );
  INV_X1 DP_mult_209_U1662 ( .A(DP_mult_209_n2292), .ZN(DP_mult_209_n2058) );
  XNOR2_X1 DP_mult_209_U1661 ( .A(DP_coeffs_ff_int[87]), .B(DP_mult_209_n2274), 
        .ZN(DP_mult_209_n1813) );
  NOR2_X1 DP_mult_209_U1660 ( .A1(DP_mult_209_n513), .A2(DP_mult_209_n520), 
        .ZN(DP_mult_209_n511) );
  NOR2_X1 DP_mult_209_U1659 ( .A1(DP_mult_209_n520), .A2(DP_mult_209_n513), 
        .ZN(DP_mult_209_n2057) );
  NAND3_X1 DP_mult_209_U1658 ( .A1(DP_mult_209_n2054), .A2(DP_mult_209_n2055), 
        .A3(DP_mult_209_n2056), .ZN(DP_mult_209_n856) );
  NAND2_X1 DP_mult_209_U1657 ( .A1(DP_mult_209_n878), .A2(DP_mult_209_n861), 
        .ZN(DP_mult_209_n2056) );
  NAND2_X1 DP_mult_209_U1656 ( .A1(DP_mult_209_n859), .A2(DP_mult_209_n861), 
        .ZN(DP_mult_209_n2055) );
  NAND2_X1 DP_mult_209_U1655 ( .A1(DP_mult_209_n859), .A2(DP_mult_209_n878), 
        .ZN(DP_mult_209_n2054) );
  XNOR2_X1 DP_mult_209_U1654 ( .A(DP_mult_209_n878), .B(DP_mult_209_n861), 
        .ZN(DP_mult_209_n2053) );
  XNOR2_X1 DP_mult_209_U1653 ( .A(DP_mult_209_n859), .B(DP_mult_209_n2053), 
        .ZN(DP_mult_209_n857) );
  NAND3_X1 DP_mult_209_U1652 ( .A1(DP_mult_209_n2049), .A2(DP_mult_209_n2050), 
        .A3(DP_mult_209_n2051), .ZN(DP_mult_209_n862) );
  NAND2_X1 DP_mult_209_U1651 ( .A1(DP_mult_209_n873), .A2(DP_mult_209_n888), 
        .ZN(DP_mult_209_n2051) );
  NAND2_X1 DP_mult_209_U1650 ( .A1(DP_mult_209_n886), .A2(DP_mult_209_n888), 
        .ZN(DP_mult_209_n2050) );
  NAND2_X1 DP_mult_209_U1649 ( .A1(DP_mult_209_n886), .A2(DP_mult_209_n873), 
        .ZN(DP_mult_209_n2049) );
  XOR2_X1 DP_mult_209_U1648 ( .A(DP_mult_209_n886), .B(DP_mult_209_n2048), .Z(
        DP_mult_209_n863) );
  XOR2_X1 DP_mult_209_U1647 ( .A(DP_mult_209_n873), .B(DP_mult_209_n888), .Z(
        DP_mult_209_n2048) );
  INV_X1 DP_mult_209_U1646 ( .A(DP_mult_209_n2117), .ZN(DP_mult_209_n2187) );
  XOR2_X1 DP_mult_209_U1645 ( .A(DP_coeffs_ff_int[81]), .B(
        DP_coeffs_ff_int[82]), .Z(DP_mult_209_n2190) );
  INV_X2 DP_mult_209_U1644 ( .A(DP_mult_209_n2255), .ZN(DP_mult_209_n2252) );
  INV_X1 DP_mult_209_U1643 ( .A(DP_mult_209_n524), .ZN(DP_mult_209_n2047) );
  XNOR2_X1 DP_mult_209_U1642 ( .A(DP_mult_209_n964), .B(DP_mult_209_n945), 
        .ZN(DP_mult_209_n2046) );
  XNOR2_X1 DP_mult_209_U1641 ( .A(DP_mult_209_n943), .B(DP_mult_209_n2046), 
        .ZN(DP_mult_209_n941) );
  XNOR2_X1 DP_mult_209_U1640 ( .A(DP_coeffs_ff_int[77]), .B(DP_mult_209_n2296), 
        .ZN(DP_mult_209_n1808) );
  XNOR2_X1 DP_mult_209_U1639 ( .A(DP_coeffs_ff_int[79]), .B(DP_mult_209_n2292), 
        .ZN(DP_mult_209_n1809) );
  NOR2_X1 DP_mult_209_U1638 ( .A1(DP_mult_209_n558), .A2(DP_mult_209_n563), 
        .ZN(DP_mult_209_n552) );
  NAND2_X1 DP_mult_209_U1637 ( .A1(DP_mult_209_n1813), .A2(DP_mult_209_n259), 
        .ZN(DP_mult_209_n283) );
  XNOR2_X1 DP_mult_209_U1636 ( .A(DP_mult_209_n2103), .B(DP_mult_209_n921), 
        .ZN(DP_mult_209_n919) );
  XNOR2_X1 DP_mult_209_U1635 ( .A(DP_coeffs_ff_int[73]), .B(
        DP_coeffs_ff_int[74]), .ZN(DP_mult_209_n2116) );
  INV_X2 DP_mult_209_U1634 ( .A(DP_mult_209_n2185), .ZN(DP_mult_209_n2045) );
  NAND2_X1 DP_mult_209_U1633 ( .A1(DP_mult_209_n2042), .A2(DP_mult_209_n2043), 
        .ZN(DP_mult_209_n1442) );
  OR2_X1 DP_mult_209_U1632 ( .A1(DP_mult_209_n1740), .A2(DP_mult_209_n2019), 
        .ZN(DP_mult_209_n2043) );
  OR2_X1 DP_mult_209_U1631 ( .A1(DP_mult_209_n2196), .A2(DP_mult_209_n1741), 
        .ZN(DP_mult_209_n2042) );
  NOR2_X1 DP_mult_209_U1630 ( .A1(DP_mult_209_n1003), .A2(DP_mult_209_n1020), 
        .ZN(DP_mult_209_n2041) );
  NAND3_X1 DP_mult_209_U1629 ( .A1(DP_mult_209_n2038), .A2(DP_mult_209_n2039), 
        .A3(DP_mult_209_n2040), .ZN(DP_mult_209_n1064) );
  NAND2_X1 DP_mult_209_U1628 ( .A1(DP_mult_209_n1332), .A2(DP_mult_209_n1354), 
        .ZN(DP_mult_209_n2040) );
  NAND2_X1 DP_mult_209_U1627 ( .A1(DP_mult_209_n1442), .A2(DP_mult_209_n1354), 
        .ZN(DP_mult_209_n2039) );
  NAND2_X1 DP_mult_209_U1626 ( .A1(DP_mult_209_n1442), .A2(DP_mult_209_n1332), 
        .ZN(DP_mult_209_n2038) );
  XOR2_X1 DP_mult_209_U1625 ( .A(DP_mult_209_n1442), .B(DP_mult_209_n2037), 
        .Z(DP_mult_209_n1065) );
  XOR2_X1 DP_mult_209_U1624 ( .A(DP_mult_209_n1332), .B(DP_mult_209_n1354), 
        .Z(DP_mult_209_n2037) );
  INV_X1 DP_mult_209_U1623 ( .A(DP_mult_209_n2270), .ZN(DP_mult_209_n2266) );
  INV_X1 DP_mult_209_U1622 ( .A(DP_mult_209_n2072), .ZN(DP_mult_209_n2188) );
  INV_X1 DP_mult_209_U1621 ( .A(DP_mult_209_n2282), .ZN(DP_mult_209_n2035) );
  INV_X2 DP_mult_209_U1620 ( .A(DP_mult_209_n2282), .ZN(DP_mult_209_n2036) );
  BUF_X1 DP_mult_209_U1619 ( .A(DP_mult_209_n490), .Z(DP_mult_209_n2108) );
  OAI22_X1 DP_mult_209_U1618 ( .A1(DP_mult_209_n2222), .A2(DP_mult_209_n1733), 
        .B1(DP_mult_209_n1732), .B2(DP_mult_209_n2019), .ZN(DP_mult_209_n2034)
         );
  NAND3_X1 DP_mult_209_U1617 ( .A1(DP_mult_209_n2105), .A2(DP_mult_209_n2106), 
        .A3(DP_mult_209_n2107), .ZN(DP_mult_209_n2032) );
  NAND3_X1 DP_mult_209_U1616 ( .A1(DP_mult_209_n2105), .A2(DP_mult_209_n2106), 
        .A3(DP_mult_209_n2107), .ZN(DP_mult_209_n2033) );
  NAND3_X1 DP_mult_209_U1615 ( .A1(DP_mult_209_n2029), .A2(DP_mult_209_n2030), 
        .A3(DP_mult_209_n2031), .ZN(DP_mult_209_n1074) );
  NAND2_X1 DP_mult_209_U1614 ( .A1(DP_mult_209_n1081), .A2(DP_mult_209_n1083), 
        .ZN(DP_mult_209_n2031) );
  NAND2_X1 DP_mult_209_U1613 ( .A1(DP_mult_209_n1079), .A2(DP_mult_209_n1083), 
        .ZN(DP_mult_209_n2030) );
  NAND2_X1 DP_mult_209_U1612 ( .A1(DP_mult_209_n1079), .A2(DP_mult_209_n1081), 
        .ZN(DP_mult_209_n2029) );
  XOR2_X1 DP_mult_209_U1611 ( .A(DP_mult_209_n1079), .B(DP_mult_209_n2028), 
        .Z(DP_mult_209_n1075) );
  XOR2_X1 DP_mult_209_U1610 ( .A(DP_mult_209_n1081), .B(DP_mult_209_n1083), 
        .Z(DP_mult_209_n2028) );
  OAI22_X1 DP_mult_209_U1609 ( .A1(DP_mult_209_n2220), .A2(DP_mult_209_n1683), 
        .B1(DP_mult_209_n1682), .B2(DP_mult_209_n2246), .ZN(DP_mult_209_n2027)
         );
  INV_X1 DP_mult_209_U1608 ( .A(DP_mult_209_n2183), .ZN(DP_mult_209_n2241) );
  INV_X2 DP_mult_209_U1607 ( .A(DP_mult_209_n2305), .ZN(DP_mult_209_n2303) );
  CLKBUF_X1 DP_mult_209_U1606 ( .A(DP_mult_209_n1027), .Z(DP_mult_209_n2026)
         );
  XOR2_X1 DP_mult_209_U1605 ( .A(DP_mult_209_n1987), .B(DP_pipe03[14]), .Z(
        DP_mult_209_n1666) );
  INV_X1 DP_mult_209_U1604 ( .A(DP_mult_209_n2078), .ZN(DP_mult_209_n2024) );
  INV_X1 DP_mult_209_U1603 ( .A(DP_mult_209_n2078), .ZN(DP_mult_209_n2025) );
  INV_X1 DP_mult_209_U1602 ( .A(DP_mult_209_n1975), .ZN(DP_mult_209_n2023) );
  CLKBUF_X3 DP_mult_209_U1601 ( .A(DP_mult_209_n279), .Z(DP_mult_209_n2022) );
  NOR2_X1 DP_mult_209_U1600 ( .A1(DP_mult_209_n2021), .A2(DP_mult_209_n596), 
        .ZN(DP_mult_209_n594) );
  AND2_X1 DP_mult_209_U1599 ( .A1(DP_mult_209_n595), .A2(DP_mult_209_n609), 
        .ZN(DP_mult_209_n2021) );
  XNOR2_X1 DP_mult_209_U1598 ( .A(DP_coeffs_ff_int[83]), .B(DP_mult_209_n2283), 
        .ZN(DP_mult_209_n1811) );
  INV_X2 DP_mult_209_U1597 ( .A(DP_mult_209_n2188), .ZN(DP_mult_209_n2248) );
  INV_X1 DP_mult_209_U1596 ( .A(DP_mult_209_n2020), .ZN(DP_mult_209_n2018) );
  XOR2_X1 DP_mult_209_U1595 ( .A(DP_coeffs_ff_int[86]), .B(
        DP_coeffs_ff_int[85]), .Z(DP_mult_209_n2183) );
  OR2_X1 DP_mult_209_U1594 ( .A1(DP_mult_209_n788), .A2(DP_mult_209_n775), 
        .ZN(DP_mult_209_n2166) );
  INV_X1 DP_mult_209_U1593 ( .A(DP_mult_209_n2063), .ZN(DP_mult_209_n2017) );
  INV_X1 DP_mult_209_U1592 ( .A(DP_mult_209_n2228), .ZN(DP_mult_209_n2016) );
  INV_X1 DP_mult_209_U1591 ( .A(DP_mult_209_n2086), .ZN(DP_mult_209_n2014) );
  INV_X1 DP_mult_209_U1590 ( .A(DP_mult_209_n2086), .ZN(DP_mult_209_n2015) );
  NOR2_X1 DP_mult_209_U1589 ( .A1(DP_mult_209_n505), .A2(DP_mult_209_n452), 
        .ZN(DP_mult_209_n2013) );
  XNOR2_X1 DP_mult_209_U1588 ( .A(DP_coeffs_ff_int[79]), .B(
        DP_coeffs_ff_int[80]), .ZN(DP_mult_209_n267) );
  INV_X2 DP_mult_209_U1587 ( .A(DP_mult_209_n2259), .ZN(DP_mult_209_n2256) );
  CLKBUF_X1 DP_mult_209_U1586 ( .A(DP_coeffs_ff_int[92]), .Z(DP_mult_209_n2020) );
  INV_X1 DP_mult_209_U1585 ( .A(DP_mult_209_n2239), .ZN(DP_mult_209_n2012) );
  INV_X1 DP_mult_209_U1584 ( .A(DP_mult_209_n2061), .ZN(DP_mult_209_n2011) );
  OR2_X1 DP_mult_209_U1583 ( .A1(DP_mult_209_n558), .A2(DP_mult_209_n563), 
        .ZN(DP_mult_209_n2010) );
  NAND3_X1 DP_mult_209_U1582 ( .A1(DP_mult_209_n2007), .A2(DP_mult_209_n2008), 
        .A3(DP_mult_209_n2009), .ZN(DP_mult_209_n834) );
  NAND2_X1 DP_mult_209_U1581 ( .A1(DP_mult_209_n1210), .A2(DP_mult_209_n1276), 
        .ZN(DP_mult_209_n2009) );
  NAND2_X1 DP_mult_209_U1580 ( .A1(DP_mult_209_n837), .A2(DP_mult_209_n1276), 
        .ZN(DP_mult_209_n2008) );
  NAND2_X1 DP_mult_209_U1579 ( .A1(DP_mult_209_n837), .A2(DP_mult_209_n1210), 
        .ZN(DP_mult_209_n2007) );
  XOR2_X1 DP_mult_209_U1578 ( .A(DP_mult_209_n837), .B(DP_mult_209_n2006), .Z(
        DP_mult_209_n835) );
  XOR2_X1 DP_mult_209_U1577 ( .A(DP_mult_209_n1210), .B(DP_mult_209_n1276), 
        .Z(DP_mult_209_n2006) );
  CLKBUF_X1 DP_mult_209_U1576 ( .A(DP_mult_209_n2166), .Z(DP_mult_209_n2005)
         );
  XOR2_X1 DP_mult_209_U1575 ( .A(DP_mult_209_n2270), .B(DP_pipe03[22]), .Z(
        DP_mult_209_n1683) );
  AND2_X1 DP_mult_209_U1574 ( .A1(DP_mult_209_n525), .A2(DP_mult_209_n511), 
        .ZN(DP_mult_209_n2004) );
  BUF_X2 DP_mult_209_U1573 ( .A(DP_mult_209_n277), .Z(DP_mult_209_n2003) );
  XOR2_X1 DP_mult_209_U1572 ( .A(DP_pipe03[23]), .B(DP_mult_209_n2259), .Z(
        DP_mult_209_n1732) );
  INV_X2 DP_mult_209_U1571 ( .A(DP_mult_209_n2018), .ZN(DP_mult_209_n2258) );
  INV_X1 DP_mult_209_U1570 ( .A(DP_mult_209_n2067), .ZN(DP_mult_209_n2189) );
  AND2_X2 DP_mult_209_U1569 ( .A1(DP_mult_209_n1811), .A2(DP_mult_209_n2236), 
        .ZN(DP_mult_209_n2062) );
  XNOR2_X1 DP_mult_209_U1568 ( .A(DP_mult_209_n1400), .B(DP_mult_209_n1467), 
        .ZN(DP_mult_209_n2002) );
  XNOR2_X1 DP_mult_209_U1567 ( .A(DP_mult_209_n2002), .B(DP_mult_209_n1186), 
        .ZN(DP_mult_209_n1095) );
  XNOR2_X1 DP_mult_209_U1566 ( .A(DP_mult_209_n1947), .B(DP_mult_209_n2278), 
        .ZN(DP_mult_209_n1812) );
  NAND3_X1 DP_mult_209_U1565 ( .A1(DP_mult_209_n1999), .A2(DP_mult_209_n2000), 
        .A3(DP_mult_209_n2001), .ZN(DP_mult_209_n962) );
  NAND2_X1 DP_mult_209_U1564 ( .A1(DP_mult_209_n984), .A2(DP_mult_209_n967), 
        .ZN(DP_mult_209_n2001) );
  NAND2_X1 DP_mult_209_U1563 ( .A1(DP_mult_209_n965), .A2(DP_mult_209_n967), 
        .ZN(DP_mult_209_n2000) );
  NAND2_X1 DP_mult_209_U1562 ( .A1(DP_mult_209_n965), .A2(DP_mult_209_n984), 
        .ZN(DP_mult_209_n1999) );
  XOR2_X1 DP_mult_209_U1561 ( .A(DP_mult_209_n965), .B(DP_mult_209_n1998), .Z(
        DP_mult_209_n963) );
  XOR2_X1 DP_mult_209_U1560 ( .A(DP_mult_209_n984), .B(DP_mult_209_n967), .Z(
        DP_mult_209_n1998) );
  INV_X1 DP_mult_209_U1559 ( .A(DP_pipe03[0]), .ZN(DP_mult_209_n1996) );
  INV_X1 DP_mult_209_U1558 ( .A(DP_pipe03[0]), .ZN(DP_mult_209_n1997) );
  INV_X1 DP_mult_209_U1557 ( .A(DP_mult_209_n2078), .ZN(DP_mult_209_n2216) );
  XOR2_X1 DP_mult_209_U1556 ( .A(DP_coeffs_ff_int[91]), .B(
        DP_coeffs_ff_int[90]), .Z(DP_mult_209_n1815) );
  INV_X2 DP_mult_209_U1555 ( .A(DP_mult_209_n1995), .ZN(DP_mult_209_n2229) );
  XOR2_X1 DP_mult_209_U1554 ( .A(DP_coeffs_ff_int[77]), .B(
        DP_coeffs_ff_int[78]), .Z(DP_mult_209_n1995) );
  BUF_X2 DP_mult_209_U1553 ( .A(DP_mult_209_n251), .Z(DP_mult_209_n2249) );
  CLKBUF_X1 DP_mult_209_U1552 ( .A(DP_mult_209_n2183), .Z(DP_mult_209_n1994)
         );
  INV_X1 DP_mult_209_U1551 ( .A(DP_mult_209_n2187), .ZN(DP_mult_209_n2246) );
  INV_X2 DP_mult_209_U1550 ( .A(DP_mult_209_n2187), .ZN(DP_mult_209_n1993) );
  INV_X2 DP_mult_209_U1549 ( .A(DP_mult_209_n1955), .ZN(DP_mult_209_n2235) );
  INV_X1 DP_mult_209_U1548 ( .A(DP_mult_209_n2061), .ZN(DP_mult_209_n2052) );
  INV_X1 DP_mult_209_U1547 ( .A(DP_mult_209_n2061), .ZN(DP_mult_209_n1991) );
  INV_X1 DP_mult_209_U1546 ( .A(DP_mult_209_n2062), .ZN(DP_mult_209_n1992) );
  AND2_X1 DP_mult_209_U1545 ( .A1(DP_mult_209_n2122), .A2(DP_mult_209_n535), 
        .ZN(DP_mult_209_n1990) );
  XNOR2_X1 DP_mult_209_U1544 ( .A(DP_mult_209_n1950), .B(DP_mult_209_n1990), 
        .ZN(DP_pipe0_coeff_pipe03[3]) );
  AND2_X2 DP_mult_209_U1543 ( .A1(DP_mult_209_n1808), .A2(DP_mult_209_n2063), 
        .ZN(DP_mult_209_n1989) );
  BUF_X1 DP_mult_209_U1542 ( .A(DP_mult_209_n1988), .Z(DP_mult_209_n1987) );
  AND2_X1 DP_mult_209_U1541 ( .A1(DP_mult_209_n675), .A2(DP_mult_209_n1983), 
        .ZN(DP_mult_209_n1986) );
  XNOR2_X1 DP_mult_209_U1540 ( .A(DP_mult_209_n560), .B(DP_mult_209_n1986), 
        .ZN(DP_pipe0_coeff_pipe03[0]) );
  AND2_X1 DP_mult_209_U1539 ( .A1(DP_mult_209_n673), .A2(DP_mult_209_n543), 
        .ZN(DP_mult_209_n1985) );
  XNOR2_X1 DP_mult_209_U1538 ( .A(DP_mult_209_n544), .B(DP_mult_209_n1985), 
        .ZN(DP_pipe0_coeff_pipe03[2]) );
  INV_X1 DP_mult_209_U1537 ( .A(DP_mult_209_n553), .ZN(DP_mult_209_n1984) );
  CLKBUF_X1 DP_mult_209_U1536 ( .A(DP_mult_209_n559), .Z(DP_mult_209_n1983) );
  OR2_X1 DP_mult_209_U1535 ( .A1(DP_mult_209_n1151), .A2(DP_mult_209_n1158), 
        .ZN(DP_mult_209_n1982) );
  AND2_X1 DP_mult_209_U1534 ( .A1(DP_mult_209_n1021), .A2(DP_mult_209_n1038), 
        .ZN(DP_mult_209_n1981) );
  AND2_X1 DP_mult_209_U1533 ( .A1(DP_mult_209_n1111), .A2(DP_mult_209_n1122), 
        .ZN(DP_mult_209_n1980) );
  AND2_X1 DP_mult_209_U1532 ( .A1(DP_mult_209_n1133), .A2(DP_mult_209_n1142), 
        .ZN(DP_mult_209_n1979) );
  AND2_X1 DP_mult_209_U1531 ( .A1(DP_mult_209_n1055), .A2(DP_mult_209_n1070), 
        .ZN(DP_mult_209_n1978) );
  AND2_X1 DP_mult_209_U1530 ( .A1(DP_mult_209_n1179), .A2(DP_mult_209_n1433), 
        .ZN(DP_mult_209_n1977) );
  AND2_X1 DP_mult_209_U1529 ( .A1(DP_mult_209_n1457), .A2(DP_mult_209_n1480), 
        .ZN(DP_mult_209_n1976) );
  AND2_X1 DP_mult_209_U1528 ( .A1(DP_mult_209_n1814), .A2(DP_mult_209_n2117), 
        .ZN(DP_mult_209_n1975) );
  AND2_X1 DP_mult_209_U1527 ( .A1(DP_mult_209_n1151), .A2(DP_mult_209_n1158), 
        .ZN(DP_mult_209_n1974) );
  AND2_X1 DP_mult_209_U1526 ( .A1(DP_mult_209_n1123), .A2(DP_mult_209_n1132), 
        .ZN(DP_mult_209_n1973) );
  AND2_X1 DP_mult_209_U1525 ( .A1(DP_mult_209_n1143), .A2(DP_mult_209_n1150), 
        .ZN(DP_mult_209_n1972) );
  OR2_X1 DP_mult_209_U1524 ( .A1(DP_mult_209_n1179), .A2(DP_mult_209_n1433), 
        .ZN(DP_mult_209_n1971) );
  OR2_X1 DP_mult_209_U1523 ( .A1(DP_mult_209_n1457), .A2(DP_mult_209_n1480), 
        .ZN(DP_mult_209_n1970) );
  AND2_X1 DP_mult_209_U1522 ( .A1(DP_mult_209_n1193), .A2(DP_mult_209_n1481), 
        .ZN(DP_mult_209_n1969) );
  OR2_X1 DP_mult_209_U1521 ( .A1(DP_mult_209_n1055), .A2(DP_mult_209_n1070), 
        .ZN(DP_mult_209_n2168) );
  AND2_X1 DP_mult_209_U1520 ( .A1(DP_mult_209_n1810), .A2(DP_mult_209_n2233), 
        .ZN(DP_mult_209_n2153) );
  INV_X1 DP_mult_209_U1519 ( .A(DP_mult_209_n2153), .ZN(DP_mult_209_n2155) );
  INV_X1 DP_mult_209_U1518 ( .A(DP_mult_209_n1975), .ZN(DP_mult_209_n2158) );
  BUF_X2 DP_mult_209_U1517 ( .A(DP_mult_209_n2203), .Z(DP_mult_209_n2192) );
  BUF_X1 DP_mult_209_U1516 ( .A(DP_mult_209_n279), .Z(DP_mult_209_n2089) );
  INV_X1 DP_mult_209_U1515 ( .A(DP_mult_209_n2205), .ZN(DP_mult_209_n2204) );
  INV_X1 DP_mult_209_U1514 ( .A(DP_mult_209_n2205), .ZN(DP_mult_209_n1968) );
  NAND3_X1 DP_mult_209_U1513 ( .A1(DP_mult_209_n1965), .A2(DP_mult_209_n1966), 
        .A3(DP_mult_209_n1967), .ZN(DP_mult_209_n858) );
  NAND2_X1 DP_mult_209_U1512 ( .A1(DP_mult_209_n882), .A2(DP_mult_209_n863), 
        .ZN(DP_mult_209_n1967) );
  NAND2_X1 DP_mult_209_U1511 ( .A1(DP_mult_209_n880), .A2(DP_mult_209_n863), 
        .ZN(DP_mult_209_n1966) );
  NAND2_X1 DP_mult_209_U1510 ( .A1(DP_mult_209_n880), .A2(DP_mult_209_n882), 
        .ZN(DP_mult_209_n1965) );
  XOR2_X1 DP_mult_209_U1509 ( .A(DP_mult_209_n880), .B(DP_mult_209_n1964), .Z(
        DP_mult_209_n859) );
  XOR2_X1 DP_mult_209_U1508 ( .A(DP_mult_209_n882), .B(DP_mult_209_n863), .Z(
        DP_mult_209_n1964) );
  AND2_X2 DP_mult_209_U1507 ( .A1(DP_mult_209_n1809), .A2(DP_mult_209_n267), 
        .ZN(DP_mult_209_n2066) );
  INV_X1 DP_mult_209_U1506 ( .A(DP_mult_209_n2066), .ZN(DP_mult_209_n2210) );
  INV_X2 DP_mult_209_U1505 ( .A(DP_mult_209_n2066), .ZN(DP_mult_209_n1962) );
  INV_X1 DP_mult_209_U1504 ( .A(DP_mult_209_n2066), .ZN(DP_mult_209_n1963) );
  XOR2_X1 DP_mult_209_U1503 ( .A(DP_coeffs_ff_int[83]), .B(
        DP_coeffs_ff_int[84]), .Z(DP_mult_209_n1961) );
  XOR2_X1 DP_mult_209_U1502 ( .A(DP_coeffs_ff_int[83]), .B(
        DP_coeffs_ff_int[84]), .Z(DP_mult_209_n1960) );
  XOR2_X1 DP_mult_209_U1501 ( .A(DP_pipe03[5]), .B(DP_mult_209_n2278), .Z(
        DP_mult_209_n1650) );
  CLKBUF_X3 DP_mult_209_U1500 ( .A(DP_mult_209_n297), .Z(DP_mult_209_n2044) );
  INV_X1 DP_mult_209_U1499 ( .A(DP_mult_209_n2189), .ZN(DP_mult_209_n2247) );
  INV_X2 DP_mult_209_U1498 ( .A(DP_mult_209_n2189), .ZN(DP_mult_209_n1958) );
  INV_X1 DP_mult_209_U1497 ( .A(DP_mult_209_n2189), .ZN(DP_mult_209_n1959) );
  XOR2_X1 DP_mult_209_U1496 ( .A(DP_coeffs_ff_int[81]), .B(
        DP_coeffs_ff_int[82]), .Z(DP_mult_209_n1955) );
  INV_X1 DP_mult_209_U1495 ( .A(DP_mult_209_n2086), .ZN(DP_mult_209_n1954) );
  INV_X2 DP_mult_209_U1494 ( .A(DP_mult_209_n2283), .ZN(DP_mult_209_n2280) );
  INV_X2 DP_mult_209_U1493 ( .A(DP_mult_209_n2269), .ZN(DP_mult_209_n2268) );
  AND2_X2 DP_mult_209_U1492 ( .A1(DP_mult_209_n1811), .A2(DP_mult_209_n2236), 
        .ZN(DP_mult_209_n2061) );
  INV_X1 DP_mult_209_U1491 ( .A(DP_mult_209_n1988), .ZN(DP_mult_209_n2272) );
  INV_X1 DP_mult_209_U1490 ( .A(DP_mult_209_n1988), .ZN(DP_mult_209_n1952) );
  INV_X1 DP_mult_209_U1489 ( .A(DP_mult_209_n1988), .ZN(DP_mult_209_n1953) );
  INV_X2 DP_mult_209_U1488 ( .A(DP_mult_209_n2087), .ZN(DP_mult_209_n2101) );
  BUF_X1 DP_mult_209_U1487 ( .A(DP_mult_209_n536), .Z(DP_mult_209_n1950) );
  BUF_X1 DP_mult_209_U1486 ( .A(DP_mult_209_n536), .Z(DP_mult_209_n1951) );
  BUF_X1 DP_mult_209_U1485 ( .A(DP_mult_209_n536), .Z(DP_mult_209_n1949) );
  CLKBUF_X1 DP_mult_209_U1484 ( .A(DP_mult_209_n568), .Z(DP_mult_209_n1948) );
  INV_X2 DP_mult_209_U1483 ( .A(DP_mult_209_n2279), .ZN(DP_mult_209_n2276) );
  BUF_X2 DP_mult_209_U1482 ( .A(DP_mult_209_n251), .Z(DP_mult_209_n2250) );
  CLKBUF_X1 DP_mult_209_U1481 ( .A(DP_coeffs_ff_int[85]), .Z(DP_mult_209_n1947) );
  BUF_X1 DP_mult_209_U1480 ( .A(DP_mult_209_n581), .Z(DP_mult_209_n1957) );
  AND2_X1 DP_mult_209_U1479 ( .A1(DP_mult_209_n550), .A2(DP_mult_209_n2100), 
        .ZN(DP_mult_209_n1946) );
  XNOR2_X1 DP_mult_209_U1478 ( .A(DP_mult_209_n551), .B(DP_mult_209_n1946), 
        .ZN(DP_pipe0_coeff_pipe03[1]) );
  BUF_X1 DP_mult_209_U1477 ( .A(DP_mult_209_n1238), .Z(DP_mult_209_n1944) );
  NAND2_X1 DP_mult_209_U1476 ( .A1(DP_mult_209_n1216), .A2(DP_mult_209_n1944), 
        .ZN(DP_mult_209_n1943) );
  INV_X1 DP_mult_209_U1475 ( .A(DP_mult_209_n1943), .ZN(DP_mult_209_n960) );
  XOR2_X1 DP_mult_209_U1474 ( .A(DP_mult_209_n1216), .B(DP_mult_209_n1238), 
        .Z(DP_mult_209_n961) );
  AND2_X2 DP_mult_209_U1473 ( .A1(DP_mult_209_n1807), .A2(DP_mult_209_n2226), 
        .ZN(DP_mult_209_n2086) );
  INV_X1 DP_mult_209_U1472 ( .A(DP_mult_209_n1939), .ZN(DP_mult_209_n1941) );
  INV_X2 DP_mult_209_U1471 ( .A(DP_mult_209_n1939), .ZN(DP_mult_209_n1942) );
  INV_X1 DP_mult_209_U1470 ( .A(DP_mult_209_n1939), .ZN(DP_mult_209_n1940) );
  INV_X1 DP_mult_209_U1469 ( .A(DP_mult_209_n2257), .ZN(DP_mult_209_n1939) );
  AND2_X1 DP_mult_209_U1468 ( .A1(DP_mult_209_n775), .A2(DP_mult_209_n788), 
        .ZN(DP_mult_209_n1956) );
  INV_X1 DP_mult_209_U1467 ( .A(DP_mult_209_n1956), .ZN(DP_mult_209_n474) );
  INV_X2 DP_mult_209_U1466 ( .A(DP_mult_209_n1989), .ZN(DP_mult_209_n2208) );
  INV_X1 DP_mult_209_U1465 ( .A(DP_mult_209_n2205), .ZN(DP_mult_209_n1938) );
  INV_X1 DP_mult_209_U1464 ( .A(DP_coeffs_ff_int[72]), .ZN(DP_mult_209_n1937)
         );
  INV_X1 DP_mult_209_U1463 ( .A(DP_mult_209_n1989), .ZN(DP_mult_209_n2097) );
  BUF_X2 DP_mult_209_U1462 ( .A(DP_mult_209_n2274), .Z(DP_mult_209_n1988) );
  NAND3_X1 DP_mult_209_U1461 ( .A1(DP_mult_209_n1934), .A2(DP_mult_209_n1935), 
        .A3(DP_mult_209_n1936), .ZN(DP_mult_209_n880) );
  NAND2_X1 DP_mult_209_U1460 ( .A1(DP_mult_209_n904), .A2(DP_mult_209_n887), 
        .ZN(DP_mult_209_n1936) );
  NAND2_X1 DP_mult_209_U1459 ( .A1(DP_mult_209_n902), .A2(DP_mult_209_n887), 
        .ZN(DP_mult_209_n1935) );
  NAND2_X1 DP_mult_209_U1458 ( .A1(DP_mult_209_n902), .A2(DP_mult_209_n904), 
        .ZN(DP_mult_209_n1934) );
  XOR2_X1 DP_mult_209_U1457 ( .A(DP_mult_209_n902), .B(DP_mult_209_n1933), .Z(
        DP_mult_209_n881) );
  XOR2_X1 DP_mult_209_U1456 ( .A(DP_mult_209_n904), .B(DP_mult_209_n887), .Z(
        DP_mult_209_n1933) );
  CLKBUF_X1 DP_mult_209_U1455 ( .A(DP_mult_209_n1237), .Z(DP_mult_209_n1945)
         );
  NAND3_X1 DP_mult_209_U1454 ( .A1(DP_mult_209_n1930), .A2(DP_mult_209_n1931), 
        .A3(DP_mult_209_n1932), .ZN(DP_mult_209_n884) );
  NAND2_X1 DP_mult_209_U1453 ( .A1(DP_mult_209_n891), .A2(DP_mult_209_n895), 
        .ZN(DP_mult_209_n1932) );
  NAND2_X1 DP_mult_209_U1452 ( .A1(DP_mult_209_n908), .A2(DP_mult_209_n895), 
        .ZN(DP_mult_209_n1931) );
  NAND2_X1 DP_mult_209_U1451 ( .A1(DP_mult_209_n908), .A2(DP_mult_209_n891), 
        .ZN(DP_mult_209_n1930) );
  XOR2_X1 DP_mult_209_U1450 ( .A(DP_mult_209_n908), .B(DP_mult_209_n1929), .Z(
        DP_mult_209_n885) );
  XOR2_X1 DP_mult_209_U1449 ( .A(DP_mult_209_n891), .B(DP_mult_209_n895), .Z(
        DP_mult_209_n1929) );
  INV_X2 DP_mult_209_U1448 ( .A(DP_mult_209_n2188), .ZN(DP_mult_209_n2019) );
  HA_X1 DP_mult_209_U798 ( .A(DP_mult_209_n1456), .B(DP_mult_209_n1479), .CO(
        DP_mult_209_n1180), .S(DP_mult_209_n1181) );
  FA_X1 DP_mult_209_U797 ( .A(DP_mult_209_n1455), .B(DP_mult_209_n1478), .CI(
        DP_mult_209_n1180), .CO(DP_mult_209_n1178), .S(DP_mult_209_n1179) );
  HA_X1 DP_mult_209_U796 ( .A(DP_mult_209_n1432), .B(DP_mult_209_n1477), .CO(
        DP_mult_209_n1176), .S(DP_mult_209_n1177) );
  FA_X1 DP_mult_209_U795 ( .A(DP_mult_209_n1191), .B(DP_mult_209_n1454), .CI(
        DP_mult_209_n1177), .CO(DP_mult_209_n1174), .S(DP_mult_209_n1175) );
  FA_X1 DP_mult_209_U794 ( .A(DP_mult_209_n1476), .B(DP_mult_209_n1453), .CI(
        DP_mult_209_n1431), .CO(DP_mult_209_n1172), .S(DP_mult_209_n1173) );
  FA_X1 DP_mult_209_U793 ( .A(DP_mult_209_n1409), .B(DP_mult_209_n1176), .CI(
        DP_mult_209_n1173), .CO(DP_mult_209_n1170), .S(DP_mult_209_n1171) );
  HA_X1 DP_mult_209_U792 ( .A(DP_mult_209_n1408), .B(DP_mult_209_n1430), .CO(
        DP_mult_209_n1168), .S(DP_mult_209_n1169) );
  FA_X1 DP_mult_209_U791 ( .A(DP_mult_209_n1452), .B(DP_mult_209_n1475), .CI(
        DP_mult_209_n1190), .CO(DP_mult_209_n1166), .S(DP_mult_209_n1167) );
  FA_X1 DP_mult_209_U790 ( .A(DP_mult_209_n1172), .B(DP_mult_209_n1169), .CI(
        DP_mult_209_n1167), .CO(DP_mult_209_n1164), .S(DP_mult_209_n1165) );
  FA_X1 DP_mult_209_U789 ( .A(DP_mult_209_n1451), .B(DP_mult_209_n1474), .CI(
        DP_mult_209_n1407), .CO(DP_mult_209_n1162), .S(DP_mult_209_n1163) );
  FA_X1 DP_mult_209_U788 ( .A(DP_mult_209_n1168), .B(DP_mult_209_n1429), .CI(
        DP_mult_209_n1166), .CO(DP_mult_209_n1160), .S(DP_mult_209_n1161) );
  FA_X1 DP_mult_209_U787 ( .A(DP_mult_209_n1163), .B(DP_mult_209_n1385), .CI(
        DP_mult_209_n1164), .CO(DP_mult_209_n1158), .S(DP_mult_209_n1159) );
  HA_X1 DP_mult_209_U786 ( .A(DP_mult_209_n1384), .B(DP_mult_209_n1406), .CO(
        DP_mult_209_n1156), .S(DP_mult_209_n1157) );
  FA_X1 DP_mult_209_U785 ( .A(DP_mult_209_n1450), .B(DP_mult_209_n1428), .CI(
        DP_mult_209_n1189), .CO(DP_mult_209_n1154), .S(DP_mult_209_n1155) );
  FA_X1 DP_mult_209_U784 ( .A(DP_mult_209_n1157), .B(DP_mult_209_n1473), .CI(
        DP_mult_209_n1162), .CO(DP_mult_209_n1152), .S(DP_mult_209_n1153) );
  FA_X1 DP_mult_209_U783 ( .A(DP_mult_209_n1160), .B(DP_mult_209_n1155), .CI(
        DP_mult_209_n1153), .CO(DP_mult_209_n1150), .S(DP_mult_209_n1151) );
  FA_X1 DP_mult_209_U782 ( .A(DP_mult_209_n1383), .B(DP_mult_209_n1472), .CI(
        DP_mult_209_n1405), .CO(DP_mult_209_n1148), .S(DP_mult_209_n1149) );
  FA_X1 DP_mult_209_U781 ( .A(DP_mult_209_n1427), .B(DP_mult_209_n1449), .CI(
        DP_mult_209_n1156), .CO(DP_mult_209_n1146), .S(DP_mult_209_n1147) );
  FA_X1 DP_mult_209_U780 ( .A(DP_mult_209_n1361), .B(DP_mult_209_n1154), .CI(
        DP_mult_209_n1149), .CO(DP_mult_209_n1144), .S(DP_mult_209_n1145) );
  FA_X1 DP_mult_209_U779 ( .A(DP_mult_209_n1152), .B(DP_mult_209_n1147), .CI(
        DP_mult_209_n1145), .CO(DP_mult_209_n1142), .S(DP_mult_209_n1143) );
  HA_X1 DP_mult_209_U778 ( .A(DP_mult_209_n1360), .B(DP_mult_209_n1382), .CO(
        DP_mult_209_n1140), .S(DP_mult_209_n1141) );
  FA_X1 DP_mult_209_U777 ( .A(DP_mult_209_n1471), .B(DP_mult_209_n1426), .CI(
        DP_mult_209_n1188), .CO(DP_mult_209_n1138), .S(DP_mult_209_n1139) );
  FA_X1 DP_mult_209_U776 ( .A(DP_mult_209_n1404), .B(DP_mult_209_n1448), .CI(
        DP_mult_209_n1141), .CO(DP_mult_209_n1136), .S(DP_mult_209_n1137) );
  FA_X1 DP_mult_209_U775 ( .A(DP_mult_209_n1146), .B(DP_mult_209_n1148), .CI(
        DP_mult_209_n1139), .CO(DP_mult_209_n1134), .S(DP_mult_209_n1135) );
  FA_X1 DP_mult_209_U774 ( .A(DP_mult_209_n1144), .B(DP_mult_209_n1137), .CI(
        DP_mult_209_n1135), .CO(DP_mult_209_n1132), .S(DP_mult_209_n1133) );
  FA_X1 DP_mult_209_U773 ( .A(DP_mult_209_n1381), .B(DP_mult_209_n1470), .CI(
        DP_mult_209_n1359), .CO(DP_mult_209_n1130), .S(DP_mult_209_n1131) );
  FA_X1 DP_mult_209_U772 ( .A(DP_mult_209_n1403), .B(DP_mult_209_n1447), .CI(
        DP_mult_209_n1425), .CO(DP_mult_209_n1128), .S(DP_mult_209_n1129) );
  FA_X1 DP_mult_209_U771 ( .A(DP_mult_209_n1138), .B(DP_mult_209_n1140), .CI(
        DP_mult_209_n1337), .CO(DP_mult_209_n1126), .S(DP_mult_209_n1127) );
  FA_X1 DP_mult_209_U770 ( .A(DP_mult_209_n1131), .B(DP_mult_209_n1129), .CI(
        DP_mult_209_n1136), .CO(DP_mult_209_n1124), .S(DP_mult_209_n1125) );
  FA_X1 DP_mult_209_U769 ( .A(DP_mult_209_n1127), .B(DP_mult_209_n1134), .CI(
        DP_mult_209_n1125), .CO(DP_mult_209_n1122), .S(DP_mult_209_n1123) );
  HA_X1 DP_mult_209_U768 ( .A(DP_mult_209_n1336), .B(DP_mult_209_n1358), .CO(
        DP_mult_209_n1120), .S(DP_mult_209_n1121) );
  FA_X1 DP_mult_209_U767 ( .A(DP_mult_209_n1380), .B(DP_mult_209_n1402), .CI(
        DP_mult_209_n1187), .CO(DP_mult_209_n1118), .S(DP_mult_209_n1119) );
  FA_X1 DP_mult_209_U766 ( .A(DP_mult_209_n1424), .B(DP_mult_209_n1469), .CI(
        DP_mult_209_n1446), .CO(DP_mult_209_n1116), .S(DP_mult_209_n1117) );
  FA_X1 DP_mult_209_U765 ( .A(DP_mult_209_n1130), .B(DP_mult_209_n1121), .CI(
        DP_mult_209_n1128), .CO(DP_mult_209_n1114), .S(DP_mult_209_n1115) );
  FA_X1 DP_mult_209_U764 ( .A(DP_mult_209_n1119), .B(DP_mult_209_n1117), .CI(
        DP_mult_209_n1126), .CO(DP_mult_209_n1112), .S(DP_mult_209_n1113) );
  FA_X1 DP_mult_209_U763 ( .A(DP_mult_209_n1124), .B(DP_mult_209_n1115), .CI(
        DP_mult_209_n1113), .CO(DP_mult_209_n1110), .S(DP_mult_209_n1111) );
  FA_X1 DP_mult_209_U762 ( .A(DP_mult_209_n1335), .B(DP_mult_209_n1468), .CI(
        DP_mult_209_n1357), .CO(DP_mult_209_n1108), .S(DP_mult_209_n1109) );
  FA_X1 DP_mult_209_U761 ( .A(DP_mult_209_n1379), .B(DP_mult_209_n1445), .CI(
        DP_mult_209_n1401), .CO(DP_mult_209_n1106), .S(DP_mult_209_n1107) );
  FA_X1 DP_mult_209_U760 ( .A(DP_mult_209_n1120), .B(DP_mult_209_n1423), .CI(
        DP_mult_209_n1118), .CO(DP_mult_209_n1104), .S(DP_mult_209_n1105) );
  FA_X1 DP_mult_209_U759 ( .A(DP_mult_209_n1313), .B(DP_mult_209_n1116), .CI(
        DP_mult_209_n1107), .CO(DP_mult_209_n1102), .S(DP_mult_209_n1103) );
  FA_X1 DP_mult_209_U758 ( .A(DP_mult_209_n1114), .B(DP_mult_209_n1109), .CI(
        DP_mult_209_n1105), .CO(DP_mult_209_n1100), .S(DP_mult_209_n1101) );
  FA_X1 DP_mult_209_U757 ( .A(DP_mult_209_n1103), .B(DP_mult_209_n1112), .CI(
        DP_mult_209_n1101), .CO(DP_mult_209_n1098), .S(DP_mult_209_n1099) );
  HA_X1 DP_mult_209_U756 ( .A(DP_mult_209_n1312), .B(DP_mult_209_n1334), .CO(
        DP_mult_209_n1096), .S(DP_mult_209_n1097) );
  FA_X1 DP_mult_209_U754 ( .A(DP_mult_209_n1444), .B(DP_mult_209_n1356), .CI(
        DP_mult_209_n1378), .CO(DP_mult_209_n1092), .S(DP_mult_209_n1093) );
  FA_X1 DP_mult_209_U753 ( .A(DP_mult_209_n1097), .B(DP_mult_209_n1422), .CI(
        DP_mult_209_n1108), .CO(DP_mult_209_n1090), .S(DP_mult_209_n1091) );
  FA_X1 DP_mult_209_U752 ( .A(DP_mult_209_n1095), .B(DP_mult_209_n1106), .CI(
        DP_mult_209_n1093), .CO(DP_mult_209_n1088), .S(DP_mult_209_n1089) );
  FA_X1 DP_mult_209_U751 ( .A(DP_mult_209_n1102), .B(DP_mult_209_n1104), .CI(
        DP_mult_209_n1091), .CO(DP_mult_209_n1086), .S(DP_mult_209_n1087) );
  FA_X1 DP_mult_209_U750 ( .A(DP_mult_209_n1100), .B(DP_mult_209_n1089), .CI(
        DP_mult_209_n1087), .CO(DP_mult_209_n1084), .S(DP_mult_209_n1085) );
  FA_X1 DP_mult_209_U749 ( .A(DP_mult_209_n1311), .B(DP_mult_209_n1466), .CI(
        DP_mult_209_n1333), .CO(DP_mult_209_n1082), .S(DP_mult_209_n1083) );
  FA_X1 DP_mult_209_U748 ( .A(DP_mult_209_n1355), .B(DP_mult_209_n1443), .CI(
        DP_mult_209_n1377), .CO(DP_mult_209_n1080), .S(DP_mult_209_n1081) );
  FA_X1 DP_mult_209_U747 ( .A(DP_mult_209_n1399), .B(DP_mult_209_n1421), .CI(
        DP_mult_209_n1096), .CO(DP_mult_209_n1078), .S(DP_mult_209_n1079) );
  FA_X1 DP_mult_209_U746 ( .A(DP_mult_209_n1289), .B(DP_mult_209_n1094), .CI(
        DP_mult_209_n1092), .CO(DP_mult_209_n1076), .S(DP_mult_209_n1077) );
  FA_X1 DP_mult_209_U744 ( .A(DP_mult_209_n1088), .B(DP_mult_209_n1090), .CI(
        DP_mult_209_n1077), .CO(DP_mult_209_n1072), .S(DP_mult_209_n1073) );
  FA_X1 DP_mult_209_U743 ( .A(DP_mult_209_n1086), .B(DP_mult_209_n1075), .CI(
        DP_mult_209_n1073), .CO(DP_mult_209_n1070), .S(DP_mult_209_n1071) );
  HA_X1 DP_mult_209_U742 ( .A(DP_mult_209_n1288), .B(DP_mult_209_n1310), .CO(
        DP_mult_209_n1068), .S(DP_mult_209_n1069) );
  FA_X1 DP_mult_209_U741 ( .A(DP_mult_209_n1465), .B(DP_mult_209_n1376), .CI(
        DP_mult_209_n1185), .CO(DP_mult_209_n1066), .S(DP_mult_209_n1067) );
  FA_X1 DP_mult_209_U739 ( .A(DP_mult_209_n1398), .B(DP_mult_209_n1420), .CI(
        DP_mult_209_n1069), .CO(DP_mult_209_n1062), .S(DP_mult_209_n1063) );
  FA_X1 DP_mult_209_U738 ( .A(DP_mult_209_n1080), .B(DP_mult_209_n1082), .CI(
        DP_mult_209_n1078), .CO(DP_mult_209_n1060), .S(DP_mult_209_n1061) );
  FA_X1 DP_mult_209_U737 ( .A(DP_mult_209_n1067), .B(DP_mult_209_n1065), .CI(
        DP_mult_209_n1076), .CO(DP_mult_209_n1058), .S(DP_mult_209_n1059) );
  FA_X1 DP_mult_209_U736 ( .A(DP_mult_209_n1074), .B(DP_mult_209_n1063), .CI(
        DP_mult_209_n1061), .CO(DP_mult_209_n1056), .S(DP_mult_209_n1057) );
  FA_X1 DP_mult_209_U735 ( .A(DP_mult_209_n1072), .B(DP_mult_209_n1059), .CI(
        DP_mult_209_n1057), .CO(DP_mult_209_n1054), .S(DP_mult_209_n1055) );
  FA_X1 DP_mult_209_U734 ( .A(DP_mult_209_n1287), .B(DP_mult_209_n1464), .CI(
        DP_mult_209_n1309), .CO(DP_mult_209_n1052), .S(DP_mult_209_n1053) );
  FA_X1 DP_mult_209_U733 ( .A(DP_mult_209_n1331), .B(DP_mult_209_n1353), .CI(
        DP_mult_209_n1375), .CO(DP_mult_209_n1050), .S(DP_mult_209_n1051) );
  FA_X1 DP_mult_209_U732 ( .A(DP_mult_209_n1397), .B(DP_mult_209_n1441), .CI(
        DP_mult_209_n1419), .CO(DP_mult_209_n1048), .S(DP_mult_209_n1049) );
  FA_X1 DP_mult_209_U731 ( .A(DP_mult_209_n1064), .B(DP_mult_209_n1068), .CI(
        DP_mult_209_n1066), .CO(DP_mult_209_n1046), .S(DP_mult_209_n1047) );
  FA_X1 DP_mult_209_U730 ( .A(DP_mult_209_n1049), .B(DP_mult_209_n1265), .CI(
        DP_mult_209_n1051), .CO(DP_mult_209_n1044), .S(DP_mult_209_n1045) );
  FA_X1 DP_mult_209_U729 ( .A(DP_mult_209_n1062), .B(DP_mult_209_n1053), .CI(
        DP_mult_209_n1060), .CO(DP_mult_209_n1042), .S(DP_mult_209_n1043) );
  FA_X1 DP_mult_209_U728 ( .A(DP_mult_209_n1045), .B(DP_mult_209_n1047), .CI(
        DP_mult_209_n1058), .CO(DP_mult_209_n1040), .S(DP_mult_209_n1041) );
  FA_X1 DP_mult_209_U727 ( .A(DP_mult_209_n1056), .B(DP_mult_209_n1043), .CI(
        DP_mult_209_n1041), .CO(DP_mult_209_n1038), .S(DP_mult_209_n1039) );
  HA_X1 DP_mult_209_U726 ( .A(DP_mult_209_n1264), .B(DP_mult_209_n1286), .CO(
        DP_mult_209_n1036), .S(DP_mult_209_n1037) );
  FA_X1 DP_mult_209_U725 ( .A(DP_mult_209_n1308), .B(DP_mult_209_n1374), .CI(
        DP_mult_209_n1184), .CO(DP_mult_209_n1034), .S(DP_mult_209_n1035) );
  FA_X1 DP_mult_209_U724 ( .A(DP_mult_209_n1463), .B(DP_mult_209_n1396), .CI(
        DP_mult_209_n1330), .CO(DP_mult_209_n1032), .S(DP_mult_209_n1033) );
  FA_X1 DP_mult_209_U723 ( .A(DP_mult_209_n1352), .B(DP_mult_209_n1418), .CI(
        DP_mult_209_n1440), .CO(DP_mult_209_n1030), .S(DP_mult_209_n1031) );
  FA_X1 DP_mult_209_U722 ( .A(DP_mult_209_n1052), .B(DP_mult_209_n1037), .CI(
        DP_mult_209_n1050), .CO(DP_mult_209_n1028), .S(DP_mult_209_n1029) );
  FA_X1 DP_mult_209_U720 ( .A(DP_mult_209_n1046), .B(DP_mult_209_n1035), .CI(
        DP_mult_209_n1029), .CO(DP_mult_209_n1024), .S(DP_mult_209_n1025) );
  FA_X1 DP_mult_209_U718 ( .A(DP_mult_209_n1040), .B(DP_mult_209_n1025), .CI(
        DP_mult_209_n1023), .CO(DP_mult_209_n1020), .S(DP_mult_209_n1021) );
  FA_X1 DP_mult_209_U716 ( .A(DP_mult_209_n1307), .B(DP_mult_209_n1329), .CI(
        DP_mult_209_n1373), .CO(DP_mult_209_n1016), .S(DP_mult_209_n1017) );
  FA_X1 DP_mult_209_U714 ( .A(DP_mult_209_n1036), .B(DP_mult_209_n1439), .CI(
        DP_mult_209_n1032), .CO(DP_mult_209_n1012), .S(DP_mult_209_n1013) );
  FA_X1 DP_mult_209_U713 ( .A(DP_mult_209_n1030), .B(DP_mult_209_n1034), .CI(
        DP_mult_209_n1241), .CO(DP_mult_209_n1010), .S(DP_mult_209_n1011) );
  FA_X1 DP_mult_209_U712 ( .A(DP_mult_209_n1019), .B(DP_mult_209_n1015), .CI(
        DP_mult_209_n1017), .CO(DP_mult_209_n1008), .S(DP_mult_209_n1009) );
  FA_X1 DP_mult_209_U711 ( .A(DP_mult_209_n1013), .B(DP_mult_209_n1028), .CI(
        DP_mult_209_n1026), .CO(DP_mult_209_n1006), .S(DP_mult_209_n1007) );
  FA_X1 DP_mult_209_U710 ( .A(DP_mult_209_n1009), .B(DP_mult_209_n1011), .CI(
        DP_mult_209_n1024), .CO(DP_mult_209_n1004), .S(DP_mult_209_n1005) );
  FA_X1 DP_mult_209_U709 ( .A(DP_mult_209_n1022), .B(DP_mult_209_n1007), .CI(
        DP_mult_209_n1005), .CO(DP_mult_209_n1002), .S(DP_mult_209_n1003) );
  HA_X1 DP_mult_209_U708 ( .A(DP_mult_209_n1240), .B(DP_mult_209_n1262), .CO(
        DP_mult_209_n1000), .S(DP_mult_209_n1001) );
  FA_X1 DP_mult_209_U707 ( .A(DP_mult_209_n1461), .B(DP_mult_209_n1350), .CI(
        DP_mult_209_n1183), .CO(DP_mult_209_n998), .S(DP_mult_209_n999) );
  FA_X1 DP_mult_209_U706 ( .A(DP_mult_209_n1438), .B(DP_mult_209_n1284), .CI(
        DP_mult_209_n1372), .CO(DP_mult_209_n996), .S(DP_mult_209_n997) );
  FA_X1 DP_mult_209_U705 ( .A(DP_mult_209_n1328), .B(DP_mult_209_n1416), .CI(
        DP_mult_209_n1306), .CO(DP_mult_209_n994), .S(DP_mult_209_n995) );
  FA_X1 DP_mult_209_U703 ( .A(DP_mult_209_n1014), .B(DP_mult_209_n1016), .CI(
        DP_mult_209_n995), .CO(DP_mult_209_n990), .S(DP_mult_209_n991) );
  FA_X1 DP_mult_209_U702 ( .A(DP_mult_209_n999), .B(DP_mult_209_n997), .CI(
        DP_mult_209_n1012), .CO(DP_mult_209_n988), .S(DP_mult_209_n989) );
  FA_X1 DP_mult_209_U701 ( .A(DP_mult_209_n993), .B(DP_mult_209_n1010), .CI(
        DP_mult_209_n1008), .CO(DP_mult_209_n986), .S(DP_mult_209_n987) );
  FA_X1 DP_mult_209_U700 ( .A(DP_mult_209_n989), .B(DP_mult_209_n991), .CI(
        DP_mult_209_n1006), .CO(DP_mult_209_n984), .S(DP_mult_209_n985) );
  FA_X1 DP_mult_209_U699 ( .A(DP_mult_209_n1004), .B(DP_mult_209_n987), .CI(
        DP_mult_209_n985), .CO(DP_mult_209_n982), .S(DP_mult_209_n983) );
  FA_X1 DP_mult_209_U698 ( .A(DP_mult_209_n1239), .B(DP_mult_209_n1349), .CI(
        DP_mult_209_n1261), .CO(DP_mult_209_n980), .S(DP_mult_209_n981) );
  FA_X1 DP_mult_209_U697 ( .A(DP_mult_209_n1460), .B(DP_mult_209_n1371), .CI(
        DP_mult_209_n1283), .CO(DP_mult_209_n978), .S(DP_mult_209_n979) );
  FA_X1 DP_mult_209_U696 ( .A(DP_mult_209_n1305), .B(DP_mult_209_n1437), .CI(
        DP_mult_209_n1327), .CO(DP_mult_209_n976), .S(DP_mult_209_n977) );
  FA_X1 DP_mult_209_U695 ( .A(DP_mult_209_n1393), .B(DP_mult_209_n1415), .CI(
        DP_mult_209_n1000), .CO(DP_mult_209_n974), .S(DP_mult_209_n975) );
  FA_X1 DP_mult_209_U694 ( .A(DP_mult_209_n994), .B(DP_mult_209_n996), .CI(
        DP_mult_209_n1217), .CO(DP_mult_209_n972), .S(DP_mult_209_n973) );
  FA_X1 DP_mult_209_U693 ( .A(DP_mult_209_n977), .B(DP_mult_209_n998), .CI(
        DP_mult_209_n979), .CO(DP_mult_209_n970), .S(DP_mult_209_n971) );
  FA_X1 DP_mult_209_U692 ( .A(DP_mult_209_n992), .B(DP_mult_209_n981), .CI(
        DP_mult_209_n975), .CO(DP_mult_209_n968), .S(DP_mult_209_n969) );
  FA_X1 DP_mult_209_U691 ( .A(DP_mult_209_n973), .B(DP_mult_209_n990), .CI(
        DP_mult_209_n988), .CO(DP_mult_209_n966), .S(DP_mult_209_n967) );
  FA_X1 DP_mult_209_U690 ( .A(DP_mult_209_n969), .B(DP_mult_209_n971), .CI(
        DP_mult_209_n986), .CO(DP_mult_209_n964), .S(DP_mult_209_n965) );
  FA_X1 DP_mult_209_U687 ( .A(DP_mult_209_n1182), .B(DP_mult_209_n1260), .CI(
        DP_mult_209_n1348), .CO(DP_mult_209_n958), .S(DP_mult_209_n959) );
  FA_X1 DP_mult_209_U686 ( .A(DP_mult_209_n1459), .B(DP_mult_209_n1370), .CI(
        DP_mult_209_n1436), .CO(DP_mult_209_n956), .S(DP_mult_209_n957) );
  FA_X1 DP_mult_209_U684 ( .A(DP_mult_209_n1326), .B(DP_mult_209_n1392), .CI(
        DP_mult_209_n961), .CO(DP_mult_209_n952), .S(DP_mult_209_n953) );
  FA_X1 DP_mult_209_U683 ( .A(DP_mult_209_n976), .B(DP_mult_209_n980), .CI(
        DP_mult_209_n978), .CO(DP_mult_209_n950), .S(DP_mult_209_n951) );
  FA_X1 DP_mult_209_U682 ( .A(DP_mult_209_n955), .B(DP_mult_209_n974), .CI(
        DP_mult_209_n957), .CO(DP_mult_209_n948), .S(DP_mult_209_n949) );
  FA_X1 DP_mult_209_U680 ( .A(DP_mult_209_n951), .B(DP_mult_209_n970), .CI(
        DP_mult_209_n968), .CO(DP_mult_209_n944), .S(DP_mult_209_n945) );
  FA_X1 DP_mult_209_U679 ( .A(DP_mult_209_n947), .B(DP_mult_209_n949), .CI(
        DP_mult_209_n966), .CO(DP_mult_209_n942), .S(DP_mult_209_n943) );
  FA_X1 DP_mult_209_U675 ( .A(DP_mult_209_n1259), .B(DP_mult_209_n1347), .CI(
        DP_mult_209_n1303), .CO(DP_mult_209_n936), .S(DP_mult_209_n937) );
  FA_X1 DP_mult_209_U674 ( .A(DP_mult_209_n1391), .B(DP_mult_209_n1369), .CI(
        DP_mult_209_n1281), .CO(DP_mult_209_n934), .S(DP_mult_209_n935) );
  FA_X1 DP_mult_209_U673 ( .A(DP_mult_209_n1325), .B(DP_mult_209_n1435), .CI(
        DP_mult_209_n1413), .CO(DP_mult_209_n932), .S(DP_mult_209_n933) );
  FA_X1 DP_mult_209_U672 ( .A(DP_mult_209_n1458), .B(DP_mult_209_n960), .CI(
        DP_mult_209_n939), .CO(DP_mult_209_n930), .S(DP_mult_209_n931) );
  FA_X1 DP_mult_209_U671 ( .A(DP_mult_209_n954), .B(DP_mult_209_n958), .CI(
        DP_mult_209_n956), .CO(DP_mult_209_n928), .S(DP_mult_209_n929) );
  FA_X1 DP_mult_209_U670 ( .A(DP_mult_209_n937), .B(DP_mult_209_n933), .CI(
        DP_mult_209_n952), .CO(DP_mult_209_n926), .S(DP_mult_209_n927) );
  FA_X1 DP_mult_209_U669 ( .A(DP_mult_209_n950), .B(DP_mult_209_n935), .CI(
        DP_mult_209_n931), .CO(DP_mult_209_n924), .S(DP_mult_209_n925) );
  FA_X1 DP_mult_209_U668 ( .A(DP_mult_209_n929), .B(DP_mult_209_n948), .CI(
        DP_mult_209_n946), .CO(DP_mult_209_n922), .S(DP_mult_209_n923) );
  FA_X1 DP_mult_209_U667 ( .A(DP_mult_209_n925), .B(DP_mult_209_n927), .CI(
        DP_mult_209_n944), .CO(DP_mult_209_n920), .S(DP_mult_209_n921) );
  FA_X1 DP_mult_209_U664 ( .A(DP_mult_209_n1214), .B(DP_mult_209_n917), .CI(
        DP_mult_209_n1302), .CO(DP_mult_209_n914), .S(DP_mult_209_n915) );
  FA_X1 DP_mult_209_U663 ( .A(DP_mult_209_n1236), .B(DP_mult_209_n1412), .CI(
        DP_mult_209_n1258), .CO(DP_mult_209_n912), .S(DP_mult_209_n913) );
  FA_X1 DP_mult_209_U662 ( .A(DP_mult_209_n1324), .B(DP_mult_209_n1280), .CI(
        DP_mult_209_n1346), .CO(DP_mult_209_n910), .S(DP_mult_209_n911) );
  FA_X1 DP_mult_209_U661 ( .A(DP_mult_209_n1368), .B(DP_mult_209_n1390), .CI(
        DP_mult_209_n938), .CO(DP_mult_209_n908), .S(DP_mult_209_n909) );
  FA_X1 DP_mult_209_U660 ( .A(DP_mult_209_n932), .B(DP_mult_209_n936), .CI(
        DP_mult_209_n934), .CO(DP_mult_209_n906), .S(DP_mult_209_n907) );
  FA_X1 DP_mult_209_U659 ( .A(DP_mult_209_n913), .B(DP_mult_209_n911), .CI(
        DP_mult_209_n915), .CO(DP_mult_209_n904), .S(DP_mult_209_n905) );
  FA_X1 DP_mult_209_U658 ( .A(DP_mult_209_n909), .B(DP_mult_209_n930), .CI(
        DP_mult_209_n928), .CO(DP_mult_209_n902), .S(DP_mult_209_n903) );
  FA_X1 DP_mult_209_U657 ( .A(DP_mult_209_n907), .B(DP_mult_209_n926), .CI(
        DP_mult_209_n905), .CO(DP_mult_209_n900), .S(DP_mult_209_n901) );
  FA_X1 DP_mult_209_U656 ( .A(DP_mult_209_n903), .B(DP_mult_209_n924), .CI(
        DP_mult_209_n922), .CO(DP_mult_209_n898), .S(DP_mult_209_n899) );
  FA_X1 DP_mult_209_U654 ( .A(DP_mult_209_n1235), .B(DP_mult_209_n1213), .CI(
        DP_mult_209_n1411), .CO(DP_mult_209_n894), .S(DP_mult_209_n895) );
  FA_X1 DP_mult_209_U653 ( .A(DP_mult_209_n2034), .B(DP_mult_209_n1323), .CI(
        DP_mult_209_n1279), .CO(DP_mult_209_n892), .S(DP_mult_209_n893) );
  FA_X1 DP_mult_209_U652 ( .A(DP_mult_209_n1257), .B(DP_mult_209_n1301), .CI(
        DP_mult_209_n1345), .CO(DP_mult_209_n890), .S(DP_mult_209_n891) );
  FA_X1 DP_mult_209_U651 ( .A(DP_mult_209_n1367), .B(DP_mult_209_n1389), .CI(
        DP_mult_209_n1434), .CO(DP_mult_209_n888), .S(DP_mult_209_n889) );
  FA_X1 DP_mult_209_U650 ( .A(DP_mult_209_n910), .B(DP_mult_209_n912), .CI(
        DP_mult_209_n914), .CO(DP_mult_209_n886), .S(DP_mult_209_n887) );
  FA_X1 DP_mult_209_U648 ( .A(DP_mult_209_n906), .B(DP_mult_209_n893), .CI(
        DP_mult_209_n889), .CO(DP_mult_209_n882), .S(DP_mult_209_n883) );
  FA_X1 DP_mult_209_U646 ( .A(DP_mult_209_n883), .B(DP_mult_209_n885), .CI(
        DP_mult_209_n900), .CO(DP_mult_209_n878), .S(DP_mult_209_n879) );
  FA_X1 DP_mult_209_U645 ( .A(DP_mult_209_n898), .B(DP_mult_209_n881), .CI(
        DP_mult_209_n879), .CO(DP_mult_209_n876), .S(DP_mult_209_n877) );
  FA_X1 DP_mult_209_U643 ( .A(DP_mult_209_n1388), .B(DP_mult_209_n1278), .CI(
        DP_mult_209_n875), .CO(DP_mult_209_n872), .S(DP_mult_209_n873) );
  FA_X1 DP_mult_209_U642 ( .A(DP_mult_209_n1366), .B(DP_mult_209_n1212), .CI(
        DP_mult_209_n1344), .CO(DP_mult_209_n870), .S(DP_mult_209_n871) );
  FA_X1 DP_mult_209_U641 ( .A(DP_mult_209_n1234), .B(DP_mult_209_n1322), .CI(
        DP_mult_209_n1256), .CO(DP_mult_209_n868), .S(DP_mult_209_n869) );
  FA_X1 DP_mult_209_U640 ( .A(DP_mult_209_n894), .B(DP_mult_209_n1300), .CI(
        DP_mult_209_n892), .CO(DP_mult_209_n866), .S(DP_mult_209_n867) );
  FA_X1 DP_mult_209_U639 ( .A(DP_mult_209_n869), .B(DP_mult_209_n890), .CI(
        DP_mult_209_n871), .CO(DP_mult_209_n864), .S(DP_mult_209_n865) );
  FA_X1 DP_mult_209_U637 ( .A(DP_mult_209_n884), .B(DP_mult_209_n867), .CI(
        DP_mult_209_n865), .CO(DP_mult_209_n860), .S(DP_mult_209_n861) );
  FA_X1 DP_mult_209_U634 ( .A(DP_mult_209_n1387), .B(DP_mult_209_n1211), .CI(
        DP_mult_209_n1233), .CO(DP_mult_209_n854), .S(DP_mult_209_n855) );
  FA_X1 DP_mult_209_U633 ( .A(DP_mult_209_n1255), .B(DP_mult_209_n1321), .CI(
        DP_mult_209_n874), .CO(DP_mult_209_n852), .S(DP_mult_209_n853) );
  FA_X1 DP_mult_209_U632 ( .A(DP_mult_209_n1299), .B(DP_mult_209_n1277), .CI(
        DP_mult_209_n1343), .CO(DP_mult_209_n850), .S(DP_mult_209_n851) );
  FA_X1 DP_mult_209_U631 ( .A(DP_mult_209_n1410), .B(DP_mult_209_n1365), .CI(
        DP_mult_209_n872), .CO(DP_mult_209_n848), .S(DP_mult_209_n849) );
  FA_X1 DP_mult_209_U630 ( .A(DP_mult_209_n868), .B(DP_mult_209_n870), .CI(
        DP_mult_209_n851), .CO(DP_mult_209_n846), .S(DP_mult_209_n847) );
  FA_X1 DP_mult_209_U629 ( .A(DP_mult_209_n855), .B(DP_mult_209_n853), .CI(
        DP_mult_209_n866), .CO(DP_mult_209_n844), .S(DP_mult_209_n845) );
  FA_X1 DP_mult_209_U627 ( .A(DP_mult_209_n845), .B(DP_mult_209_n847), .CI(
        DP_mult_209_n860), .CO(DP_mult_209_n840), .S(DP_mult_209_n841) );
  FA_X1 DP_mult_209_U626 ( .A(DP_mult_209_n858), .B(DP_mult_209_n843), .CI(
        DP_mult_209_n841), .CO(DP_mult_209_n838), .S(DP_mult_209_n839) );
  FA_X1 DP_mult_209_U623 ( .A(DP_mult_209_n1232), .B(DP_mult_209_n1364), .CI(
        DP_mult_209_n1342), .CO(DP_mult_209_n832), .S(DP_mult_209_n833) );
  FA_X1 DP_mult_209_U622 ( .A(DP_mult_209_n1320), .B(DP_mult_209_n1254), .CI(
        DP_mult_209_n1298), .CO(DP_mult_209_n830), .S(DP_mult_209_n831) );
  FA_X1 DP_mult_209_U621 ( .A(DP_mult_209_n852), .B(DP_mult_209_n854), .CI(
        DP_mult_209_n850), .CO(DP_mult_209_n828), .S(DP_mult_209_n829) );
  FA_X1 DP_mult_209_U620 ( .A(DP_mult_209_n835), .B(DP_mult_209_n831), .CI(
        DP_mult_209_n833), .CO(DP_mult_209_n826), .S(DP_mult_209_n827) );
  FA_X1 DP_mult_209_U619 ( .A(DP_mult_209_n846), .B(DP_mult_209_n848), .CI(
        DP_mult_209_n829), .CO(DP_mult_209_n824), .S(DP_mult_209_n825) );
  FA_X1 DP_mult_209_U617 ( .A(DP_mult_209_n840), .B(DP_mult_209_n825), .CI(
        DP_mult_209_n823), .CO(DP_mult_209_n820), .S(DP_mult_209_n821) );
  FA_X1 DP_mult_209_U616 ( .A(DP_mult_209_n836), .B(DP_mult_209_n1209), .CI(
        DP_mult_209_n1363), .CO(DP_mult_209_n818), .S(DP_mult_209_n819) );
  FA_X1 DP_mult_209_U615 ( .A(DP_mult_209_n1231), .B(DP_mult_209_n1297), .CI(
        DP_mult_209_n1275), .CO(DP_mult_209_n816), .S(DP_mult_209_n817) );
  FA_X1 DP_mult_209_U614 ( .A(DP_mult_209_n1319), .B(DP_mult_209_n1253), .CI(
        DP_mult_209_n1341), .CO(DP_mult_209_n814), .S(DP_mult_209_n815) );
  FA_X1 DP_mult_209_U613 ( .A(DP_mult_209_n834), .B(DP_mult_209_n1386), .CI(
        DP_mult_209_n830), .CO(DP_mult_209_n812), .S(DP_mult_209_n813) );
  FA_X1 DP_mult_209_U612 ( .A(DP_mult_209_n815), .B(DP_mult_209_n832), .CI(
        DP_mult_209_n817), .CO(DP_mult_209_n810), .S(DP_mult_209_n811) );
  FA_X1 DP_mult_209_U611 ( .A(DP_mult_209_n828), .B(DP_mult_209_n819), .CI(
        DP_mult_209_n813), .CO(DP_mult_209_n808), .S(DP_mult_209_n809) );
  FA_X1 DP_mult_209_U610 ( .A(DP_mult_209_n811), .B(DP_mult_209_n826), .CI(
        DP_mult_209_n824), .CO(DP_mult_209_n806), .S(DP_mult_209_n807) );
  FA_X1 DP_mult_209_U609 ( .A(DP_mult_209_n822), .B(DP_mult_209_n809), .CI(
        DP_mult_209_n807), .CO(DP_mult_209_n804), .S(DP_mult_209_n805) );
  FA_X1 DP_mult_209_U607 ( .A(DP_mult_209_n1340), .B(DP_mult_209_n1252), .CI(
        DP_mult_209_n803), .CO(DP_mult_209_n800), .S(DP_mult_209_n801) );
  FA_X1 DP_mult_209_U606 ( .A(DP_mult_209_n1208), .B(DP_mult_209_n1318), .CI(
        DP_mult_209_n1230), .CO(DP_mult_209_n798), .S(DP_mult_209_n799) );
  FA_X1 DP_mult_209_U605 ( .A(DP_mult_209_n1274), .B(DP_mult_209_n1296), .CI(
        DP_mult_209_n818), .CO(DP_mult_209_n796), .S(DP_mult_209_n797) );
  FA_X1 DP_mult_209_U604 ( .A(DP_mult_209_n814), .B(DP_mult_209_n816), .CI(
        DP_mult_209_n799), .CO(DP_mult_209_n794), .S(DP_mult_209_n795) );
  FA_X1 DP_mult_209_U603 ( .A(DP_mult_209_n812), .B(DP_mult_209_n801), .CI(
        DP_mult_209_n797), .CO(DP_mult_209_n792), .S(DP_mult_209_n793) );
  FA_X1 DP_mult_209_U602 ( .A(DP_mult_209_n795), .B(DP_mult_209_n810), .CI(
        DP_mult_209_n808), .CO(DP_mult_209_n790), .S(DP_mult_209_n791) );
  FA_X1 DP_mult_209_U601 ( .A(DP_mult_209_n806), .B(DP_mult_209_n793), .CI(
        DP_mult_209_n791), .CO(DP_mult_209_n788), .S(DP_mult_209_n789) );
  FA_X1 DP_mult_209_U600 ( .A(DP_mult_209_n802), .B(DP_mult_209_n1207), .CI(
        DP_mult_209_n1251), .CO(DP_mult_209_n786), .S(DP_mult_209_n787) );
  FA_X1 DP_mult_209_U599 ( .A(DP_mult_209_n1273), .B(DP_mult_209_n1317), .CI(
        DP_mult_209_n1295), .CO(DP_mult_209_n784), .S(DP_mult_209_n785) );
  FA_X1 DP_mult_209_U598 ( .A(DP_mult_209_n1339), .B(DP_mult_209_n1229), .CI(
        DP_mult_209_n1362), .CO(DP_mult_209_n782), .S(DP_mult_209_n783) );
  FA_X1 DP_mult_209_U597 ( .A(DP_mult_209_n798), .B(DP_mult_209_n800), .CI(
        DP_mult_209_n785), .CO(DP_mult_209_n780), .S(DP_mult_209_n781) );
  FA_X1 DP_mult_209_U596 ( .A(DP_mult_209_n796), .B(DP_mult_209_n787), .CI(
        DP_mult_209_n783), .CO(DP_mult_209_n778), .S(DP_mult_209_n779) );
  FA_X1 DP_mult_209_U595 ( .A(DP_mult_209_n781), .B(DP_mult_209_n794), .CI(
        DP_mult_209_n792), .CO(DP_mult_209_n776), .S(DP_mult_209_n777) );
  FA_X1 DP_mult_209_U594 ( .A(DP_mult_209_n790), .B(DP_mult_209_n779), .CI(
        DP_mult_209_n777), .CO(DP_mult_209_n774), .S(DP_mult_209_n775) );
  FA_X1 DP_mult_209_U592 ( .A(DP_mult_209_n1316), .B(DP_mult_209_n1250), .CI(
        DP_mult_209_n773), .CO(DP_mult_209_n770), .S(DP_mult_209_n771) );
  FA_X1 DP_mult_209_U591 ( .A(DP_mult_209_n1294), .B(DP_mult_209_n1206), .CI(
        DP_mult_209_n1272), .CO(DP_mult_209_n768), .S(DP_mult_209_n769) );
  FA_X1 DP_mult_209_U590 ( .A(DP_mult_209_n786), .B(DP_mult_209_n1228), .CI(
        DP_mult_209_n784), .CO(DP_mult_209_n766), .S(DP_mult_209_n767) );
  FA_X1 DP_mult_209_U589 ( .A(DP_mult_209_n771), .B(DP_mult_209_n769), .CI(
        DP_mult_209_n782), .CO(DP_mult_209_n764), .S(DP_mult_209_n765) );
  FA_X1 DP_mult_209_U588 ( .A(DP_mult_209_n767), .B(DP_mult_209_n780), .CI(
        DP_mult_209_n778), .CO(DP_mult_209_n762), .S(DP_mult_209_n763) );
  FA_X1 DP_mult_209_U587 ( .A(DP_mult_209_n776), .B(DP_mult_209_n765), .CI(
        DP_mult_209_n763), .CO(DP_mult_209_n760), .S(DP_mult_209_n761) );
  FA_X1 DP_mult_209_U586 ( .A(DP_mult_209_n772), .B(DP_mult_209_n1205), .CI(
        DP_mult_209_n1227), .CO(DP_mult_209_n758), .S(DP_mult_209_n759) );
  FA_X1 DP_mult_209_U585 ( .A(DP_mult_209_n1249), .B(DP_mult_209_n1293), .CI(
        DP_mult_209_n1315), .CO(DP_mult_209_n756), .S(DP_mult_209_n757) );
  FA_X1 DP_mult_209_U584 ( .A(DP_mult_209_n1338), .B(DP_mult_209_n1271), .CI(
        DP_mult_209_n770), .CO(DP_mult_209_n754), .S(DP_mult_209_n755) );
  FA_X1 DP_mult_209_U583 ( .A(DP_mult_209_n757), .B(DP_mult_209_n768), .CI(
        DP_mult_209_n759), .CO(DP_mult_209_n752), .S(DP_mult_209_n753) );
  FA_X1 DP_mult_209_U582 ( .A(DP_mult_209_n755), .B(DP_mult_209_n766), .CI(
        DP_mult_209_n764), .CO(DP_mult_209_n750), .S(DP_mult_209_n751) );
  FA_X1 DP_mult_209_U581 ( .A(DP_mult_209_n762), .B(DP_mult_209_n753), .CI(
        DP_mult_209_n751), .CO(DP_mult_209_n748), .S(DP_mult_209_n749) );
  FA_X1 DP_mult_209_U579 ( .A(DP_mult_209_n1292), .B(DP_mult_209_n1248), .CI(
        DP_mult_209_n747), .CO(DP_mult_209_n744), .S(DP_mult_209_n745) );
  FA_X1 DP_mult_209_U578 ( .A(DP_mult_209_n1226), .B(DP_mult_209_n1204), .CI(
        DP_mult_209_n1270), .CO(DP_mult_209_n742), .S(DP_mult_209_n743) );
  FA_X1 DP_mult_209_U577 ( .A(DP_mult_209_n756), .B(DP_mult_209_n758), .CI(
        DP_mult_209_n743), .CO(DP_mult_209_n740), .S(DP_mult_209_n741) );
  FA_X1 DP_mult_209_U576 ( .A(DP_mult_209_n754), .B(DP_mult_209_n745), .CI(
        DP_mult_209_n752), .CO(DP_mult_209_n738), .S(DP_mult_209_n739) );
  FA_X1 DP_mult_209_U575 ( .A(DP_mult_209_n750), .B(DP_mult_209_n741), .CI(
        DP_mult_209_n739), .CO(DP_mult_209_n736), .S(DP_mult_209_n737) );
  FA_X1 DP_mult_209_U574 ( .A(DP_mult_209_n746), .B(DP_mult_209_n1203), .CI(
        DP_mult_209_n1247), .CO(DP_mult_209_n734), .S(DP_mult_209_n735) );
  FA_X1 DP_mult_209_U573 ( .A(DP_mult_209_n1225), .B(DP_mult_209_n1291), .CI(
        DP_mult_209_n1269), .CO(DP_mult_209_n732), .S(DP_mult_209_n733) );
  FA_X1 DP_mult_209_U572 ( .A(DP_mult_209_n744), .B(DP_mult_209_n1314), .CI(
        DP_mult_209_n742), .CO(DP_mult_209_n730), .S(DP_mult_209_n731) );
  FA_X1 DP_mult_209_U571 ( .A(DP_mult_209_n735), .B(DP_mult_209_n733), .CI(
        DP_mult_209_n740), .CO(DP_mult_209_n728), .S(DP_mult_209_n729) );
  FA_X1 DP_mult_209_U570 ( .A(DP_mult_209_n738), .B(DP_mult_209_n731), .CI(
        DP_mult_209_n729), .CO(DP_mult_209_n726), .S(DP_mult_209_n727) );
  FA_X1 DP_mult_209_U568 ( .A(DP_mult_209_n1268), .B(DP_mult_209_n1224), .CI(
        DP_mult_209_n725), .CO(DP_mult_209_n722), .S(DP_mult_209_n723) );
  FA_X1 DP_mult_209_U567 ( .A(DP_mult_209_n1202), .B(DP_mult_209_n1246), .CI(
        DP_mult_209_n734), .CO(DP_mult_209_n720), .S(DP_mult_209_n721) );
  FA_X1 DP_mult_209_U566 ( .A(DP_mult_209_n723), .B(DP_mult_209_n732), .CI(
        DP_mult_209_n730), .CO(DP_mult_209_n718), .S(DP_mult_209_n719) );
  FA_X1 DP_mult_209_U565 ( .A(DP_mult_209_n728), .B(DP_mult_209_n721), .CI(
        DP_mult_209_n719), .CO(DP_mult_209_n716), .S(DP_mult_209_n717) );
  FA_X1 DP_mult_209_U564 ( .A(DP_mult_209_n1267), .B(DP_mult_209_n1201), .CI(
        DP_mult_209_n724), .CO(DP_mult_209_n714), .S(DP_mult_209_n715) );
  FA_X1 DP_mult_209_U563 ( .A(DP_mult_209_n1245), .B(DP_mult_209_n1223), .CI(
        DP_mult_209_n1290), .CO(DP_mult_209_n712), .S(DP_mult_209_n713) );
  FA_X1 DP_mult_209_U562 ( .A(DP_mult_209_n715), .B(DP_mult_209_n722), .CI(
        DP_mult_209_n720), .CO(DP_mult_209_n710), .S(DP_mult_209_n711) );
  FA_X1 DP_mult_209_U561 ( .A(DP_mult_209_n718), .B(DP_mult_209_n713), .CI(
        DP_mult_209_n711), .CO(DP_mult_209_n708), .S(DP_mult_209_n709) );
  FA_X1 DP_mult_209_U559 ( .A(DP_mult_209_n1222), .B(DP_mult_209_n1200), .CI(
        DP_mult_209_n707), .CO(DP_mult_209_n704), .S(DP_mult_209_n705) );
  FA_X1 DP_mult_209_U558 ( .A(DP_mult_209_n714), .B(DP_mult_209_n1244), .CI(
        DP_mult_209_n705), .CO(DP_mult_209_n702), .S(DP_mult_209_n703) );
  FA_X1 DP_mult_209_U557 ( .A(DP_mult_209_n710), .B(DP_mult_209_n712), .CI(
        DP_mult_209_n703), .CO(DP_mult_209_n700), .S(DP_mult_209_n701) );
  FA_X1 DP_mult_209_U556 ( .A(DP_mult_209_n1221), .B(DP_mult_209_n1199), .CI(
        DP_mult_209_n706), .CO(DP_mult_209_n698), .S(DP_mult_209_n699) );
  FA_X1 DP_mult_209_U555 ( .A(DP_mult_209_n1266), .B(DP_mult_209_n1243), .CI(
        DP_mult_209_n704), .CO(DP_mult_209_n696), .S(DP_mult_209_n697) );
  FA_X1 DP_mult_209_U554 ( .A(DP_mult_209_n702), .B(DP_mult_209_n699), .CI(
        DP_mult_209_n697), .CO(DP_mult_209_n694), .S(DP_mult_209_n695) );
  FA_X1 DP_mult_209_U552 ( .A(DP_mult_209_n1198), .B(DP_mult_209_n1220), .CI(
        DP_mult_209_n693), .CO(DP_mult_209_n690), .S(DP_mult_209_n691) );
  FA_X1 DP_mult_209_U551 ( .A(DP_mult_209_n691), .B(DP_mult_209_n698), .CI(
        DP_mult_209_n696), .CO(DP_mult_209_n688), .S(DP_mult_209_n689) );
  FA_X1 DP_mult_209_U550 ( .A(DP_mult_209_n1219), .B(DP_mult_209_n692), .CI(
        DP_mult_209_n1197), .CO(DP_mult_209_n686), .S(DP_mult_209_n687) );
  FA_X1 DP_mult_209_U549 ( .A(DP_mult_209_n690), .B(DP_mult_209_n1242), .CI(
        DP_mult_209_n687), .CO(DP_mult_209_n684), .S(DP_mult_209_n685) );
  FA_X1 DP_mult_209_U547 ( .A(DP_mult_209_n683), .B(DP_mult_209_n1196), .CI(
        DP_mult_209_n686), .CO(DP_mult_209_n680), .S(DP_mult_209_n681) );
  FA_X1 DP_mult_209_U546 ( .A(DP_mult_209_n1195), .B(DP_mult_209_n682), .CI(
        DP_mult_209_n1218), .CO(DP_mult_209_n678), .S(DP_mult_209_n679) );
  XNOR2_X1 CU_U5 ( .A(vIn), .B(CU_n3), .ZN(CU_nextState_0_) );
  INV_X1 CU_U4 ( .A(CU_n3), .ZN(sw_regs_en_int) );
  XNOR2_X1 CU_U3 ( .A(CU_n1), .B(CU_n2), .ZN(CU_n3) );
  DFFR_X1 CU_presentState_reg_1_ ( .D(sw_regs_en_int), .CK(clk), .RN(rst_n), 
        .Q(delayed_controls_0__1_), .QN(CU_n2) );
  DFFR_X1 CU_presentState_reg_0_ ( .D(CU_nextState_0_), .CK(clk), .RN(rst_n), 
        .QN(CU_n1) );
  MUX2_X1 reg_delay_0_U3 ( .A(delayed_controls_1__0_), .B(sw_regs_en_int), .S(
        1'b1), .Z(reg_delay_0_n6) );
  MUX2_X1 reg_delay_0_U2 ( .A(delayed_controls_1__1_), .B(
        delayed_controls_0__1_), .S(1'b1), .Z(reg_delay_0_n5) );
  DFFR_X1 reg_delay_0_Q_reg_1_ ( .D(reg_delay_0_n6), .CK(clk), .RN(rst_n), .Q(
        delayed_controls_1__0_) );
  DFFR_X1 reg_delay_0_Q_reg_0_ ( .D(reg_delay_0_n5), .CK(clk), .RN(rst_n), .Q(
        delayed_controls_1__1_) );
  MUX2_X1 reg_delay_1_U3 ( .A(delayed_controls_2__0_), .B(
        delayed_controls_1__0_), .S(1'b1), .Z(reg_delay_1_n3) );
  MUX2_X1 reg_delay_1_U2 ( .A(vOut), .B(delayed_controls_1__1_), .S(1'b1), .Z(
        reg_delay_1_n4) );
  DFFR_X1 reg_delay_1_Q_reg_0_ ( .D(reg_delay_1_n4), .CK(clk), .RN(rst_n), .Q(
        vOut) );
  DFFR_X1 reg_delay_1_Q_reg_1_ ( .D(reg_delay_1_n3), .CK(clk), .RN(rst_n), .Q(
        delayed_controls_2__0_) );
endmodule

