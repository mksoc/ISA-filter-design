
module iir_filter ( clk, rst_n, vIn, dIn, a, b, dOut, vOut );
  input [11:0] dIn;
  input [23:0] a;
  input [35:0] b;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   sw_out_regs_en_int, DP_n17, DP_n16, DP_n15, DP_n14, DP_n13, DP_n12,
         DP_n11, DP_n10, DP_n9, DP_n8, DP_n7, DP_n6, DP_n5, DP_n4, DP_n3,
         DP_n2, DP_n1, DP_fb_0_, DP_fb_10_, DP_fb_11_, DP_fb_12_, DP_fb_1_,
         DP_fb_2_, DP_fb_3_, DP_fb_4_, DP_fb_5_, DP_fb_6_, DP_fb_7_, DP_fb_8_,
         DP_fb_9_, DP_ff_0_, DP_ff_10_, DP_ff_11_, DP_ff_12_, DP_ff_1_,
         DP_ff_2_, DP_ff_3_, DP_ff_4_, DP_ff_5_, DP_ff_6_, DP_ff_7_, DP_ff_8_,
         DP_ff_9_, DP_w_b0_0_, DP_w_b0_1_, DP_w_b0_2_, DP_w_b0_3_, DP_w_b0_4_,
         DP_w_b0_5_, DP_w_b0_6_, DP_w_b0_7_, DP_w_b0_8_, DP_w_b0_9_,
         DP_w_b0_10_, DP_w_b0_11_, DP_sw1_b2_0_, DP_sw1_b2_1_, DP_sw1_b2_2_,
         DP_sw1_b2_3_, DP_sw1_b2_4_, DP_sw1_b2_5_, DP_sw1_b2_6_, DP_sw1_b2_7_,
         DP_sw1_b2_8_, DP_sw1_b2_9_, DP_sw1_b2_10_, DP_sw1_b2_11_,
         DP_sw0_b1_0_, DP_sw0_b1_1_, DP_sw0_b1_2_, DP_sw0_b1_3_, DP_sw0_b1_4_,
         DP_sw0_b1_5_, DP_sw0_b1_6_, DP_sw0_b1_7_, DP_sw0_b1_8_, DP_sw0_b1_9_,
         DP_sw0_b1_10_, DP_sw0_b1_11_, DP_sw1_a2_0_, DP_sw1_a2_1_,
         DP_sw1_a2_2_, DP_sw1_a2_3_, DP_sw1_a2_4_, DP_sw1_a2_5_, DP_sw1_a2_6_,
         DP_sw1_a2_7_, DP_sw1_a2_8_, DP_sw1_a2_9_, DP_sw1_a2_10_,
         DP_sw1_a2_11_, DP_sw0_a1_0_, DP_sw0_a1_1_, DP_sw0_a1_2_, DP_sw0_a1_3_,
         DP_sw0_a1_4_, DP_sw0_a1_5_, DP_sw0_a1_6_, DP_sw0_a1_7_, DP_sw0_a1_8_,
         DP_sw0_a1_9_, DP_sw0_a1_10_, DP_sw0_a1_11_, DP_y_out_0_, DP_y_out_1_,
         DP_y_out_2_, DP_y_out_3_, DP_y_out_4_, DP_y_out_5_, DP_y_out_6_,
         DP_y_out_7_, DP_y_out_8_, DP_y_out_9_, DP_y_out_10_, DP_y_out_11_,
         DP_sw1_0_, DP_sw1_1_, DP_sw1_2_, DP_sw1_3_, DP_sw1_4_, DP_sw1_5_,
         DP_sw1_6_, DP_sw1_7_, DP_sw1_8_, DP_sw1_9_, DP_sw1_10_, DP_sw1_11_,
         DP_sw1_12_, DP_sw0_0_, DP_sw0_1_, DP_sw0_2_, DP_sw0_3_, DP_sw0_4_,
         DP_sw0_5_, DP_sw0_6_, DP_sw0_7_, DP_sw0_8_, DP_sw0_9_, DP_sw0_10_,
         DP_sw0_11_, DP_sw0_12_, DP_w_0_, DP_w_1_, DP_w_2_, DP_w_3_, DP_w_4_,
         DP_w_5_, DP_w_6_, DP_w_7_, DP_w_8_, DP_w_9_, DP_w_10_, DP_w_11_,
         DP_w_12_, DP_x_0_, DP_x_1_, DP_x_2_, DP_x_3_, DP_x_4_, DP_x_5_,
         DP_x_6_, DP_x_7_, DP_x_8_, DP_x_9_, DP_x_10_, DP_x_11_, DP_reg_in_n39,
         DP_reg_in_n38, DP_reg_in_n37, DP_reg_in_n36, DP_reg_in_n35,
         DP_reg_in_n34, DP_reg_in_n33, DP_reg_in_n32, DP_reg_in_n31,
         DP_reg_in_n30, DP_reg_in_n29, DP_reg_in_n28, DP_reg_in_n27,
         DP_reg_in_n26, DP_reg_in_n25, DP_reg_in_n24, DP_reg_in_n23,
         DP_reg_in_n22, DP_reg_in_n21, DP_reg_in_n20, DP_reg_in_n19,
         DP_reg_in_n18, DP_reg_in_n17, DP_reg_in_n16, DP_reg_in_n15,
         DP_reg_in_n14, DP_reg_in_n13, DP_reg_in_n12, DP_reg_in_n11,
         DP_reg_in_n10, DP_reg_in_n9, DP_reg_in_n8, DP_reg_in_n7, DP_reg_in_n6,
         DP_reg_in_n5, DP_reg_in_n4, DP_reg_in_n3, DP_reg_in_n2, DP_reg_in_n1,
         DP_reg_a_i_1_n74, DP_reg_a_i_1_n73, DP_reg_a_i_1_n72,
         DP_reg_a_i_1_n71, DP_reg_a_i_1_n70, DP_reg_a_i_1_n69,
         DP_reg_a_i_1_n68, DP_reg_a_i_1_n67, DP_reg_a_i_1_n66,
         DP_reg_a_i_1_n65, DP_reg_a_i_1_n64, DP_reg_a_i_1_n63,
         DP_reg_a_i_1_n62, DP_reg_a_i_1_n61, DP_reg_a_i_1_n60,
         DP_reg_a_i_1_n59, DP_reg_a_i_1_n58, DP_reg_a_i_1_n57,
         DP_reg_a_i_1_n56, DP_reg_a_i_1_n55, DP_reg_a_i_1_n54,
         DP_reg_a_i_1_n53, DP_reg_a_i_1_n52, DP_reg_a_i_1_n51,
         DP_reg_a_i_1_n50, DP_reg_a_i_1_n49, DP_reg_a_i_1_n48,
         DP_reg_a_i_1_n47, DP_reg_a_i_1_n46, DP_reg_a_i_1_n45,
         DP_reg_a_i_1_n44, DP_reg_a_i_1_n43, DP_reg_a_i_1_n42,
         DP_reg_a_i_1_n41, DP_reg_a_i_1_n40, DP_reg_a_i_1_n39,
         DP_reg_a_i_1_n38, DP_reg_a_i_1_n37, DP_reg_a_i_2_n74,
         DP_reg_a_i_2_n73, DP_reg_a_i_2_n72, DP_reg_a_i_2_n71,
         DP_reg_a_i_2_n70, DP_reg_a_i_2_n69, DP_reg_a_i_2_n68,
         DP_reg_a_i_2_n67, DP_reg_a_i_2_n66, DP_reg_a_i_2_n65,
         DP_reg_a_i_2_n64, DP_reg_a_i_2_n63, DP_reg_a_i_2_n62,
         DP_reg_a_i_2_n61, DP_reg_a_i_2_n60, DP_reg_a_i_2_n59,
         DP_reg_a_i_2_n58, DP_reg_a_i_2_n57, DP_reg_a_i_2_n56,
         DP_reg_a_i_2_n55, DP_reg_a_i_2_n54, DP_reg_a_i_2_n53,
         DP_reg_a_i_2_n52, DP_reg_a_i_2_n51, DP_reg_a_i_2_n50,
         DP_reg_a_i_2_n49, DP_reg_a_i_2_n48, DP_reg_a_i_2_n47,
         DP_reg_a_i_2_n46, DP_reg_a_i_2_n45, DP_reg_a_i_2_n44,
         DP_reg_a_i_2_n43, DP_reg_a_i_2_n42, DP_reg_a_i_2_n41,
         DP_reg_a_i_2_n40, DP_reg_a_i_2_n39, DP_reg_a_i_2_n38,
         DP_reg_a_i_2_n37, DP_reg_b_i_0_n74, DP_reg_b_i_0_n73,
         DP_reg_b_i_0_n72, DP_reg_b_i_0_n71, DP_reg_b_i_0_n70,
         DP_reg_b_i_0_n69, DP_reg_b_i_0_n68, DP_reg_b_i_0_n67,
         DP_reg_b_i_0_n66, DP_reg_b_i_0_n65, DP_reg_b_i_0_n64,
         DP_reg_b_i_0_n63, DP_reg_b_i_0_n62, DP_reg_b_i_0_n61,
         DP_reg_b_i_0_n60, DP_reg_b_i_0_n59, DP_reg_b_i_0_n58,
         DP_reg_b_i_0_n57, DP_reg_b_i_0_n56, DP_reg_b_i_0_n55,
         DP_reg_b_i_0_n54, DP_reg_b_i_0_n53, DP_reg_b_i_0_n52,
         DP_reg_b_i_0_n51, DP_reg_b_i_0_n50, DP_reg_b_i_0_n49,
         DP_reg_b_i_0_n48, DP_reg_b_i_0_n47, DP_reg_b_i_0_n46,
         DP_reg_b_i_0_n45, DP_reg_b_i_0_n44, DP_reg_b_i_0_n43,
         DP_reg_b_i_0_n42, DP_reg_b_i_0_n41, DP_reg_b_i_0_n40,
         DP_reg_b_i_0_n39, DP_reg_b_i_0_n38, DP_reg_b_i_0_n37,
         DP_reg_b_i_1_n74, DP_reg_b_i_1_n73, DP_reg_b_i_1_n72,
         DP_reg_b_i_1_n71, DP_reg_b_i_1_n70, DP_reg_b_i_1_n69,
         DP_reg_b_i_1_n68, DP_reg_b_i_1_n67, DP_reg_b_i_1_n66,
         DP_reg_b_i_1_n65, DP_reg_b_i_1_n64, DP_reg_b_i_1_n63,
         DP_reg_b_i_1_n62, DP_reg_b_i_1_n61, DP_reg_b_i_1_n60,
         DP_reg_b_i_1_n59, DP_reg_b_i_1_n58, DP_reg_b_i_1_n57,
         DP_reg_b_i_1_n56, DP_reg_b_i_1_n55, DP_reg_b_i_1_n54,
         DP_reg_b_i_1_n53, DP_reg_b_i_1_n52, DP_reg_b_i_1_n51,
         DP_reg_b_i_1_n50, DP_reg_b_i_1_n49, DP_reg_b_i_1_n48,
         DP_reg_b_i_1_n47, DP_reg_b_i_1_n46, DP_reg_b_i_1_n45,
         DP_reg_b_i_1_n44, DP_reg_b_i_1_n43, DP_reg_b_i_1_n42,
         DP_reg_b_i_1_n41, DP_reg_b_i_1_n40, DP_reg_b_i_1_n39,
         DP_reg_b_i_1_n38, DP_reg_b_i_1_n37, DP_reg_b_i_2_n74,
         DP_reg_b_i_2_n73, DP_reg_b_i_2_n72, DP_reg_b_i_2_n71,
         DP_reg_b_i_2_n70, DP_reg_b_i_2_n69, DP_reg_b_i_2_n68,
         DP_reg_b_i_2_n67, DP_reg_b_i_2_n66, DP_reg_b_i_2_n65,
         DP_reg_b_i_2_n64, DP_reg_b_i_2_n63, DP_reg_b_i_2_n62,
         DP_reg_b_i_2_n61, DP_reg_b_i_2_n60, DP_reg_b_i_2_n59,
         DP_reg_b_i_2_n58, DP_reg_b_i_2_n57, DP_reg_b_i_2_n56,
         DP_reg_b_i_2_n55, DP_reg_b_i_2_n54, DP_reg_b_i_2_n53,
         DP_reg_b_i_2_n52, DP_reg_b_i_2_n51, DP_reg_b_i_2_n50,
         DP_reg_b_i_2_n49, DP_reg_b_i_2_n48, DP_reg_b_i_2_n47,
         DP_reg_b_i_2_n46, DP_reg_b_i_2_n45, DP_reg_b_i_2_n44,
         DP_reg_b_i_2_n43, DP_reg_b_i_2_n42, DP_reg_b_i_2_n41,
         DP_reg_b_i_2_n40, DP_reg_b_i_2_n39, DP_reg_b_i_2_n38,
         DP_reg_b_i_2_n37, DP_reg_sw0_n42, DP_reg_sw0_n41, DP_reg_sw0_n40,
         DP_reg_sw0_n39, DP_reg_sw0_n38, DP_reg_sw0_n37, DP_reg_sw0_n36,
         DP_reg_sw0_n35, DP_reg_sw0_n34, DP_reg_sw0_n33, DP_reg_sw0_n32,
         DP_reg_sw0_n31, DP_reg_sw0_n30, DP_reg_sw0_n29, DP_reg_sw0_n28,
         DP_reg_sw0_n27, DP_reg_sw0_n26, DP_reg_sw0_n25, DP_reg_sw0_n24,
         DP_reg_sw0_n23, DP_reg_sw0_n22, DP_reg_sw0_n21, DP_reg_sw0_n20,
         DP_reg_sw0_n19, DP_reg_sw0_n18, DP_reg_sw0_n17, DP_reg_sw0_n16,
         DP_reg_sw0_n15, DP_reg_sw0_n14, DP_reg_sw0_n13, DP_reg_sw0_n12,
         DP_reg_sw0_n11, DP_reg_sw0_n10, DP_reg_sw0_n9, DP_reg_sw0_n8,
         DP_reg_sw0_n7, DP_reg_sw0_n6, DP_reg_sw0_n5, DP_reg_sw0_n4,
         DP_reg_sw0_n3, DP_reg_sw0_n2, DP_reg_sw0_n1, DP_reg_sw1_n80,
         DP_reg_sw1_n79, DP_reg_sw1_n78, DP_reg_sw1_n77, DP_reg_sw1_n76,
         DP_reg_sw1_n75, DP_reg_sw1_n74, DP_reg_sw1_n73, DP_reg_sw1_n72,
         DP_reg_sw1_n71, DP_reg_sw1_n70, DP_reg_sw1_n69, DP_reg_sw1_n68,
         DP_reg_sw1_n67, DP_reg_sw1_n66, DP_reg_sw1_n65, DP_reg_sw1_n64,
         DP_reg_sw1_n63, DP_reg_sw1_n62, DP_reg_sw1_n61, DP_reg_sw1_n60,
         DP_reg_sw1_n59, DP_reg_sw1_n58, DP_reg_sw1_n57, DP_reg_sw1_n56,
         DP_reg_sw1_n55, DP_reg_sw1_n54, DP_reg_sw1_n53, DP_reg_sw1_n52,
         DP_reg_sw1_n51, DP_reg_sw1_n50, DP_reg_sw1_n49, DP_reg_sw1_n48,
         DP_reg_sw1_n47, DP_reg_sw1_n46, DP_reg_sw1_n45, DP_reg_sw1_n44,
         DP_reg_sw1_n43, DP_reg_sw1_n42, DP_reg_sw1_n41, DP_reg_sw1_n40,
         DP_reg_out_n74, DP_reg_out_n73, DP_reg_out_n72, DP_reg_out_n71,
         DP_reg_out_n70, DP_reg_out_n69, DP_reg_out_n68, DP_reg_out_n67,
         DP_reg_out_n66, DP_reg_out_n65, DP_reg_out_n64, DP_reg_out_n63,
         DP_reg_out_n62, DP_reg_out_n61, DP_reg_out_n60, DP_reg_out_n59,
         DP_reg_out_n58, DP_reg_out_n57, DP_reg_out_n56, DP_reg_out_n55,
         DP_reg_out_n54, DP_reg_out_n53, DP_reg_out_n52, DP_reg_out_n51,
         DP_reg_out_n50, DP_reg_out_n49, DP_reg_out_n48, DP_reg_out_n47,
         DP_reg_out_n46, DP_reg_out_n45, DP_reg_out_n44, DP_reg_out_n43,
         DP_reg_out_n42, DP_reg_out_n41, DP_reg_out_n40, DP_reg_out_n39,
         DP_reg_out_n38, DP_reg_out_n37,
         DP_add_1_root_add_0_root_add_107_carry_1_,
         DP_add_1_root_add_0_root_add_107_carry_2_,
         DP_add_1_root_add_0_root_add_107_carry_3_,
         DP_add_1_root_add_0_root_add_107_carry_4_,
         DP_add_1_root_add_0_root_add_107_carry_5_,
         DP_add_1_root_add_0_root_add_107_carry_6_,
         DP_add_1_root_add_0_root_add_107_carry_7_,
         DP_add_1_root_add_0_root_add_107_carry_8_,
         DP_add_1_root_add_0_root_add_107_carry_9_,
         DP_add_1_root_add_0_root_add_107_carry_10_,
         DP_add_1_root_add_0_root_add_107_carry_11_,
         DP_add_1_root_add_0_root_add_107_carry_12_,
         DP_add_0_root_add_0_root_add_107_carry_1_,
         DP_add_0_root_add_0_root_add_107_carry_2_,
         DP_add_0_root_add_0_root_add_107_carry_3_,
         DP_add_0_root_add_0_root_add_107_carry_4_,
         DP_add_0_root_add_0_root_add_107_carry_5_,
         DP_add_0_root_add_0_root_add_107_carry_6_,
         DP_add_0_root_add_0_root_add_107_carry_7_,
         DP_add_0_root_add_0_root_add_107_carry_8_,
         DP_add_0_root_add_0_root_add_107_carry_9_,
         DP_add_0_root_add_0_root_add_107_carry_10_,
         DP_add_0_root_add_0_root_add_107_carry_11_,
         DP_add_0_root_add_0_root_add_107_carry_12_, DP_mult_105_n660,
         DP_mult_105_n659, DP_mult_105_n658, DP_mult_105_n657,
         DP_mult_105_n656, DP_mult_105_n655, DP_mult_105_n654,
         DP_mult_105_n653, DP_mult_105_n652, DP_mult_105_n651,
         DP_mult_105_n650, DP_mult_105_n649, DP_mult_105_n648,
         DP_mult_105_n647, DP_mult_105_n646, DP_mult_105_n645,
         DP_mult_105_n644, DP_mult_105_n643, DP_mult_105_n642,
         DP_mult_105_n641, DP_mult_105_n640, DP_mult_105_n639,
         DP_mult_105_n638, DP_mult_105_n637, DP_mult_105_n636,
         DP_mult_105_n635, DP_mult_105_n634, DP_mult_105_n633,
         DP_mult_105_n632, DP_mult_105_n631, DP_mult_105_n630,
         DP_mult_105_n629, DP_mult_105_n628, DP_mult_105_n627,
         DP_mult_105_n626, DP_mult_105_n625, DP_mult_105_n624,
         DP_mult_105_n623, DP_mult_105_n622, DP_mult_105_n621,
         DP_mult_105_n620, DP_mult_105_n619, DP_mult_105_n618,
         DP_mult_105_n617, DP_mult_105_n616, DP_mult_105_n615,
         DP_mult_105_n614, DP_mult_105_n613, DP_mult_105_n612,
         DP_mult_105_n611, DP_mult_105_n610, DP_mult_105_n609,
         DP_mult_105_n608, DP_mult_105_n607, DP_mult_105_n606,
         DP_mult_105_n605, DP_mult_105_n604, DP_mult_105_n603,
         DP_mult_105_n602, DP_mult_105_n601, DP_mult_105_n600,
         DP_mult_105_n599, DP_mult_105_n598, DP_mult_105_n597,
         DP_mult_105_n596, DP_mult_105_n595, DP_mult_105_n594,
         DP_mult_105_n593, DP_mult_105_n592, DP_mult_105_n591,
         DP_mult_105_n590, DP_mult_105_n589, DP_mult_105_n588,
         DP_mult_105_n587, DP_mult_105_n586, DP_mult_105_n585,
         DP_mult_105_n584, DP_mult_105_n583, DP_mult_105_n582,
         DP_mult_105_n581, DP_mult_105_n580, DP_mult_105_n579,
         DP_mult_105_n578, DP_mult_105_n577, DP_mult_105_n576,
         DP_mult_105_n575, DP_mult_105_n574, DP_mult_105_n573,
         DP_mult_105_n572, DP_mult_105_n571, DP_mult_105_n570,
         DP_mult_105_n569, DP_mult_105_n568, DP_mult_105_n567,
         DP_mult_105_n566, DP_mult_105_n565, DP_mult_105_n564,
         DP_mult_105_n563, DP_mult_105_n562, DP_mult_105_n561,
         DP_mult_105_n560, DP_mult_105_n559, DP_mult_105_n558,
         DP_mult_105_n557, DP_mult_105_n556, DP_mult_105_n555,
         DP_mult_105_n554, DP_mult_105_n553, DP_mult_105_n552,
         DP_mult_105_n551, DP_mult_105_n550, DP_mult_105_n549,
         DP_mult_105_n548, DP_mult_105_n547, DP_mult_105_n546,
         DP_mult_105_n545, DP_mult_105_n544, DP_mult_105_n543,
         DP_mult_105_n542, DP_mult_105_n541, DP_mult_105_n540,
         DP_mult_105_n539, DP_mult_105_n538, DP_mult_105_n537,
         DP_mult_105_n536, DP_mult_105_n535, DP_mult_105_n534,
         DP_mult_105_n533, DP_mult_105_n532, DP_mult_105_n531,
         DP_mult_105_n530, DP_mult_105_n529, DP_mult_105_n528,
         DP_mult_105_n527, DP_mult_105_n526, DP_mult_105_n525,
         DP_mult_105_n524, DP_mult_105_n523, DP_mult_105_n522,
         DP_mult_105_n521, DP_mult_105_n520, DP_mult_105_n519,
         DP_mult_105_n337, DP_mult_105_n336, DP_mult_105_n335,
         DP_mult_105_n334, DP_mult_105_n333, DP_mult_105_n332,
         DP_mult_105_n331, DP_mult_105_n330, DP_mult_105_n329,
         DP_mult_105_n328, DP_mult_105_n327, DP_mult_105_n325,
         DP_mult_105_n324, DP_mult_105_n323, DP_mult_105_n322,
         DP_mult_105_n321, DP_mult_105_n320, DP_mult_105_n319,
         DP_mult_105_n318, DP_mult_105_n317, DP_mult_105_n316,
         DP_mult_105_n315, DP_mult_105_n314, DP_mult_105_n313,
         DP_mult_105_n312, DP_mult_105_n311, DP_mult_105_n310,
         DP_mult_105_n309, DP_mult_105_n308, DP_mult_105_n307,
         DP_mult_105_n306, DP_mult_105_n305, DP_mult_105_n303,
         DP_mult_105_n302, DP_mult_105_n301, DP_mult_105_n300,
         DP_mult_105_n299, DP_mult_105_n298, DP_mult_105_n297,
         DP_mult_105_n296, DP_mult_105_n295, DP_mult_105_n294,
         DP_mult_105_n293, DP_mult_105_n292, DP_mult_105_n291,
         DP_mult_105_n290, DP_mult_105_n289, DP_mult_105_n288,
         DP_mult_105_n287, DP_mult_105_n286, DP_mult_105_n285,
         DP_mult_105_n284, DP_mult_105_n283, DP_mult_105_n281,
         DP_mult_105_n280, DP_mult_105_n279, DP_mult_105_n278,
         DP_mult_105_n277, DP_mult_105_n276, DP_mult_105_n275,
         DP_mult_105_n274, DP_mult_105_n273, DP_mult_105_n272,
         DP_mult_105_n271, DP_mult_105_n270, DP_mult_105_n269,
         DP_mult_105_n268, DP_mult_105_n267, DP_mult_105_n266,
         DP_mult_105_n265, DP_mult_105_n264, DP_mult_105_n263,
         DP_mult_105_n259, DP_mult_105_n258, DP_mult_105_n257,
         DP_mult_105_n256, DP_mult_105_n255, DP_mult_105_n254,
         DP_mult_105_n253, DP_mult_105_n252, DP_mult_105_n251,
         DP_mult_105_n250, DP_mult_105_n249, DP_mult_105_n248,
         DP_mult_105_n247, DP_mult_105_n246, DP_mult_105_n245,
         DP_mult_105_n244, DP_mult_105_n243, DP_mult_105_n242,
         DP_mult_105_n241, DP_mult_105_n240, DP_mult_105_n239,
         DP_mult_105_n238, DP_mult_105_n237, DP_mult_105_n236,
         DP_mult_105_n235, DP_mult_105_n234, DP_mult_105_n233,
         DP_mult_105_n232, DP_mult_105_n231, DP_mult_105_n230,
         DP_mult_105_n229, DP_mult_105_n228, DP_mult_105_n227,
         DP_mult_105_n226, DP_mult_105_n225, DP_mult_105_n224,
         DP_mult_105_n223, DP_mult_105_n222, DP_mult_105_n221,
         DP_mult_105_n220, DP_mult_105_n219, DP_mult_105_n218,
         DP_mult_105_n217, DP_mult_105_n216, DP_mult_105_n215,
         DP_mult_105_n214, DP_mult_105_n213, DP_mult_105_n212,
         DP_mult_105_n211, DP_mult_105_n210, DP_mult_105_n209,
         DP_mult_105_n208, DP_mult_105_n207, DP_mult_105_n206,
         DP_mult_105_n205, DP_mult_105_n204, DP_mult_105_n203,
         DP_mult_105_n202, DP_mult_105_n201, DP_mult_105_n200,
         DP_mult_105_n199, DP_mult_105_n198, DP_mult_105_n197,
         DP_mult_105_n196, DP_mult_105_n195, DP_mult_105_n194,
         DP_mult_105_n193, DP_mult_105_n192, DP_mult_105_n191,
         DP_mult_105_n190, DP_mult_105_n189, DP_mult_105_n188,
         DP_mult_105_n187, DP_mult_105_n186, DP_mult_105_n185,
         DP_mult_105_n184, DP_mult_105_n183, DP_mult_105_n182,
         DP_mult_105_n181, DP_mult_105_n180, DP_mult_105_n179,
         DP_mult_105_n178, DP_mult_105_n177, DP_mult_105_n176,
         DP_mult_105_n175, DP_mult_105_n174, DP_mult_105_n173,
         DP_mult_105_n172, DP_mult_105_n171, DP_mult_105_n170,
         DP_mult_105_n169, DP_mult_105_n168, DP_mult_105_n167,
         DP_mult_105_n166, DP_mult_105_n165, DP_mult_105_n164,
         DP_mult_105_n163, DP_mult_105_n162, DP_mult_105_n161,
         DP_mult_105_n160, DP_mult_105_n159, DP_mult_105_n158,
         DP_mult_105_n157, DP_mult_105_n156, DP_mult_105_n155,
         DP_mult_105_n154, DP_mult_105_n153, DP_mult_105_n152,
         DP_mult_105_n151, DP_mult_105_n150, DP_mult_105_n149,
         DP_mult_105_n148, DP_mult_105_n147, DP_mult_105_n146,
         DP_mult_105_n145, DP_mult_105_n144, DP_mult_105_n143,
         DP_mult_105_n142, DP_mult_105_n141, DP_mult_105_n140,
         DP_mult_105_n139, DP_mult_105_n138, DP_mult_105_n126,
         DP_mult_105_n125, DP_mult_105_n124, DP_mult_105_n123,
         DP_mult_105_n122, DP_mult_105_n121, DP_mult_105_n120,
         DP_mult_105_n119, DP_mult_105_n118, DP_mult_105_n117,
         DP_mult_105_n116, DP_mult_105_n115,
         DP_sub_1_root_sub_0_root_sub_104_B_not_0_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_1_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_2_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_3_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_4_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_5_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_6_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_7_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_8_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_9_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_10_,
         DP_sub_1_root_sub_0_root_sub_104_B_not_12_,
         DP_sub_1_root_sub_0_root_sub_104_carry_1_,
         DP_sub_1_root_sub_0_root_sub_104_carry_2_,
         DP_sub_1_root_sub_0_root_sub_104_carry_3_,
         DP_sub_1_root_sub_0_root_sub_104_carry_4_,
         DP_sub_1_root_sub_0_root_sub_104_carry_5_,
         DP_sub_1_root_sub_0_root_sub_104_carry_6_,
         DP_sub_1_root_sub_0_root_sub_104_carry_7_,
         DP_sub_1_root_sub_0_root_sub_104_carry_8_,
         DP_sub_1_root_sub_0_root_sub_104_carry_9_,
         DP_sub_1_root_sub_0_root_sub_104_carry_10_,
         DP_sub_1_root_sub_0_root_sub_104_carry_11_,
         DP_sub_1_root_sub_0_root_sub_104_carry_12_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_0_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_1_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_2_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_3_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_4_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_5_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_6_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_7_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_8_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_9_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_10_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_12_,
         DP_sub_0_root_sub_0_root_sub_104_carry_1_,
         DP_sub_0_root_sub_0_root_sub_104_carry_2_,
         DP_sub_0_root_sub_0_root_sub_104_carry_3_,
         DP_sub_0_root_sub_0_root_sub_104_carry_4_,
         DP_sub_0_root_sub_0_root_sub_104_carry_5_,
         DP_sub_0_root_sub_0_root_sub_104_carry_6_,
         DP_sub_0_root_sub_0_root_sub_104_carry_7_,
         DP_sub_0_root_sub_0_root_sub_104_carry_8_,
         DP_sub_0_root_sub_0_root_sub_104_carry_9_,
         DP_sub_0_root_sub_0_root_sub_104_carry_10_,
         DP_sub_0_root_sub_0_root_sub_104_carry_11_,
         DP_sub_0_root_sub_0_root_sub_104_carry_12_, DP_mult_97_n660,
         DP_mult_97_n659, DP_mult_97_n658, DP_mult_97_n657, DP_mult_97_n656,
         DP_mult_97_n655, DP_mult_97_n654, DP_mult_97_n653, DP_mult_97_n652,
         DP_mult_97_n651, DP_mult_97_n650, DP_mult_97_n649, DP_mult_97_n648,
         DP_mult_97_n647, DP_mult_97_n646, DP_mult_97_n645, DP_mult_97_n644,
         DP_mult_97_n643, DP_mult_97_n642, DP_mult_97_n641, DP_mult_97_n640,
         DP_mult_97_n639, DP_mult_97_n638, DP_mult_97_n637, DP_mult_97_n636,
         DP_mult_97_n635, DP_mult_97_n634, DP_mult_97_n633, DP_mult_97_n632,
         DP_mult_97_n631, DP_mult_97_n630, DP_mult_97_n629, DP_mult_97_n628,
         DP_mult_97_n627, DP_mult_97_n626, DP_mult_97_n625, DP_mult_97_n624,
         DP_mult_97_n623, DP_mult_97_n622, DP_mult_97_n621, DP_mult_97_n620,
         DP_mult_97_n619, DP_mult_97_n618, DP_mult_97_n617, DP_mult_97_n616,
         DP_mult_97_n615, DP_mult_97_n614, DP_mult_97_n613, DP_mult_97_n612,
         DP_mult_97_n611, DP_mult_97_n610, DP_mult_97_n609, DP_mult_97_n608,
         DP_mult_97_n607, DP_mult_97_n606, DP_mult_97_n605, DP_mult_97_n604,
         DP_mult_97_n603, DP_mult_97_n602, DP_mult_97_n601, DP_mult_97_n600,
         DP_mult_97_n599, DP_mult_97_n598, DP_mult_97_n597, DP_mult_97_n596,
         DP_mult_97_n595, DP_mult_97_n594, DP_mult_97_n593, DP_mult_97_n592,
         DP_mult_97_n591, DP_mult_97_n590, DP_mult_97_n589, DP_mult_97_n588,
         DP_mult_97_n587, DP_mult_97_n586, DP_mult_97_n585, DP_mult_97_n584,
         DP_mult_97_n583, DP_mult_97_n582, DP_mult_97_n581, DP_mult_97_n580,
         DP_mult_97_n579, DP_mult_97_n578, DP_mult_97_n577, DP_mult_97_n576,
         DP_mult_97_n575, DP_mult_97_n574, DP_mult_97_n573, DP_mult_97_n572,
         DP_mult_97_n571, DP_mult_97_n570, DP_mult_97_n569, DP_mult_97_n568,
         DP_mult_97_n567, DP_mult_97_n566, DP_mult_97_n565, DP_mult_97_n564,
         DP_mult_97_n563, DP_mult_97_n562, DP_mult_97_n561, DP_mult_97_n560,
         DP_mult_97_n559, DP_mult_97_n558, DP_mult_97_n557, DP_mult_97_n556,
         DP_mult_97_n555, DP_mult_97_n554, DP_mult_97_n553, DP_mult_97_n552,
         DP_mult_97_n551, DP_mult_97_n550, DP_mult_97_n549, DP_mult_97_n548,
         DP_mult_97_n547, DP_mult_97_n546, DP_mult_97_n545, DP_mult_97_n544,
         DP_mult_97_n543, DP_mult_97_n542, DP_mult_97_n541, DP_mult_97_n540,
         DP_mult_97_n539, DP_mult_97_n538, DP_mult_97_n537, DP_mult_97_n536,
         DP_mult_97_n535, DP_mult_97_n534, DP_mult_97_n533, DP_mult_97_n532,
         DP_mult_97_n531, DP_mult_97_n530, DP_mult_97_n529, DP_mult_97_n528,
         DP_mult_97_n527, DP_mult_97_n526, DP_mult_97_n525, DP_mult_97_n524,
         DP_mult_97_n523, DP_mult_97_n522, DP_mult_97_n521, DP_mult_97_n520,
         DP_mult_97_n519, DP_mult_97_n337, DP_mult_97_n336, DP_mult_97_n335,
         DP_mult_97_n334, DP_mult_97_n333, DP_mult_97_n332, DP_mult_97_n331,
         DP_mult_97_n330, DP_mult_97_n329, DP_mult_97_n328, DP_mult_97_n327,
         DP_mult_97_n325, DP_mult_97_n324, DP_mult_97_n323, DP_mult_97_n322,
         DP_mult_97_n321, DP_mult_97_n320, DP_mult_97_n319, DP_mult_97_n318,
         DP_mult_97_n317, DP_mult_97_n316, DP_mult_97_n315, DP_mult_97_n314,
         DP_mult_97_n313, DP_mult_97_n312, DP_mult_97_n311, DP_mult_97_n310,
         DP_mult_97_n309, DP_mult_97_n308, DP_mult_97_n307, DP_mult_97_n306,
         DP_mult_97_n305, DP_mult_97_n303, DP_mult_97_n302, DP_mult_97_n301,
         DP_mult_97_n300, DP_mult_97_n299, DP_mult_97_n298, DP_mult_97_n297,
         DP_mult_97_n296, DP_mult_97_n295, DP_mult_97_n294, DP_mult_97_n293,
         DP_mult_97_n292, DP_mult_97_n291, DP_mult_97_n290, DP_mult_97_n289,
         DP_mult_97_n288, DP_mult_97_n287, DP_mult_97_n286, DP_mult_97_n285,
         DP_mult_97_n284, DP_mult_97_n283, DP_mult_97_n281, DP_mult_97_n280,
         DP_mult_97_n279, DP_mult_97_n278, DP_mult_97_n277, DP_mult_97_n276,
         DP_mult_97_n275, DP_mult_97_n274, DP_mult_97_n273, DP_mult_97_n272,
         DP_mult_97_n271, DP_mult_97_n270, DP_mult_97_n269, DP_mult_97_n268,
         DP_mult_97_n267, DP_mult_97_n266, DP_mult_97_n265, DP_mult_97_n264,
         DP_mult_97_n263, DP_mult_97_n259, DP_mult_97_n258, DP_mult_97_n257,
         DP_mult_97_n256, DP_mult_97_n255, DP_mult_97_n254, DP_mult_97_n253,
         DP_mult_97_n252, DP_mult_97_n251, DP_mult_97_n250, DP_mult_97_n249,
         DP_mult_97_n248, DP_mult_97_n247, DP_mult_97_n246, DP_mult_97_n245,
         DP_mult_97_n244, DP_mult_97_n243, DP_mult_97_n242, DP_mult_97_n241,
         DP_mult_97_n240, DP_mult_97_n239, DP_mult_97_n238, DP_mult_97_n237,
         DP_mult_97_n236, DP_mult_97_n235, DP_mult_97_n234, DP_mult_97_n233,
         DP_mult_97_n232, DP_mult_97_n231, DP_mult_97_n230, DP_mult_97_n229,
         DP_mult_97_n228, DP_mult_97_n227, DP_mult_97_n226, DP_mult_97_n225,
         DP_mult_97_n224, DP_mult_97_n223, DP_mult_97_n222, DP_mult_97_n221,
         DP_mult_97_n220, DP_mult_97_n219, DP_mult_97_n218, DP_mult_97_n217,
         DP_mult_97_n216, DP_mult_97_n215, DP_mult_97_n214, DP_mult_97_n213,
         DP_mult_97_n212, DP_mult_97_n211, DP_mult_97_n210, DP_mult_97_n209,
         DP_mult_97_n208, DP_mult_97_n207, DP_mult_97_n206, DP_mult_97_n205,
         DP_mult_97_n204, DP_mult_97_n203, DP_mult_97_n202, DP_mult_97_n201,
         DP_mult_97_n200, DP_mult_97_n199, DP_mult_97_n198, DP_mult_97_n197,
         DP_mult_97_n196, DP_mult_97_n195, DP_mult_97_n194, DP_mult_97_n193,
         DP_mult_97_n192, DP_mult_97_n191, DP_mult_97_n190, DP_mult_97_n189,
         DP_mult_97_n188, DP_mult_97_n187, DP_mult_97_n186, DP_mult_97_n185,
         DP_mult_97_n184, DP_mult_97_n183, DP_mult_97_n182, DP_mult_97_n181,
         DP_mult_97_n180, DP_mult_97_n179, DP_mult_97_n178, DP_mult_97_n177,
         DP_mult_97_n176, DP_mult_97_n175, DP_mult_97_n174, DP_mult_97_n173,
         DP_mult_97_n172, DP_mult_97_n171, DP_mult_97_n170, DP_mult_97_n169,
         DP_mult_97_n168, DP_mult_97_n167, DP_mult_97_n166, DP_mult_97_n165,
         DP_mult_97_n164, DP_mult_97_n163, DP_mult_97_n162, DP_mult_97_n161,
         DP_mult_97_n160, DP_mult_97_n159, DP_mult_97_n158, DP_mult_97_n157,
         DP_mult_97_n156, DP_mult_97_n155, DP_mult_97_n154, DP_mult_97_n153,
         DP_mult_97_n152, DP_mult_97_n151, DP_mult_97_n150, DP_mult_97_n149,
         DP_mult_97_n148, DP_mult_97_n147, DP_mult_97_n146, DP_mult_97_n145,
         DP_mult_97_n144, DP_mult_97_n143, DP_mult_97_n142, DP_mult_97_n141,
         DP_mult_97_n140, DP_mult_97_n139, DP_mult_97_n138, DP_mult_97_n126,
         DP_mult_97_n125, DP_mult_97_n124, DP_mult_97_n123, DP_mult_97_n122,
         DP_mult_97_n121, DP_mult_97_n120, DP_mult_97_n119, DP_mult_97_n118,
         DP_mult_97_n117, DP_mult_97_n116, DP_mult_97_n115, DP_mult_99_n660,
         DP_mult_99_n659, DP_mult_99_n658, DP_mult_99_n657, DP_mult_99_n656,
         DP_mult_99_n655, DP_mult_99_n654, DP_mult_99_n653, DP_mult_99_n652,
         DP_mult_99_n651, DP_mult_99_n650, DP_mult_99_n649, DP_mult_99_n648,
         DP_mult_99_n647, DP_mult_99_n646, DP_mult_99_n645, DP_mult_99_n644,
         DP_mult_99_n643, DP_mult_99_n642, DP_mult_99_n641, DP_mult_99_n640,
         DP_mult_99_n639, DP_mult_99_n638, DP_mult_99_n637, DP_mult_99_n636,
         DP_mult_99_n635, DP_mult_99_n634, DP_mult_99_n633, DP_mult_99_n632,
         DP_mult_99_n631, DP_mult_99_n630, DP_mult_99_n629, DP_mult_99_n628,
         DP_mult_99_n627, DP_mult_99_n626, DP_mult_99_n625, DP_mult_99_n624,
         DP_mult_99_n623, DP_mult_99_n622, DP_mult_99_n621, DP_mult_99_n620,
         DP_mult_99_n619, DP_mult_99_n618, DP_mult_99_n617, DP_mult_99_n616,
         DP_mult_99_n615, DP_mult_99_n614, DP_mult_99_n613, DP_mult_99_n612,
         DP_mult_99_n611, DP_mult_99_n610, DP_mult_99_n609, DP_mult_99_n608,
         DP_mult_99_n607, DP_mult_99_n606, DP_mult_99_n605, DP_mult_99_n604,
         DP_mult_99_n603, DP_mult_99_n602, DP_mult_99_n601, DP_mult_99_n600,
         DP_mult_99_n599, DP_mult_99_n598, DP_mult_99_n597, DP_mult_99_n596,
         DP_mult_99_n595, DP_mult_99_n594, DP_mult_99_n593, DP_mult_99_n592,
         DP_mult_99_n591, DP_mult_99_n590, DP_mult_99_n589, DP_mult_99_n588,
         DP_mult_99_n587, DP_mult_99_n586, DP_mult_99_n585, DP_mult_99_n584,
         DP_mult_99_n583, DP_mult_99_n582, DP_mult_99_n581, DP_mult_99_n580,
         DP_mult_99_n579, DP_mult_99_n578, DP_mult_99_n577, DP_mult_99_n576,
         DP_mult_99_n575, DP_mult_99_n574, DP_mult_99_n573, DP_mult_99_n572,
         DP_mult_99_n571, DP_mult_99_n570, DP_mult_99_n569, DP_mult_99_n568,
         DP_mult_99_n567, DP_mult_99_n566, DP_mult_99_n565, DP_mult_99_n564,
         DP_mult_99_n563, DP_mult_99_n562, DP_mult_99_n561, DP_mult_99_n560,
         DP_mult_99_n559, DP_mult_99_n558, DP_mult_99_n557, DP_mult_99_n556,
         DP_mult_99_n555, DP_mult_99_n554, DP_mult_99_n553, DP_mult_99_n552,
         DP_mult_99_n551, DP_mult_99_n550, DP_mult_99_n549, DP_mult_99_n548,
         DP_mult_99_n547, DP_mult_99_n546, DP_mult_99_n545, DP_mult_99_n544,
         DP_mult_99_n543, DP_mult_99_n542, DP_mult_99_n541, DP_mult_99_n540,
         DP_mult_99_n539, DP_mult_99_n538, DP_mult_99_n537, DP_mult_99_n536,
         DP_mult_99_n535, DP_mult_99_n534, DP_mult_99_n533, DP_mult_99_n532,
         DP_mult_99_n531, DP_mult_99_n530, DP_mult_99_n529, DP_mult_99_n528,
         DP_mult_99_n527, DP_mult_99_n526, DP_mult_99_n525, DP_mult_99_n524,
         DP_mult_99_n523, DP_mult_99_n522, DP_mult_99_n521, DP_mult_99_n520,
         DP_mult_99_n519, DP_mult_99_n337, DP_mult_99_n336, DP_mult_99_n335,
         DP_mult_99_n334, DP_mult_99_n333, DP_mult_99_n332, DP_mult_99_n331,
         DP_mult_99_n330, DP_mult_99_n329, DP_mult_99_n328, DP_mult_99_n327,
         DP_mult_99_n325, DP_mult_99_n324, DP_mult_99_n323, DP_mult_99_n322,
         DP_mult_99_n321, DP_mult_99_n320, DP_mult_99_n319, DP_mult_99_n318,
         DP_mult_99_n317, DP_mult_99_n316, DP_mult_99_n315, DP_mult_99_n314,
         DP_mult_99_n313, DP_mult_99_n312, DP_mult_99_n311, DP_mult_99_n310,
         DP_mult_99_n309, DP_mult_99_n308, DP_mult_99_n307, DP_mult_99_n306,
         DP_mult_99_n305, DP_mult_99_n303, DP_mult_99_n302, DP_mult_99_n301,
         DP_mult_99_n300, DP_mult_99_n299, DP_mult_99_n298, DP_mult_99_n297,
         DP_mult_99_n296, DP_mult_99_n295, DP_mult_99_n294, DP_mult_99_n293,
         DP_mult_99_n292, DP_mult_99_n291, DP_mult_99_n290, DP_mult_99_n289,
         DP_mult_99_n288, DP_mult_99_n287, DP_mult_99_n286, DP_mult_99_n285,
         DP_mult_99_n284, DP_mult_99_n283, DP_mult_99_n281, DP_mult_99_n280,
         DP_mult_99_n279, DP_mult_99_n278, DP_mult_99_n277, DP_mult_99_n276,
         DP_mult_99_n275, DP_mult_99_n274, DP_mult_99_n273, DP_mult_99_n272,
         DP_mult_99_n271, DP_mult_99_n270, DP_mult_99_n269, DP_mult_99_n268,
         DP_mult_99_n267, DP_mult_99_n266, DP_mult_99_n265, DP_mult_99_n264,
         DP_mult_99_n263, DP_mult_99_n259, DP_mult_99_n258, DP_mult_99_n257,
         DP_mult_99_n256, DP_mult_99_n255, DP_mult_99_n254, DP_mult_99_n253,
         DP_mult_99_n252, DP_mult_99_n251, DP_mult_99_n250, DP_mult_99_n249,
         DP_mult_99_n248, DP_mult_99_n247, DP_mult_99_n246, DP_mult_99_n245,
         DP_mult_99_n244, DP_mult_99_n243, DP_mult_99_n242, DP_mult_99_n241,
         DP_mult_99_n240, DP_mult_99_n239, DP_mult_99_n238, DP_mult_99_n237,
         DP_mult_99_n236, DP_mult_99_n235, DP_mult_99_n234, DP_mult_99_n233,
         DP_mult_99_n232, DP_mult_99_n231, DP_mult_99_n230, DP_mult_99_n229,
         DP_mult_99_n228, DP_mult_99_n227, DP_mult_99_n226, DP_mult_99_n225,
         DP_mult_99_n224, DP_mult_99_n223, DP_mult_99_n222, DP_mult_99_n221,
         DP_mult_99_n220, DP_mult_99_n219, DP_mult_99_n218, DP_mult_99_n217,
         DP_mult_99_n216, DP_mult_99_n215, DP_mult_99_n214, DP_mult_99_n213,
         DP_mult_99_n212, DP_mult_99_n211, DP_mult_99_n210, DP_mult_99_n209,
         DP_mult_99_n208, DP_mult_99_n207, DP_mult_99_n206, DP_mult_99_n205,
         DP_mult_99_n204, DP_mult_99_n203, DP_mult_99_n202, DP_mult_99_n201,
         DP_mult_99_n200, DP_mult_99_n199, DP_mult_99_n198, DP_mult_99_n197,
         DP_mult_99_n196, DP_mult_99_n195, DP_mult_99_n194, DP_mult_99_n193,
         DP_mult_99_n192, DP_mult_99_n191, DP_mult_99_n190, DP_mult_99_n189,
         DP_mult_99_n188, DP_mult_99_n187, DP_mult_99_n186, DP_mult_99_n185,
         DP_mult_99_n184, DP_mult_99_n183, DP_mult_99_n182, DP_mult_99_n181,
         DP_mult_99_n180, DP_mult_99_n179, DP_mult_99_n178, DP_mult_99_n177,
         DP_mult_99_n176, DP_mult_99_n175, DP_mult_99_n174, DP_mult_99_n173,
         DP_mult_99_n172, DP_mult_99_n171, DP_mult_99_n170, DP_mult_99_n169,
         DP_mult_99_n168, DP_mult_99_n167, DP_mult_99_n166, DP_mult_99_n165,
         DP_mult_99_n164, DP_mult_99_n163, DP_mult_99_n162, DP_mult_99_n161,
         DP_mult_99_n160, DP_mult_99_n159, DP_mult_99_n158, DP_mult_99_n157,
         DP_mult_99_n156, DP_mult_99_n155, DP_mult_99_n154, DP_mult_99_n153,
         DP_mult_99_n152, DP_mult_99_n151, DP_mult_99_n150, DP_mult_99_n149,
         DP_mult_99_n148, DP_mult_99_n147, DP_mult_99_n146, DP_mult_99_n145,
         DP_mult_99_n144, DP_mult_99_n143, DP_mult_99_n142, DP_mult_99_n141,
         DP_mult_99_n140, DP_mult_99_n139, DP_mult_99_n138, DP_mult_99_n126,
         DP_mult_99_n125, DP_mult_99_n124, DP_mult_99_n123, DP_mult_99_n122,
         DP_mult_99_n121, DP_mult_99_n120, DP_mult_99_n119, DP_mult_99_n118,
         DP_mult_99_n117, DP_mult_99_n116, DP_mult_99_n115, DP_mult_96_n660,
         DP_mult_96_n659, DP_mult_96_n658, DP_mult_96_n657, DP_mult_96_n656,
         DP_mult_96_n655, DP_mult_96_n654, DP_mult_96_n653, DP_mult_96_n652,
         DP_mult_96_n651, DP_mult_96_n650, DP_mult_96_n649, DP_mult_96_n648,
         DP_mult_96_n647, DP_mult_96_n646, DP_mult_96_n645, DP_mult_96_n644,
         DP_mult_96_n643, DP_mult_96_n642, DP_mult_96_n641, DP_mult_96_n640,
         DP_mult_96_n639, DP_mult_96_n638, DP_mult_96_n637, DP_mult_96_n636,
         DP_mult_96_n635, DP_mult_96_n634, DP_mult_96_n633, DP_mult_96_n632,
         DP_mult_96_n631, DP_mult_96_n630, DP_mult_96_n629, DP_mult_96_n628,
         DP_mult_96_n627, DP_mult_96_n626, DP_mult_96_n625, DP_mult_96_n624,
         DP_mult_96_n623, DP_mult_96_n622, DP_mult_96_n621, DP_mult_96_n620,
         DP_mult_96_n619, DP_mult_96_n618, DP_mult_96_n617, DP_mult_96_n616,
         DP_mult_96_n615, DP_mult_96_n614, DP_mult_96_n613, DP_mult_96_n612,
         DP_mult_96_n611, DP_mult_96_n610, DP_mult_96_n609, DP_mult_96_n608,
         DP_mult_96_n607, DP_mult_96_n606, DP_mult_96_n605, DP_mult_96_n604,
         DP_mult_96_n603, DP_mult_96_n602, DP_mult_96_n601, DP_mult_96_n600,
         DP_mult_96_n599, DP_mult_96_n598, DP_mult_96_n597, DP_mult_96_n596,
         DP_mult_96_n595, DP_mult_96_n594, DP_mult_96_n593, DP_mult_96_n592,
         DP_mult_96_n591, DP_mult_96_n590, DP_mult_96_n589, DP_mult_96_n588,
         DP_mult_96_n587, DP_mult_96_n586, DP_mult_96_n585, DP_mult_96_n584,
         DP_mult_96_n583, DP_mult_96_n582, DP_mult_96_n581, DP_mult_96_n580,
         DP_mult_96_n579, DP_mult_96_n578, DP_mult_96_n577, DP_mult_96_n576,
         DP_mult_96_n575, DP_mult_96_n574, DP_mult_96_n573, DP_mult_96_n572,
         DP_mult_96_n571, DP_mult_96_n570, DP_mult_96_n569, DP_mult_96_n568,
         DP_mult_96_n567, DP_mult_96_n566, DP_mult_96_n565, DP_mult_96_n564,
         DP_mult_96_n563, DP_mult_96_n562, DP_mult_96_n561, DP_mult_96_n560,
         DP_mult_96_n559, DP_mult_96_n558, DP_mult_96_n557, DP_mult_96_n556,
         DP_mult_96_n555, DP_mult_96_n554, DP_mult_96_n553, DP_mult_96_n552,
         DP_mult_96_n551, DP_mult_96_n550, DP_mult_96_n549, DP_mult_96_n548,
         DP_mult_96_n547, DP_mult_96_n546, DP_mult_96_n545, DP_mult_96_n544,
         DP_mult_96_n543, DP_mult_96_n542, DP_mult_96_n541, DP_mult_96_n540,
         DP_mult_96_n539, DP_mult_96_n538, DP_mult_96_n537, DP_mult_96_n536,
         DP_mult_96_n535, DP_mult_96_n534, DP_mult_96_n533, DP_mult_96_n532,
         DP_mult_96_n531, DP_mult_96_n530, DP_mult_96_n529, DP_mult_96_n528,
         DP_mult_96_n527, DP_mult_96_n526, DP_mult_96_n525, DP_mult_96_n524,
         DP_mult_96_n523, DP_mult_96_n522, DP_mult_96_n521, DP_mult_96_n520,
         DP_mult_96_n519, DP_mult_96_n337, DP_mult_96_n336, DP_mult_96_n335,
         DP_mult_96_n334, DP_mult_96_n333, DP_mult_96_n332, DP_mult_96_n331,
         DP_mult_96_n330, DP_mult_96_n329, DP_mult_96_n328, DP_mult_96_n327,
         DP_mult_96_n325, DP_mult_96_n324, DP_mult_96_n323, DP_mult_96_n322,
         DP_mult_96_n321, DP_mult_96_n320, DP_mult_96_n319, DP_mult_96_n318,
         DP_mult_96_n317, DP_mult_96_n316, DP_mult_96_n315, DP_mult_96_n314,
         DP_mult_96_n313, DP_mult_96_n312, DP_mult_96_n311, DP_mult_96_n310,
         DP_mult_96_n309, DP_mult_96_n308, DP_mult_96_n307, DP_mult_96_n306,
         DP_mult_96_n305, DP_mult_96_n303, DP_mult_96_n302, DP_mult_96_n301,
         DP_mult_96_n300, DP_mult_96_n299, DP_mult_96_n298, DP_mult_96_n297,
         DP_mult_96_n296, DP_mult_96_n295, DP_mult_96_n294, DP_mult_96_n293,
         DP_mult_96_n292, DP_mult_96_n291, DP_mult_96_n290, DP_mult_96_n289,
         DP_mult_96_n288, DP_mult_96_n287, DP_mult_96_n286, DP_mult_96_n285,
         DP_mult_96_n284, DP_mult_96_n283, DP_mult_96_n281, DP_mult_96_n280,
         DP_mult_96_n279, DP_mult_96_n278, DP_mult_96_n277, DP_mult_96_n276,
         DP_mult_96_n275, DP_mult_96_n274, DP_mult_96_n273, DP_mult_96_n272,
         DP_mult_96_n271, DP_mult_96_n270, DP_mult_96_n269, DP_mult_96_n268,
         DP_mult_96_n267, DP_mult_96_n266, DP_mult_96_n265, DP_mult_96_n264,
         DP_mult_96_n263, DP_mult_96_n259, DP_mult_96_n258, DP_mult_96_n257,
         DP_mult_96_n256, DP_mult_96_n255, DP_mult_96_n254, DP_mult_96_n253,
         DP_mult_96_n252, DP_mult_96_n251, DP_mult_96_n250, DP_mult_96_n249,
         DP_mult_96_n248, DP_mult_96_n247, DP_mult_96_n246, DP_mult_96_n245,
         DP_mult_96_n244, DP_mult_96_n243, DP_mult_96_n242, DP_mult_96_n241,
         DP_mult_96_n240, DP_mult_96_n239, DP_mult_96_n238, DP_mult_96_n237,
         DP_mult_96_n236, DP_mult_96_n235, DP_mult_96_n234, DP_mult_96_n233,
         DP_mult_96_n232, DP_mult_96_n231, DP_mult_96_n230, DP_mult_96_n229,
         DP_mult_96_n228, DP_mult_96_n227, DP_mult_96_n226, DP_mult_96_n225,
         DP_mult_96_n224, DP_mult_96_n223, DP_mult_96_n222, DP_mult_96_n221,
         DP_mult_96_n220, DP_mult_96_n219, DP_mult_96_n218, DP_mult_96_n217,
         DP_mult_96_n216, DP_mult_96_n215, DP_mult_96_n214, DP_mult_96_n213,
         DP_mult_96_n212, DP_mult_96_n211, DP_mult_96_n210, DP_mult_96_n209,
         DP_mult_96_n208, DP_mult_96_n207, DP_mult_96_n206, DP_mult_96_n205,
         DP_mult_96_n204, DP_mult_96_n203, DP_mult_96_n202, DP_mult_96_n201,
         DP_mult_96_n200, DP_mult_96_n199, DP_mult_96_n198, DP_mult_96_n197,
         DP_mult_96_n196, DP_mult_96_n195, DP_mult_96_n194, DP_mult_96_n193,
         DP_mult_96_n192, DP_mult_96_n191, DP_mult_96_n190, DP_mult_96_n189,
         DP_mult_96_n188, DP_mult_96_n187, DP_mult_96_n186, DP_mult_96_n185,
         DP_mult_96_n184, DP_mult_96_n183, DP_mult_96_n182, DP_mult_96_n181,
         DP_mult_96_n180, DP_mult_96_n179, DP_mult_96_n178, DP_mult_96_n177,
         DP_mult_96_n176, DP_mult_96_n175, DP_mult_96_n174, DP_mult_96_n173,
         DP_mult_96_n172, DP_mult_96_n171, DP_mult_96_n170, DP_mult_96_n169,
         DP_mult_96_n168, DP_mult_96_n167, DP_mult_96_n166, DP_mult_96_n165,
         DP_mult_96_n164, DP_mult_96_n163, DP_mult_96_n162, DP_mult_96_n161,
         DP_mult_96_n160, DP_mult_96_n159, DP_mult_96_n158, DP_mult_96_n157,
         DP_mult_96_n156, DP_mult_96_n155, DP_mult_96_n154, DP_mult_96_n153,
         DP_mult_96_n152, DP_mult_96_n151, DP_mult_96_n150, DP_mult_96_n149,
         DP_mult_96_n148, DP_mult_96_n147, DP_mult_96_n146, DP_mult_96_n145,
         DP_mult_96_n144, DP_mult_96_n143, DP_mult_96_n142, DP_mult_96_n141,
         DP_mult_96_n140, DP_mult_96_n139, DP_mult_96_n138, DP_mult_96_n126,
         DP_mult_96_n125, DP_mult_96_n124, DP_mult_96_n123, DP_mult_96_n122,
         DP_mult_96_n121, DP_mult_96_n120, DP_mult_96_n119, DP_mult_96_n118,
         DP_mult_96_n117, DP_mult_96_n116, DP_mult_96_n115, DP_mult_98_n660,
         DP_mult_98_n659, DP_mult_98_n658, DP_mult_98_n657, DP_mult_98_n656,
         DP_mult_98_n655, DP_mult_98_n654, DP_mult_98_n653, DP_mult_98_n652,
         DP_mult_98_n651, DP_mult_98_n650, DP_mult_98_n649, DP_mult_98_n648,
         DP_mult_98_n647, DP_mult_98_n646, DP_mult_98_n645, DP_mult_98_n644,
         DP_mult_98_n643, DP_mult_98_n642, DP_mult_98_n641, DP_mult_98_n640,
         DP_mult_98_n639, DP_mult_98_n638, DP_mult_98_n637, DP_mult_98_n636,
         DP_mult_98_n635, DP_mult_98_n634, DP_mult_98_n633, DP_mult_98_n632,
         DP_mult_98_n631, DP_mult_98_n630, DP_mult_98_n629, DP_mult_98_n628,
         DP_mult_98_n627, DP_mult_98_n626, DP_mult_98_n625, DP_mult_98_n624,
         DP_mult_98_n623, DP_mult_98_n622, DP_mult_98_n621, DP_mult_98_n620,
         DP_mult_98_n619, DP_mult_98_n618, DP_mult_98_n617, DP_mult_98_n616,
         DP_mult_98_n615, DP_mult_98_n614, DP_mult_98_n613, DP_mult_98_n612,
         DP_mult_98_n611, DP_mult_98_n610, DP_mult_98_n609, DP_mult_98_n608,
         DP_mult_98_n607, DP_mult_98_n606, DP_mult_98_n605, DP_mult_98_n604,
         DP_mult_98_n603, DP_mult_98_n602, DP_mult_98_n601, DP_mult_98_n600,
         DP_mult_98_n599, DP_mult_98_n598, DP_mult_98_n597, DP_mult_98_n596,
         DP_mult_98_n595, DP_mult_98_n594, DP_mult_98_n593, DP_mult_98_n592,
         DP_mult_98_n591, DP_mult_98_n590, DP_mult_98_n589, DP_mult_98_n588,
         DP_mult_98_n587, DP_mult_98_n586, DP_mult_98_n585, DP_mult_98_n584,
         DP_mult_98_n583, DP_mult_98_n582, DP_mult_98_n581, DP_mult_98_n580,
         DP_mult_98_n579, DP_mult_98_n578, DP_mult_98_n577, DP_mult_98_n576,
         DP_mult_98_n575, DP_mult_98_n574, DP_mult_98_n573, DP_mult_98_n572,
         DP_mult_98_n571, DP_mult_98_n570, DP_mult_98_n569, DP_mult_98_n568,
         DP_mult_98_n567, DP_mult_98_n566, DP_mult_98_n565, DP_mult_98_n564,
         DP_mult_98_n563, DP_mult_98_n562, DP_mult_98_n561, DP_mult_98_n560,
         DP_mult_98_n559, DP_mult_98_n558, DP_mult_98_n557, DP_mult_98_n556,
         DP_mult_98_n555, DP_mult_98_n554, DP_mult_98_n553, DP_mult_98_n552,
         DP_mult_98_n551, DP_mult_98_n550, DP_mult_98_n549, DP_mult_98_n548,
         DP_mult_98_n547, DP_mult_98_n546, DP_mult_98_n545, DP_mult_98_n544,
         DP_mult_98_n543, DP_mult_98_n542, DP_mult_98_n541, DP_mult_98_n540,
         DP_mult_98_n539, DP_mult_98_n538, DP_mult_98_n537, DP_mult_98_n536,
         DP_mult_98_n535, DP_mult_98_n534, DP_mult_98_n533, DP_mult_98_n532,
         DP_mult_98_n531, DP_mult_98_n530, DP_mult_98_n529, DP_mult_98_n528,
         DP_mult_98_n527, DP_mult_98_n526, DP_mult_98_n525, DP_mult_98_n524,
         DP_mult_98_n523, DP_mult_98_n522, DP_mult_98_n521, DP_mult_98_n520,
         DP_mult_98_n519, DP_mult_98_n337, DP_mult_98_n336, DP_mult_98_n335,
         DP_mult_98_n334, DP_mult_98_n333, DP_mult_98_n332, DP_mult_98_n331,
         DP_mult_98_n330, DP_mult_98_n329, DP_mult_98_n328, DP_mult_98_n327,
         DP_mult_98_n325, DP_mult_98_n324, DP_mult_98_n323, DP_mult_98_n322,
         DP_mult_98_n321, DP_mult_98_n320, DP_mult_98_n319, DP_mult_98_n318,
         DP_mult_98_n317, DP_mult_98_n316, DP_mult_98_n315, DP_mult_98_n314,
         DP_mult_98_n313, DP_mult_98_n312, DP_mult_98_n311, DP_mult_98_n310,
         DP_mult_98_n309, DP_mult_98_n308, DP_mult_98_n307, DP_mult_98_n306,
         DP_mult_98_n305, DP_mult_98_n303, DP_mult_98_n302, DP_mult_98_n301,
         DP_mult_98_n300, DP_mult_98_n299, DP_mult_98_n298, DP_mult_98_n297,
         DP_mult_98_n296, DP_mult_98_n295, DP_mult_98_n294, DP_mult_98_n293,
         DP_mult_98_n292, DP_mult_98_n291, DP_mult_98_n290, DP_mult_98_n289,
         DP_mult_98_n288, DP_mult_98_n287, DP_mult_98_n286, DP_mult_98_n285,
         DP_mult_98_n284, DP_mult_98_n283, DP_mult_98_n281, DP_mult_98_n280,
         DP_mult_98_n279, DP_mult_98_n278, DP_mult_98_n277, DP_mult_98_n276,
         DP_mult_98_n275, DP_mult_98_n274, DP_mult_98_n273, DP_mult_98_n272,
         DP_mult_98_n271, DP_mult_98_n270, DP_mult_98_n269, DP_mult_98_n268,
         DP_mult_98_n267, DP_mult_98_n266, DP_mult_98_n265, DP_mult_98_n264,
         DP_mult_98_n263, DP_mult_98_n259, DP_mult_98_n258, DP_mult_98_n257,
         DP_mult_98_n256, DP_mult_98_n255, DP_mult_98_n254, DP_mult_98_n253,
         DP_mult_98_n252, DP_mult_98_n251, DP_mult_98_n250, DP_mult_98_n249,
         DP_mult_98_n248, DP_mult_98_n247, DP_mult_98_n246, DP_mult_98_n245,
         DP_mult_98_n244, DP_mult_98_n243, DP_mult_98_n242, DP_mult_98_n241,
         DP_mult_98_n240, DP_mult_98_n239, DP_mult_98_n238, DP_mult_98_n237,
         DP_mult_98_n236, DP_mult_98_n235, DP_mult_98_n234, DP_mult_98_n233,
         DP_mult_98_n232, DP_mult_98_n231, DP_mult_98_n230, DP_mult_98_n229,
         DP_mult_98_n228, DP_mult_98_n227, DP_mult_98_n226, DP_mult_98_n225,
         DP_mult_98_n224, DP_mult_98_n223, DP_mult_98_n222, DP_mult_98_n221,
         DP_mult_98_n220, DP_mult_98_n219, DP_mult_98_n218, DP_mult_98_n217,
         DP_mult_98_n216, DP_mult_98_n215, DP_mult_98_n214, DP_mult_98_n213,
         DP_mult_98_n212, DP_mult_98_n211, DP_mult_98_n210, DP_mult_98_n209,
         DP_mult_98_n208, DP_mult_98_n207, DP_mult_98_n206, DP_mult_98_n205,
         DP_mult_98_n204, DP_mult_98_n203, DP_mult_98_n202, DP_mult_98_n201,
         DP_mult_98_n200, DP_mult_98_n199, DP_mult_98_n198, DP_mult_98_n197,
         DP_mult_98_n196, DP_mult_98_n195, DP_mult_98_n194, DP_mult_98_n193,
         DP_mult_98_n192, DP_mult_98_n191, DP_mult_98_n190, DP_mult_98_n189,
         DP_mult_98_n188, DP_mult_98_n187, DP_mult_98_n186, DP_mult_98_n185,
         DP_mult_98_n184, DP_mult_98_n183, DP_mult_98_n182, DP_mult_98_n181,
         DP_mult_98_n180, DP_mult_98_n179, DP_mult_98_n178, DP_mult_98_n177,
         DP_mult_98_n176, DP_mult_98_n175, DP_mult_98_n174, DP_mult_98_n173,
         DP_mult_98_n172, DP_mult_98_n171, DP_mult_98_n170, DP_mult_98_n169,
         DP_mult_98_n168, DP_mult_98_n167, DP_mult_98_n166, DP_mult_98_n165,
         DP_mult_98_n164, DP_mult_98_n163, DP_mult_98_n162, DP_mult_98_n161,
         DP_mult_98_n160, DP_mult_98_n159, DP_mult_98_n158, DP_mult_98_n157,
         DP_mult_98_n156, DP_mult_98_n155, DP_mult_98_n154, DP_mult_98_n153,
         DP_mult_98_n152, DP_mult_98_n151, DP_mult_98_n150, DP_mult_98_n149,
         DP_mult_98_n148, DP_mult_98_n147, DP_mult_98_n146, DP_mult_98_n145,
         DP_mult_98_n144, DP_mult_98_n143, DP_mult_98_n142, DP_mult_98_n141,
         DP_mult_98_n140, DP_mult_98_n139, DP_mult_98_n138, DP_mult_98_n126,
         DP_mult_98_n125, DP_mult_98_n124, DP_mult_98_n123, DP_mult_98_n122,
         DP_mult_98_n121, DP_mult_98_n120, DP_mult_98_n119, DP_mult_98_n118,
         DP_mult_98_n117, DP_mult_98_n116, DP_mult_98_n115, CU_nextState_0_,
         CU_presentState_0_;
  wire   [0:11] DP_y;
  wire   [35:0] DP_b_int;
  wire   [23:0] DP_a_int;

  INV_X1 DP_U30 ( .A(DP_y[11]), .ZN(DP_n17) );
  NAND2_X1 DP_U29 ( .A1(DP_y[0]), .A2(DP_n6), .ZN(DP_n16) );
  NAND2_X1 DP_U28 ( .A1(DP_n4), .A2(DP_n16), .ZN(DP_y_out_0_) );
  NAND2_X1 DP_U27 ( .A1(DP_y[10]), .A2(DP_n6), .ZN(DP_n15) );
  NAND2_X1 DP_U26 ( .A1(DP_n4), .A2(DP_n15), .ZN(DP_y_out_10_) );
  NAND2_X1 DP_U25 ( .A1(DP_y[1]), .A2(DP_n6), .ZN(DP_n14) );
  NAND2_X1 DP_U24 ( .A1(DP_n4), .A2(DP_n14), .ZN(DP_y_out_1_) );
  NAND2_X1 DP_U23 ( .A1(DP_y[2]), .A2(DP_n6), .ZN(DP_n13) );
  NAND2_X1 DP_U22 ( .A1(DP_n4), .A2(DP_n13), .ZN(DP_y_out_2_) );
  NAND2_X1 DP_U21 ( .A1(DP_y[3]), .A2(DP_n6), .ZN(DP_n12) );
  NAND2_X1 DP_U20 ( .A1(DP_n4), .A2(DP_n12), .ZN(DP_y_out_3_) );
  NAND2_X1 DP_U19 ( .A1(DP_y[4]), .A2(DP_n6), .ZN(DP_n11) );
  NAND2_X1 DP_U18 ( .A1(DP_n4), .A2(DP_n11), .ZN(DP_y_out_4_) );
  NAND2_X1 DP_U17 ( .A1(DP_y[5]), .A2(DP_n6), .ZN(DP_n10) );
  NAND2_X1 DP_U16 ( .A1(DP_n4), .A2(DP_n10), .ZN(DP_y_out_5_) );
  NAND2_X1 DP_U15 ( .A1(DP_y[6]), .A2(DP_n6), .ZN(DP_n9) );
  NAND2_X1 DP_U14 ( .A1(DP_n4), .A2(DP_n9), .ZN(DP_y_out_6_) );
  NAND2_X1 DP_U13 ( .A1(DP_y[7]), .A2(DP_n6), .ZN(DP_n8) );
  NAND2_X1 DP_U12 ( .A1(DP_n4), .A2(DP_n8), .ZN(DP_y_out_7_) );
  NAND2_X1 DP_U11 ( .A1(DP_y[8]), .A2(DP_n6), .ZN(DP_n7) );
  NAND2_X1 DP_U10 ( .A1(DP_n4), .A2(DP_n7), .ZN(DP_y_out_8_) );
  NAND2_X1 DP_U9 ( .A1(DP_y[9]), .A2(DP_n6), .ZN(DP_n5) );
  NAND2_X1 DP_U8 ( .A1(DP_n4), .A2(DP_n5), .ZN(DP_y_out_9_) );
  OR2_X1 DP_U7 ( .A1(DP_n17), .A2(DP_y_out_11_), .ZN(DP_n4) );
  NAND2_X1 DP_U6 ( .A1(DP_y_out_11_), .A2(DP_n17), .ZN(DP_n6) );
  CLKBUF_X2 DP_U5 ( .A(rst_n), .Z(DP_n3) );
  CLKBUF_X2 DP_U4 ( .A(rst_n), .Z(DP_n1) );
  CLKBUF_X2 DP_U3 ( .A(rst_n), .Z(DP_n2) );
  NAND2_X1 DP_reg_in_U28 ( .A1(dIn[11]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n12) );
  OAI21_X1 DP_reg_in_U27 ( .B1(DP_reg_in_n37), .B2(DP_reg_in_n24), .A(
        DP_reg_in_n12), .ZN(DP_reg_in_n36) );
  NAND2_X1 DP_reg_in_U26 ( .A1(dIn[10]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n11) );
  OAI21_X1 DP_reg_in_U25 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n23), .A(
        DP_reg_in_n11), .ZN(DP_reg_in_n35) );
  NAND2_X1 DP_reg_in_U24 ( .A1(dIn[9]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n10)
         );
  OAI21_X1 DP_reg_in_U23 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n22), .A(
        DP_reg_in_n10), .ZN(DP_reg_in_n34) );
  NAND2_X1 DP_reg_in_U22 ( .A1(dIn[8]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n9)
         );
  OAI21_X1 DP_reg_in_U21 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n21), .A(
        DP_reg_in_n9), .ZN(DP_reg_in_n33) );
  NAND2_X1 DP_reg_in_U20 ( .A1(dIn[7]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n8)
         );
  OAI21_X1 DP_reg_in_U19 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n20), .A(
        DP_reg_in_n8), .ZN(DP_reg_in_n32) );
  NAND2_X1 DP_reg_in_U18 ( .A1(dIn[6]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n7)
         );
  OAI21_X1 DP_reg_in_U17 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n19), .A(
        DP_reg_in_n7), .ZN(DP_reg_in_n31) );
  NAND2_X1 DP_reg_in_U16 ( .A1(dIn[5]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n6)
         );
  OAI21_X1 DP_reg_in_U15 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n18), .A(
        DP_reg_in_n6), .ZN(DP_reg_in_n30) );
  NAND2_X1 DP_reg_in_U14 ( .A1(dIn[4]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n5)
         );
  OAI21_X1 DP_reg_in_U13 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n17), .A(
        DP_reg_in_n5), .ZN(DP_reg_in_n29) );
  NAND2_X1 DP_reg_in_U12 ( .A1(dIn[3]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n4)
         );
  OAI21_X1 DP_reg_in_U11 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n16), .A(
        DP_reg_in_n4), .ZN(DP_reg_in_n28) );
  NAND2_X1 DP_reg_in_U10 ( .A1(dIn[2]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n3)
         );
  OAI21_X1 DP_reg_in_U9 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n15), .A(
        DP_reg_in_n3), .ZN(DP_reg_in_n27) );
  NAND2_X1 DP_reg_in_U8 ( .A1(dIn[1]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n2)
         );
  OAI21_X1 DP_reg_in_U7 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n14), .A(
        DP_reg_in_n2), .ZN(DP_reg_in_n26) );
  NAND2_X1 DP_reg_in_U6 ( .A1(DP_reg_in_n38), .A2(dIn[0]), .ZN(DP_reg_in_n1)
         );
  OAI21_X1 DP_reg_in_U5 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n13), .A(
        DP_reg_in_n1), .ZN(DP_reg_in_n25) );
  BUF_X1 DP_reg_in_U4 ( .A(vIn), .Z(DP_reg_in_n38) );
  BUF_X1 DP_reg_in_U3 ( .A(vIn), .Z(DP_reg_in_n37) );
  BUF_X1 DP_reg_in_U2 ( .A(DP_n2), .Z(DP_reg_in_n39) );
  DFFR_X1 DP_reg_in_Q_reg_0_ ( .D(DP_reg_in_n25), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_0_), .QN(DP_reg_in_n13) );
  DFFR_X1 DP_reg_in_Q_reg_1_ ( .D(DP_reg_in_n26), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_1_), .QN(DP_reg_in_n14) );
  DFFR_X1 DP_reg_in_Q_reg_2_ ( .D(DP_reg_in_n27), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_2_), .QN(DP_reg_in_n15) );
  DFFR_X1 DP_reg_in_Q_reg_3_ ( .D(DP_reg_in_n28), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_3_), .QN(DP_reg_in_n16) );
  DFFR_X1 DP_reg_in_Q_reg_4_ ( .D(DP_reg_in_n29), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_4_), .QN(DP_reg_in_n17) );
  DFFR_X1 DP_reg_in_Q_reg_5_ ( .D(DP_reg_in_n30), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_5_), .QN(DP_reg_in_n18) );
  DFFR_X1 DP_reg_in_Q_reg_6_ ( .D(DP_reg_in_n31), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_6_), .QN(DP_reg_in_n19) );
  DFFR_X1 DP_reg_in_Q_reg_7_ ( .D(DP_reg_in_n32), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_7_), .QN(DP_reg_in_n20) );
  DFFR_X1 DP_reg_in_Q_reg_8_ ( .D(DP_reg_in_n33), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_8_), .QN(DP_reg_in_n21) );
  DFFR_X1 DP_reg_in_Q_reg_9_ ( .D(DP_reg_in_n34), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_9_), .QN(DP_reg_in_n22) );
  DFFR_X1 DP_reg_in_Q_reg_10_ ( .D(DP_reg_in_n35), .CK(clk), .RN(DP_reg_in_n39), .Q(DP_x_10_), .QN(DP_reg_in_n23) );
  DFFR_X1 DP_reg_in_Q_reg_11_ ( .D(DP_reg_in_n36), .CK(clk), .RN(DP_reg_in_n39), .Q(DP_x_11_), .QN(DP_reg_in_n24) );
  NAND2_X1 DP_reg_a_i_1_U27 ( .A1(a[23]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n63) );
  OAI21_X1 DP_reg_a_i_1_U26 ( .B1(DP_reg_a_i_1_n37), .B2(DP_reg_a_i_1_n51), 
        .A(DP_reg_a_i_1_n63), .ZN(DP_reg_a_i_1_n39) );
  NAND2_X1 DP_reg_a_i_1_U25 ( .A1(a[22]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n64) );
  OAI21_X1 DP_reg_a_i_1_U24 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n52), 
        .A(DP_reg_a_i_1_n64), .ZN(DP_reg_a_i_1_n40) );
  NAND2_X1 DP_reg_a_i_1_U23 ( .A1(a[21]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n65) );
  OAI21_X1 DP_reg_a_i_1_U22 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n53), 
        .A(DP_reg_a_i_1_n65), .ZN(DP_reg_a_i_1_n41) );
  NAND2_X1 DP_reg_a_i_1_U21 ( .A1(a[20]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n66) );
  OAI21_X1 DP_reg_a_i_1_U20 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n54), 
        .A(DP_reg_a_i_1_n66), .ZN(DP_reg_a_i_1_n42) );
  NAND2_X1 DP_reg_a_i_1_U19 ( .A1(a[19]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n67) );
  OAI21_X1 DP_reg_a_i_1_U18 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n55), 
        .A(DP_reg_a_i_1_n67), .ZN(DP_reg_a_i_1_n43) );
  NAND2_X1 DP_reg_a_i_1_U17 ( .A1(a[18]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n68) );
  OAI21_X1 DP_reg_a_i_1_U16 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n56), 
        .A(DP_reg_a_i_1_n68), .ZN(DP_reg_a_i_1_n44) );
  NAND2_X1 DP_reg_a_i_1_U15 ( .A1(a[17]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n69) );
  OAI21_X1 DP_reg_a_i_1_U14 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n57), 
        .A(DP_reg_a_i_1_n69), .ZN(DP_reg_a_i_1_n45) );
  NAND2_X1 DP_reg_a_i_1_U13 ( .A1(a[16]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n70) );
  OAI21_X1 DP_reg_a_i_1_U12 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n58), 
        .A(DP_reg_a_i_1_n70), .ZN(DP_reg_a_i_1_n46) );
  NAND2_X1 DP_reg_a_i_1_U11 ( .A1(a[15]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n71) );
  OAI21_X1 DP_reg_a_i_1_U10 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n59), 
        .A(DP_reg_a_i_1_n71), .ZN(DP_reg_a_i_1_n47) );
  NAND2_X1 DP_reg_a_i_1_U9 ( .A1(a[14]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n72) );
  OAI21_X1 DP_reg_a_i_1_U8 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n60), .A(
        DP_reg_a_i_1_n72), .ZN(DP_reg_a_i_1_n48) );
  NAND2_X1 DP_reg_a_i_1_U7 ( .A1(a[13]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n73) );
  OAI21_X1 DP_reg_a_i_1_U6 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n61), .A(
        DP_reg_a_i_1_n73), .ZN(DP_reg_a_i_1_n49) );
  NAND2_X1 DP_reg_a_i_1_U5 ( .A1(DP_reg_a_i_1_n38), .A2(a[12]), .ZN(
        DP_reg_a_i_1_n74) );
  OAI21_X1 DP_reg_a_i_1_U4 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n62), .A(
        DP_reg_a_i_1_n74), .ZN(DP_reg_a_i_1_n50) );
  BUF_X1 DP_reg_a_i_1_U3 ( .A(vIn), .Z(DP_reg_a_i_1_n38) );
  BUF_X1 DP_reg_a_i_1_U2 ( .A(vIn), .Z(DP_reg_a_i_1_n37) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_0_ ( .D(DP_reg_a_i_1_n50), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[11]), .QN(DP_reg_a_i_1_n62) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_11_ ( .D(DP_reg_a_i_1_n39), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[0]), .QN(DP_reg_a_i_1_n51) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_1_ ( .D(DP_reg_a_i_1_n49), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[10]), .QN(DP_reg_a_i_1_n61) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_2_ ( .D(DP_reg_a_i_1_n48), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[9]), .QN(DP_reg_a_i_1_n60) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_3_ ( .D(DP_reg_a_i_1_n47), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[8]), .QN(DP_reg_a_i_1_n59) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_4_ ( .D(DP_reg_a_i_1_n46), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[7]), .QN(DP_reg_a_i_1_n58) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_5_ ( .D(DP_reg_a_i_1_n45), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[6]), .QN(DP_reg_a_i_1_n57) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_6_ ( .D(DP_reg_a_i_1_n44), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[5]), .QN(DP_reg_a_i_1_n56) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_7_ ( .D(DP_reg_a_i_1_n43), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[4]), .QN(DP_reg_a_i_1_n55) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_8_ ( .D(DP_reg_a_i_1_n42), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[3]), .QN(DP_reg_a_i_1_n54) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_9_ ( .D(DP_reg_a_i_1_n41), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[2]), .QN(DP_reg_a_i_1_n53) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_10_ ( .D(DP_reg_a_i_1_n40), .CK(clk), .RN(DP_n1), 
        .Q(DP_a_int[1]), .QN(DP_reg_a_i_1_n52) );
  NAND2_X1 DP_reg_a_i_2_U27 ( .A1(a[11]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n63) );
  OAI21_X1 DP_reg_a_i_2_U26 ( .B1(DP_reg_a_i_2_n37), .B2(DP_reg_a_i_2_n51), 
        .A(DP_reg_a_i_2_n63), .ZN(DP_reg_a_i_2_n39) );
  NAND2_X1 DP_reg_a_i_2_U25 ( .A1(a[10]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n64) );
  OAI21_X1 DP_reg_a_i_2_U24 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n52), 
        .A(DP_reg_a_i_2_n64), .ZN(DP_reg_a_i_2_n40) );
  NAND2_X1 DP_reg_a_i_2_U23 ( .A1(a[9]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n65) );
  OAI21_X1 DP_reg_a_i_2_U22 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n53), 
        .A(DP_reg_a_i_2_n65), .ZN(DP_reg_a_i_2_n41) );
  NAND2_X1 DP_reg_a_i_2_U21 ( .A1(a[8]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n66) );
  OAI21_X1 DP_reg_a_i_2_U20 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n54), 
        .A(DP_reg_a_i_2_n66), .ZN(DP_reg_a_i_2_n42) );
  NAND2_X1 DP_reg_a_i_2_U19 ( .A1(a[7]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n67) );
  OAI21_X1 DP_reg_a_i_2_U18 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n55), 
        .A(DP_reg_a_i_2_n67), .ZN(DP_reg_a_i_2_n43) );
  NAND2_X1 DP_reg_a_i_2_U17 ( .A1(a[6]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n68) );
  OAI21_X1 DP_reg_a_i_2_U16 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n56), 
        .A(DP_reg_a_i_2_n68), .ZN(DP_reg_a_i_2_n44) );
  NAND2_X1 DP_reg_a_i_2_U15 ( .A1(a[5]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n69) );
  OAI21_X1 DP_reg_a_i_2_U14 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n57), 
        .A(DP_reg_a_i_2_n69), .ZN(DP_reg_a_i_2_n45) );
  NAND2_X1 DP_reg_a_i_2_U13 ( .A1(a[4]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n70) );
  OAI21_X1 DP_reg_a_i_2_U12 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n58), 
        .A(DP_reg_a_i_2_n70), .ZN(DP_reg_a_i_2_n46) );
  NAND2_X1 DP_reg_a_i_2_U11 ( .A1(a[3]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n71) );
  OAI21_X1 DP_reg_a_i_2_U10 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n59), 
        .A(DP_reg_a_i_2_n71), .ZN(DP_reg_a_i_2_n47) );
  NAND2_X1 DP_reg_a_i_2_U9 ( .A1(a[2]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n72) );
  OAI21_X1 DP_reg_a_i_2_U8 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n60), .A(
        DP_reg_a_i_2_n72), .ZN(DP_reg_a_i_2_n48) );
  NAND2_X1 DP_reg_a_i_2_U7 ( .A1(a[1]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n73) );
  OAI21_X1 DP_reg_a_i_2_U6 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n61), .A(
        DP_reg_a_i_2_n73), .ZN(DP_reg_a_i_2_n49) );
  NAND2_X1 DP_reg_a_i_2_U5 ( .A1(DP_reg_a_i_2_n38), .A2(a[0]), .ZN(
        DP_reg_a_i_2_n74) );
  OAI21_X1 DP_reg_a_i_2_U4 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n62), .A(
        DP_reg_a_i_2_n74), .ZN(DP_reg_a_i_2_n50) );
  BUF_X1 DP_reg_a_i_2_U3 ( .A(vIn), .Z(DP_reg_a_i_2_n38) );
  BUF_X1 DP_reg_a_i_2_U2 ( .A(vIn), .Z(DP_reg_a_i_2_n37) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_0_ ( .D(DP_reg_a_i_2_n50), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[23]), .QN(DP_reg_a_i_2_n62) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_11_ ( .D(DP_reg_a_i_2_n39), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[12]), .QN(DP_reg_a_i_2_n51) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_1_ ( .D(DP_reg_a_i_2_n49), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[22]), .QN(DP_reg_a_i_2_n61) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_2_ ( .D(DP_reg_a_i_2_n48), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[21]), .QN(DP_reg_a_i_2_n60) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_3_ ( .D(DP_reg_a_i_2_n47), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[20]), .QN(DP_reg_a_i_2_n59) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_4_ ( .D(DP_reg_a_i_2_n46), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[19]), .QN(DP_reg_a_i_2_n58) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_5_ ( .D(DP_reg_a_i_2_n45), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[18]), .QN(DP_reg_a_i_2_n57) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_6_ ( .D(DP_reg_a_i_2_n44), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[17]), .QN(DP_reg_a_i_2_n56) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_7_ ( .D(DP_reg_a_i_2_n43), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[16]), .QN(DP_reg_a_i_2_n55) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_8_ ( .D(DP_reg_a_i_2_n42), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[15]), .QN(DP_reg_a_i_2_n54) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_9_ ( .D(DP_reg_a_i_2_n41), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[14]), .QN(DP_reg_a_i_2_n53) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_10_ ( .D(DP_reg_a_i_2_n40), .CK(clk), .RN(DP_n3), 
        .Q(DP_a_int[13]), .QN(DP_reg_a_i_2_n52) );
  NAND2_X1 DP_reg_b_i_0_U27 ( .A1(b[35]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n63) );
  OAI21_X1 DP_reg_b_i_0_U26 ( .B1(DP_reg_b_i_0_n37), .B2(DP_reg_b_i_0_n51), 
        .A(DP_reg_b_i_0_n63), .ZN(DP_reg_b_i_0_n39) );
  NAND2_X1 DP_reg_b_i_0_U25 ( .A1(b[34]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n64) );
  OAI21_X1 DP_reg_b_i_0_U24 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n52), 
        .A(DP_reg_b_i_0_n64), .ZN(DP_reg_b_i_0_n40) );
  NAND2_X1 DP_reg_b_i_0_U23 ( .A1(b[33]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n65) );
  OAI21_X1 DP_reg_b_i_0_U22 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n53), 
        .A(DP_reg_b_i_0_n65), .ZN(DP_reg_b_i_0_n41) );
  NAND2_X1 DP_reg_b_i_0_U21 ( .A1(b[32]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n66) );
  OAI21_X1 DP_reg_b_i_0_U20 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n54), 
        .A(DP_reg_b_i_0_n66), .ZN(DP_reg_b_i_0_n42) );
  NAND2_X1 DP_reg_b_i_0_U19 ( .A1(b[31]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n67) );
  OAI21_X1 DP_reg_b_i_0_U18 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n55), 
        .A(DP_reg_b_i_0_n67), .ZN(DP_reg_b_i_0_n43) );
  NAND2_X1 DP_reg_b_i_0_U17 ( .A1(b[30]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n68) );
  OAI21_X1 DP_reg_b_i_0_U16 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n56), 
        .A(DP_reg_b_i_0_n68), .ZN(DP_reg_b_i_0_n44) );
  NAND2_X1 DP_reg_b_i_0_U15 ( .A1(b[29]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n69) );
  OAI21_X1 DP_reg_b_i_0_U14 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n57), 
        .A(DP_reg_b_i_0_n69), .ZN(DP_reg_b_i_0_n45) );
  NAND2_X1 DP_reg_b_i_0_U13 ( .A1(b[28]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n70) );
  OAI21_X1 DP_reg_b_i_0_U12 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n58), 
        .A(DP_reg_b_i_0_n70), .ZN(DP_reg_b_i_0_n46) );
  NAND2_X1 DP_reg_b_i_0_U11 ( .A1(b[27]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n71) );
  OAI21_X1 DP_reg_b_i_0_U10 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n59), 
        .A(DP_reg_b_i_0_n71), .ZN(DP_reg_b_i_0_n47) );
  NAND2_X1 DP_reg_b_i_0_U9 ( .A1(b[26]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n72) );
  OAI21_X1 DP_reg_b_i_0_U8 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n60), .A(
        DP_reg_b_i_0_n72), .ZN(DP_reg_b_i_0_n48) );
  NAND2_X1 DP_reg_b_i_0_U7 ( .A1(b[25]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n73) );
  OAI21_X1 DP_reg_b_i_0_U6 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n61), .A(
        DP_reg_b_i_0_n73), .ZN(DP_reg_b_i_0_n49) );
  NAND2_X1 DP_reg_b_i_0_U5 ( .A1(DP_reg_b_i_0_n38), .A2(b[24]), .ZN(
        DP_reg_b_i_0_n74) );
  OAI21_X1 DP_reg_b_i_0_U4 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n62), .A(
        DP_reg_b_i_0_n74), .ZN(DP_reg_b_i_0_n50) );
  BUF_X1 DP_reg_b_i_0_U3 ( .A(vIn), .Z(DP_reg_b_i_0_n38) );
  BUF_X1 DP_reg_b_i_0_U2 ( .A(vIn), .Z(DP_reg_b_i_0_n37) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_0_ ( .D(DP_reg_b_i_0_n50), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[11]), .QN(DP_reg_b_i_0_n62) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_11_ ( .D(DP_reg_b_i_0_n39), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[0]), .QN(DP_reg_b_i_0_n51) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_1_ ( .D(DP_reg_b_i_0_n49), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[10]), .QN(DP_reg_b_i_0_n61) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_2_ ( .D(DP_reg_b_i_0_n48), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[9]), .QN(DP_reg_b_i_0_n60) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_3_ ( .D(DP_reg_b_i_0_n47), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[8]), .QN(DP_reg_b_i_0_n59) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_4_ ( .D(DP_reg_b_i_0_n46), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[7]), .QN(DP_reg_b_i_0_n58) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_5_ ( .D(DP_reg_b_i_0_n45), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[6]), .QN(DP_reg_b_i_0_n57) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_6_ ( .D(DP_reg_b_i_0_n44), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[5]), .QN(DP_reg_b_i_0_n56) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_7_ ( .D(DP_reg_b_i_0_n43), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[4]), .QN(DP_reg_b_i_0_n55) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_8_ ( .D(DP_reg_b_i_0_n42), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[3]), .QN(DP_reg_b_i_0_n54) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_9_ ( .D(DP_reg_b_i_0_n41), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[2]), .QN(DP_reg_b_i_0_n53) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_10_ ( .D(DP_reg_b_i_0_n40), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[1]), .QN(DP_reg_b_i_0_n52) );
  NAND2_X1 DP_reg_b_i_1_U27 ( .A1(b[23]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n63) );
  OAI21_X1 DP_reg_b_i_1_U26 ( .B1(DP_reg_b_i_1_n37), .B2(DP_reg_b_i_1_n51), 
        .A(DP_reg_b_i_1_n63), .ZN(DP_reg_b_i_1_n39) );
  NAND2_X1 DP_reg_b_i_1_U25 ( .A1(b[22]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n64) );
  OAI21_X1 DP_reg_b_i_1_U24 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n52), 
        .A(DP_reg_b_i_1_n64), .ZN(DP_reg_b_i_1_n40) );
  NAND2_X1 DP_reg_b_i_1_U23 ( .A1(b[21]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n65) );
  OAI21_X1 DP_reg_b_i_1_U22 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n53), 
        .A(DP_reg_b_i_1_n65), .ZN(DP_reg_b_i_1_n41) );
  NAND2_X1 DP_reg_b_i_1_U21 ( .A1(b[20]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n66) );
  OAI21_X1 DP_reg_b_i_1_U20 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n54), 
        .A(DP_reg_b_i_1_n66), .ZN(DP_reg_b_i_1_n42) );
  NAND2_X1 DP_reg_b_i_1_U19 ( .A1(b[19]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n67) );
  OAI21_X1 DP_reg_b_i_1_U18 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n55), 
        .A(DP_reg_b_i_1_n67), .ZN(DP_reg_b_i_1_n43) );
  NAND2_X1 DP_reg_b_i_1_U17 ( .A1(b[18]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n68) );
  OAI21_X1 DP_reg_b_i_1_U16 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n56), 
        .A(DP_reg_b_i_1_n68), .ZN(DP_reg_b_i_1_n44) );
  NAND2_X1 DP_reg_b_i_1_U15 ( .A1(b[17]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n69) );
  OAI21_X1 DP_reg_b_i_1_U14 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n57), 
        .A(DP_reg_b_i_1_n69), .ZN(DP_reg_b_i_1_n45) );
  NAND2_X1 DP_reg_b_i_1_U13 ( .A1(b[16]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n70) );
  OAI21_X1 DP_reg_b_i_1_U12 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n58), 
        .A(DP_reg_b_i_1_n70), .ZN(DP_reg_b_i_1_n46) );
  NAND2_X1 DP_reg_b_i_1_U11 ( .A1(b[15]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n71) );
  OAI21_X1 DP_reg_b_i_1_U10 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n59), 
        .A(DP_reg_b_i_1_n71), .ZN(DP_reg_b_i_1_n47) );
  NAND2_X1 DP_reg_b_i_1_U9 ( .A1(b[14]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n72) );
  OAI21_X1 DP_reg_b_i_1_U8 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n60), .A(
        DP_reg_b_i_1_n72), .ZN(DP_reg_b_i_1_n48) );
  NAND2_X1 DP_reg_b_i_1_U7 ( .A1(b[13]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n73) );
  OAI21_X1 DP_reg_b_i_1_U6 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n61), .A(
        DP_reg_b_i_1_n73), .ZN(DP_reg_b_i_1_n49) );
  NAND2_X1 DP_reg_b_i_1_U5 ( .A1(DP_reg_b_i_1_n38), .A2(b[12]), .ZN(
        DP_reg_b_i_1_n74) );
  OAI21_X1 DP_reg_b_i_1_U4 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n62), .A(
        DP_reg_b_i_1_n74), .ZN(DP_reg_b_i_1_n50) );
  BUF_X1 DP_reg_b_i_1_U3 ( .A(vIn), .Z(DP_reg_b_i_1_n38) );
  BUF_X1 DP_reg_b_i_1_U2 ( .A(vIn), .Z(DP_reg_b_i_1_n37) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_0_ ( .D(DP_reg_b_i_1_n50), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[23]), .QN(DP_reg_b_i_1_n62) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_11_ ( .D(DP_reg_b_i_1_n39), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[12]), .QN(DP_reg_b_i_1_n51) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_1_ ( .D(DP_reg_b_i_1_n49), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[22]), .QN(DP_reg_b_i_1_n61) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_2_ ( .D(DP_reg_b_i_1_n48), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[21]), .QN(DP_reg_b_i_1_n60) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_3_ ( .D(DP_reg_b_i_1_n47), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[20]), .QN(DP_reg_b_i_1_n59) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_4_ ( .D(DP_reg_b_i_1_n46), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[19]), .QN(DP_reg_b_i_1_n58) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_5_ ( .D(DP_reg_b_i_1_n45), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[18]), .QN(DP_reg_b_i_1_n57) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_6_ ( .D(DP_reg_b_i_1_n44), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[17]), .QN(DP_reg_b_i_1_n56) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_7_ ( .D(DP_reg_b_i_1_n43), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[16]), .QN(DP_reg_b_i_1_n55) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_8_ ( .D(DP_reg_b_i_1_n42), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[15]), .QN(DP_reg_b_i_1_n54) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_9_ ( .D(DP_reg_b_i_1_n41), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[14]), .QN(DP_reg_b_i_1_n53) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_10_ ( .D(DP_reg_b_i_1_n40), .CK(clk), .RN(DP_n3), 
        .Q(DP_b_int[13]), .QN(DP_reg_b_i_1_n52) );
  NAND2_X1 DP_reg_b_i_2_U27 ( .A1(b[11]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n63) );
  OAI21_X1 DP_reg_b_i_2_U26 ( .B1(DP_reg_b_i_2_n37), .B2(DP_reg_b_i_2_n51), 
        .A(DP_reg_b_i_2_n63), .ZN(DP_reg_b_i_2_n39) );
  NAND2_X1 DP_reg_b_i_2_U25 ( .A1(b[10]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n64) );
  OAI21_X1 DP_reg_b_i_2_U24 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n52), 
        .A(DP_reg_b_i_2_n64), .ZN(DP_reg_b_i_2_n40) );
  NAND2_X1 DP_reg_b_i_2_U23 ( .A1(b[9]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n65) );
  OAI21_X1 DP_reg_b_i_2_U22 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n53), 
        .A(DP_reg_b_i_2_n65), .ZN(DP_reg_b_i_2_n41) );
  NAND2_X1 DP_reg_b_i_2_U21 ( .A1(b[8]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n66) );
  OAI21_X1 DP_reg_b_i_2_U20 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n54), 
        .A(DP_reg_b_i_2_n66), .ZN(DP_reg_b_i_2_n42) );
  NAND2_X1 DP_reg_b_i_2_U19 ( .A1(b[7]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n67) );
  OAI21_X1 DP_reg_b_i_2_U18 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n55), 
        .A(DP_reg_b_i_2_n67), .ZN(DP_reg_b_i_2_n43) );
  NAND2_X1 DP_reg_b_i_2_U17 ( .A1(b[6]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n68) );
  OAI21_X1 DP_reg_b_i_2_U16 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n56), 
        .A(DP_reg_b_i_2_n68), .ZN(DP_reg_b_i_2_n44) );
  NAND2_X1 DP_reg_b_i_2_U15 ( .A1(b[5]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n69) );
  OAI21_X1 DP_reg_b_i_2_U14 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n57), 
        .A(DP_reg_b_i_2_n69), .ZN(DP_reg_b_i_2_n45) );
  NAND2_X1 DP_reg_b_i_2_U13 ( .A1(b[4]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n70) );
  OAI21_X1 DP_reg_b_i_2_U12 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n58), 
        .A(DP_reg_b_i_2_n70), .ZN(DP_reg_b_i_2_n46) );
  NAND2_X1 DP_reg_b_i_2_U11 ( .A1(b[3]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n71) );
  OAI21_X1 DP_reg_b_i_2_U10 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n59), 
        .A(DP_reg_b_i_2_n71), .ZN(DP_reg_b_i_2_n47) );
  NAND2_X1 DP_reg_b_i_2_U9 ( .A1(b[2]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n72) );
  OAI21_X1 DP_reg_b_i_2_U8 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n60), .A(
        DP_reg_b_i_2_n72), .ZN(DP_reg_b_i_2_n48) );
  NAND2_X1 DP_reg_b_i_2_U7 ( .A1(b[1]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n73) );
  OAI21_X1 DP_reg_b_i_2_U6 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n61), .A(
        DP_reg_b_i_2_n73), .ZN(DP_reg_b_i_2_n49) );
  NAND2_X1 DP_reg_b_i_2_U5 ( .A1(DP_reg_b_i_2_n38), .A2(b[0]), .ZN(
        DP_reg_b_i_2_n74) );
  OAI21_X1 DP_reg_b_i_2_U4 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n62), .A(
        DP_reg_b_i_2_n74), .ZN(DP_reg_b_i_2_n50) );
  BUF_X1 DP_reg_b_i_2_U3 ( .A(vIn), .Z(DP_reg_b_i_2_n38) );
  BUF_X1 DP_reg_b_i_2_U2 ( .A(vIn), .Z(DP_reg_b_i_2_n37) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_0_ ( .D(DP_reg_b_i_2_n50), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[35]), .QN(DP_reg_b_i_2_n62) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_11_ ( .D(DP_reg_b_i_2_n39), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[24]), .QN(DP_reg_b_i_2_n51) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_1_ ( .D(DP_reg_b_i_2_n49), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[34]), .QN(DP_reg_b_i_2_n61) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_2_ ( .D(DP_reg_b_i_2_n48), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[33]), .QN(DP_reg_b_i_2_n60) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_3_ ( .D(DP_reg_b_i_2_n47), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[32]), .QN(DP_reg_b_i_2_n59) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_4_ ( .D(DP_reg_b_i_2_n46), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[31]), .QN(DP_reg_b_i_2_n58) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_5_ ( .D(DP_reg_b_i_2_n45), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[30]), .QN(DP_reg_b_i_2_n57) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_6_ ( .D(DP_reg_b_i_2_n44), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[29]), .QN(DP_reg_b_i_2_n56) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_7_ ( .D(DP_reg_b_i_2_n43), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[28]), .QN(DP_reg_b_i_2_n55) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_8_ ( .D(DP_reg_b_i_2_n42), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[27]), .QN(DP_reg_b_i_2_n54) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_9_ ( .D(DP_reg_b_i_2_n41), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[26]), .QN(DP_reg_b_i_2_n53) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_10_ ( .D(DP_reg_b_i_2_n40), .CK(clk), .RN(DP_n2), 
        .Q(DP_b_int[25]), .QN(DP_reg_b_i_2_n52) );
  NAND2_X1 DP_reg_sw0_U30 ( .A1(sw_out_regs_en_int), .A2(DP_w_0_), .ZN(
        DP_reg_sw0_n1) );
  OAI21_X1 DP_reg_sw0_U29 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n14), .A(
        DP_reg_sw0_n1), .ZN(DP_reg_sw0_n27) );
  NAND2_X1 DP_reg_sw0_U28 ( .A1(DP_w_10_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n11) );
  OAI21_X1 DP_reg_sw0_U27 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n24), .A(
        DP_reg_sw0_n11), .ZN(DP_reg_sw0_n37) );
  NAND2_X1 DP_reg_sw0_U26 ( .A1(DP_w_7_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n8) );
  OAI21_X1 DP_reg_sw0_U25 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n21), .A(
        DP_reg_sw0_n8), .ZN(DP_reg_sw0_n34) );
  NAND2_X1 DP_reg_sw0_U24 ( .A1(DP_w_4_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n5) );
  OAI21_X1 DP_reg_sw0_U23 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n18), .A(
        DP_reg_sw0_n5), .ZN(DP_reg_sw0_n31) );
  NAND2_X1 DP_reg_sw0_U22 ( .A1(DP_w_3_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n4) );
  OAI21_X1 DP_reg_sw0_U21 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n17), .A(
        DP_reg_sw0_n4), .ZN(DP_reg_sw0_n30) );
  NAND2_X1 DP_reg_sw0_U20 ( .A1(DP_w_1_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n2) );
  OAI21_X1 DP_reg_sw0_U19 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n15), .A(
        DP_reg_sw0_n2), .ZN(DP_reg_sw0_n28) );
  NAND2_X1 DP_reg_sw0_U18 ( .A1(DP_w_9_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n10) );
  OAI21_X1 DP_reg_sw0_U17 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n23), .A(
        DP_reg_sw0_n10), .ZN(DP_reg_sw0_n36) );
  NAND2_X1 DP_reg_sw0_U16 ( .A1(DP_w_8_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n9) );
  OAI21_X1 DP_reg_sw0_U15 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n22), .A(
        DP_reg_sw0_n9), .ZN(DP_reg_sw0_n35) );
  NAND2_X1 DP_reg_sw0_U14 ( .A1(DP_w_6_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n7) );
  OAI21_X1 DP_reg_sw0_U13 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n20), .A(
        DP_reg_sw0_n7), .ZN(DP_reg_sw0_n33) );
  NAND2_X1 DP_reg_sw0_U12 ( .A1(DP_w_5_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n6) );
  OAI21_X1 DP_reg_sw0_U11 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n19), .A(
        DP_reg_sw0_n6), .ZN(DP_reg_sw0_n32) );
  NAND2_X1 DP_reg_sw0_U10 ( .A1(DP_w_2_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n3) );
  OAI21_X1 DP_reg_sw0_U9 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n16), .A(
        DP_reg_sw0_n3), .ZN(DP_reg_sw0_n29) );
  NAND2_X1 DP_reg_sw0_U8 ( .A1(DP_w_11_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n12) );
  OAI21_X1 DP_reg_sw0_U7 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n25), .A(
        DP_reg_sw0_n12), .ZN(DP_reg_sw0_n38) );
  NAND2_X1 DP_reg_sw0_U6 ( .A1(DP_w_12_), .A2(DP_reg_sw0_n40), .ZN(
        DP_reg_sw0_n13) );
  OAI21_X1 DP_reg_sw0_U5 ( .B1(DP_reg_sw0_n41), .B2(DP_reg_sw0_n26), .A(
        DP_reg_sw0_n13), .ZN(DP_reg_sw0_n39) );
  BUF_X1 DP_reg_sw0_U4 ( .A(DP_n1), .Z(DP_reg_sw0_n42) );
  BUF_X1 DP_reg_sw0_U3 ( .A(sw_out_regs_en_int), .Z(DP_reg_sw0_n41) );
  BUF_X1 DP_reg_sw0_U2 ( .A(sw_out_regs_en_int), .Z(DP_reg_sw0_n40) );
  DFFR_X1 DP_reg_sw0_Q_reg_0_ ( .D(DP_reg_sw0_n27), .CK(clk), .RN(DP_n1), .Q(
        DP_sw0_0_), .QN(DP_reg_sw0_n14) );
  DFFR_X1 DP_reg_sw0_Q_reg_1_ ( .D(DP_reg_sw0_n28), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_1_), .QN(DP_reg_sw0_n15) );
  DFFR_X1 DP_reg_sw0_Q_reg_2_ ( .D(DP_reg_sw0_n29), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_2_), .QN(DP_reg_sw0_n16) );
  DFFR_X1 DP_reg_sw0_Q_reg_3_ ( .D(DP_reg_sw0_n30), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_3_), .QN(DP_reg_sw0_n17) );
  DFFR_X1 DP_reg_sw0_Q_reg_4_ ( .D(DP_reg_sw0_n31), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_4_), .QN(DP_reg_sw0_n18) );
  DFFR_X1 DP_reg_sw0_Q_reg_5_ ( .D(DP_reg_sw0_n32), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_5_), .QN(DP_reg_sw0_n19) );
  DFFR_X1 DP_reg_sw0_Q_reg_6_ ( .D(DP_reg_sw0_n33), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_6_), .QN(DP_reg_sw0_n20) );
  DFFR_X1 DP_reg_sw0_Q_reg_7_ ( .D(DP_reg_sw0_n34), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_7_), .QN(DP_reg_sw0_n21) );
  DFFR_X1 DP_reg_sw0_Q_reg_8_ ( .D(DP_reg_sw0_n35), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_8_), .QN(DP_reg_sw0_n22) );
  DFFR_X1 DP_reg_sw0_Q_reg_9_ ( .D(DP_reg_sw0_n36), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_9_), .QN(DP_reg_sw0_n23) );
  DFFR_X1 DP_reg_sw0_Q_reg_10_ ( .D(DP_reg_sw0_n37), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_10_), .QN(DP_reg_sw0_n24) );
  DFFR_X1 DP_reg_sw0_Q_reg_11_ ( .D(DP_reg_sw0_n38), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_11_), .QN(DP_reg_sw0_n25) );
  DFFR_X1 DP_reg_sw0_Q_reg_12_ ( .D(DP_reg_sw0_n39), .CK(clk), .RN(
        DP_reg_sw0_n42), .Q(DP_sw0_12_), .QN(DP_reg_sw0_n26) );
  NAND2_X1 DP_reg_sw1_U29 ( .A1(DP_sw0_12_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n68) );
  OAI21_X1 DP_reg_sw1_U28 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n55), .A(
        DP_reg_sw1_n68), .ZN(DP_reg_sw1_n42) );
  NAND2_X1 DP_reg_sw1_U27 ( .A1(DP_sw0_11_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n69) );
  OAI21_X1 DP_reg_sw1_U26 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n56), .A(
        DP_reg_sw1_n69), .ZN(DP_reg_sw1_n43) );
  NAND2_X1 DP_reg_sw1_U25 ( .A1(DP_sw0_10_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n70) );
  OAI21_X1 DP_reg_sw1_U24 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n57), .A(
        DP_reg_sw1_n70), .ZN(DP_reg_sw1_n44) );
  NAND2_X1 DP_reg_sw1_U23 ( .A1(DP_sw0_9_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n71) );
  OAI21_X1 DP_reg_sw1_U22 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n58), .A(
        DP_reg_sw1_n71), .ZN(DP_reg_sw1_n45) );
  NAND2_X1 DP_reg_sw1_U21 ( .A1(DP_sw0_8_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n72) );
  OAI21_X1 DP_reg_sw1_U20 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n59), .A(
        DP_reg_sw1_n72), .ZN(DP_reg_sw1_n46) );
  NAND2_X1 DP_reg_sw1_U19 ( .A1(DP_sw0_7_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n73) );
  OAI21_X1 DP_reg_sw1_U18 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n60), .A(
        DP_reg_sw1_n73), .ZN(DP_reg_sw1_n47) );
  NAND2_X1 DP_reg_sw1_U17 ( .A1(DP_sw0_6_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n74) );
  OAI21_X1 DP_reg_sw1_U16 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n61), .A(
        DP_reg_sw1_n74), .ZN(DP_reg_sw1_n48) );
  NAND2_X1 DP_reg_sw1_U15 ( .A1(DP_sw0_5_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n75) );
  OAI21_X1 DP_reg_sw1_U14 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n62), .A(
        DP_reg_sw1_n75), .ZN(DP_reg_sw1_n49) );
  NAND2_X1 DP_reg_sw1_U13 ( .A1(DP_sw0_4_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n76) );
  OAI21_X1 DP_reg_sw1_U12 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n63), .A(
        DP_reg_sw1_n76), .ZN(DP_reg_sw1_n50) );
  NAND2_X1 DP_reg_sw1_U11 ( .A1(DP_sw0_3_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n77) );
  OAI21_X1 DP_reg_sw1_U10 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n64), .A(
        DP_reg_sw1_n77), .ZN(DP_reg_sw1_n51) );
  NAND2_X1 DP_reg_sw1_U9 ( .A1(DP_sw0_2_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n78) );
  OAI21_X1 DP_reg_sw1_U8 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n65), .A(
        DP_reg_sw1_n78), .ZN(DP_reg_sw1_n52) );
  NAND2_X1 DP_reg_sw1_U7 ( .A1(DP_sw0_1_), .A2(DP_reg_sw1_n40), .ZN(
        DP_reg_sw1_n79) );
  OAI21_X1 DP_reg_sw1_U6 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n66), .A(
        DP_reg_sw1_n79), .ZN(DP_reg_sw1_n53) );
  NAND2_X1 DP_reg_sw1_U5 ( .A1(DP_reg_sw1_n41), .A2(DP_sw0_0_), .ZN(
        DP_reg_sw1_n80) );
  OAI21_X1 DP_reg_sw1_U4 ( .B1(DP_reg_sw1_n41), .B2(DP_reg_sw1_n67), .A(
        DP_reg_sw1_n80), .ZN(DP_reg_sw1_n54) );
  BUF_X1 DP_reg_sw1_U3 ( .A(sw_out_regs_en_int), .Z(DP_reg_sw1_n41) );
  BUF_X1 DP_reg_sw1_U2 ( .A(sw_out_regs_en_int), .Z(DP_reg_sw1_n40) );
  DFFR_X1 DP_reg_sw1_Q_reg_2_ ( .D(DP_reg_sw1_n52), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_2_), .QN(DP_reg_sw1_n65) );
  DFFR_X1 DP_reg_sw1_Q_reg_3_ ( .D(DP_reg_sw1_n51), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_3_), .QN(DP_reg_sw1_n64) );
  DFFR_X1 DP_reg_sw1_Q_reg_4_ ( .D(DP_reg_sw1_n50), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_4_), .QN(DP_reg_sw1_n63) );
  DFFR_X1 DP_reg_sw1_Q_reg_5_ ( .D(DP_reg_sw1_n49), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_5_), .QN(DP_reg_sw1_n62) );
  DFFR_X1 DP_reg_sw1_Q_reg_6_ ( .D(DP_reg_sw1_n48), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_6_), .QN(DP_reg_sw1_n61) );
  DFFR_X1 DP_reg_sw1_Q_reg_7_ ( .D(DP_reg_sw1_n47), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_7_), .QN(DP_reg_sw1_n60) );
  DFFR_X1 DP_reg_sw1_Q_reg_8_ ( .D(DP_reg_sw1_n46), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_8_), .QN(DP_reg_sw1_n59) );
  DFFR_X1 DP_reg_sw1_Q_reg_9_ ( .D(DP_reg_sw1_n45), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_9_), .QN(DP_reg_sw1_n58) );
  DFFR_X1 DP_reg_sw1_Q_reg_10_ ( .D(DP_reg_sw1_n44), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_10_), .QN(DP_reg_sw1_n57) );
  DFFR_X1 DP_reg_sw1_Q_reg_11_ ( .D(DP_reg_sw1_n43), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_11_), .QN(DP_reg_sw1_n56) );
  DFFR_X1 DP_reg_sw1_Q_reg_12_ ( .D(DP_reg_sw1_n42), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_12_), .QN(DP_reg_sw1_n55) );
  DFFR_X1 DP_reg_sw1_Q_reg_1_ ( .D(DP_reg_sw1_n53), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_1_), .QN(DP_reg_sw1_n66) );
  DFFR_X1 DP_reg_sw1_Q_reg_0_ ( .D(DP_reg_sw1_n54), .CK(clk), .RN(DP_n1), .Q(
        DP_sw1_0_), .QN(DP_reg_sw1_n67) );
  NAND2_X1 DP_reg_out_U27 ( .A1(DP_reg_out_n38), .A2(DP_y_out_0_), .ZN(
        DP_reg_out_n74) );
  OAI21_X1 DP_reg_out_U26 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n62), .A(
        DP_reg_out_n74), .ZN(DP_reg_out_n50) );
  NAND2_X1 DP_reg_out_U25 ( .A1(DP_y_out_10_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n64) );
  OAI21_X1 DP_reg_out_U24 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n52), .A(
        DP_reg_out_n64), .ZN(DP_reg_out_n40) );
  NAND2_X1 DP_reg_out_U23 ( .A1(DP_y_out_9_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n65) );
  OAI21_X1 DP_reg_out_U22 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n53), .A(
        DP_reg_out_n65), .ZN(DP_reg_out_n41) );
  NAND2_X1 DP_reg_out_U21 ( .A1(DP_y_out_8_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n66) );
  OAI21_X1 DP_reg_out_U20 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n54), .A(
        DP_reg_out_n66), .ZN(DP_reg_out_n42) );
  NAND2_X1 DP_reg_out_U19 ( .A1(DP_y_out_7_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n67) );
  OAI21_X1 DP_reg_out_U18 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n55), .A(
        DP_reg_out_n67), .ZN(DP_reg_out_n43) );
  NAND2_X1 DP_reg_out_U17 ( .A1(DP_y_out_6_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n68) );
  OAI21_X1 DP_reg_out_U16 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n56), .A(
        DP_reg_out_n68), .ZN(DP_reg_out_n44) );
  NAND2_X1 DP_reg_out_U15 ( .A1(DP_y_out_5_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n69) );
  OAI21_X1 DP_reg_out_U14 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n57), .A(
        DP_reg_out_n69), .ZN(DP_reg_out_n45) );
  NAND2_X1 DP_reg_out_U13 ( .A1(DP_y_out_4_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n70) );
  OAI21_X1 DP_reg_out_U12 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n58), .A(
        DP_reg_out_n70), .ZN(DP_reg_out_n46) );
  NAND2_X1 DP_reg_out_U11 ( .A1(DP_y_out_3_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n71) );
  OAI21_X1 DP_reg_out_U10 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n59), .A(
        DP_reg_out_n71), .ZN(DP_reg_out_n47) );
  NAND2_X1 DP_reg_out_U9 ( .A1(DP_y_out_2_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n72) );
  OAI21_X1 DP_reg_out_U8 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n60), .A(
        DP_reg_out_n72), .ZN(DP_reg_out_n48) );
  NAND2_X1 DP_reg_out_U7 ( .A1(DP_y_out_1_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n73) );
  OAI21_X1 DP_reg_out_U6 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n61), .A(
        DP_reg_out_n73), .ZN(DP_reg_out_n49) );
  NAND2_X1 DP_reg_out_U5 ( .A1(DP_y_out_11_), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n63) );
  OAI21_X1 DP_reg_out_U4 ( .B1(DP_reg_out_n37), .B2(DP_reg_out_n51), .A(
        DP_reg_out_n63), .ZN(DP_reg_out_n39) );
  BUF_X1 DP_reg_out_U3 ( .A(sw_out_regs_en_int), .Z(DP_reg_out_n38) );
  BUF_X1 DP_reg_out_U2 ( .A(sw_out_regs_en_int), .Z(DP_reg_out_n37) );
  DFFR_X1 DP_reg_out_Q_reg_0_ ( .D(DP_reg_out_n50), .CK(clk), .RN(DP_n2), .Q(
        dOut[0]), .QN(DP_reg_out_n62) );
  DFFR_X1 DP_reg_out_Q_reg_1_ ( .D(DP_reg_out_n49), .CK(clk), .RN(DP_n2), .Q(
        dOut[1]), .QN(DP_reg_out_n61) );
  DFFR_X1 DP_reg_out_Q_reg_2_ ( .D(DP_reg_out_n48), .CK(clk), .RN(DP_n2), .Q(
        dOut[2]), .QN(DP_reg_out_n60) );
  DFFR_X1 DP_reg_out_Q_reg_3_ ( .D(DP_reg_out_n47), .CK(clk), .RN(DP_n2), .Q(
        dOut[3]), .QN(DP_reg_out_n59) );
  DFFR_X1 DP_reg_out_Q_reg_4_ ( .D(DP_reg_out_n46), .CK(clk), .RN(DP_n2), .Q(
        dOut[4]), .QN(DP_reg_out_n58) );
  DFFR_X1 DP_reg_out_Q_reg_5_ ( .D(DP_reg_out_n45), .CK(clk), .RN(DP_n2), .Q(
        dOut[5]), .QN(DP_reg_out_n57) );
  DFFR_X1 DP_reg_out_Q_reg_6_ ( .D(DP_reg_out_n44), .CK(clk), .RN(DP_n2), .Q(
        dOut[6]), .QN(DP_reg_out_n56) );
  DFFR_X1 DP_reg_out_Q_reg_7_ ( .D(DP_reg_out_n43), .CK(clk), .RN(DP_n2), .Q(
        dOut[7]), .QN(DP_reg_out_n55) );
  DFFR_X1 DP_reg_out_Q_reg_8_ ( .D(DP_reg_out_n42), .CK(clk), .RN(DP_n2), .Q(
        dOut[8]), .QN(DP_reg_out_n54) );
  DFFR_X1 DP_reg_out_Q_reg_9_ ( .D(DP_reg_out_n41), .CK(clk), .RN(DP_n2), .Q(
        dOut[9]), .QN(DP_reg_out_n53) );
  DFFR_X1 DP_reg_out_Q_reg_10_ ( .D(DP_reg_out_n40), .CK(clk), .RN(DP_n2), .Q(
        dOut[10]), .QN(DP_reg_out_n52) );
  DFFR_X1 DP_reg_out_Q_reg_11_ ( .D(DP_reg_out_n39), .CK(clk), .RN(DP_n2), .Q(
        dOut[11]), .QN(DP_reg_out_n51) );
  XOR2_X1 DP_add_1_root_add_0_root_add_107_U2 ( .A(DP_sw0_b1_0_), .B(
        DP_sw1_b2_0_), .Z(DP_ff_0_) );
  AND2_X1 DP_add_1_root_add_0_root_add_107_U1 ( .A1(DP_sw1_b2_0_), .A2(
        DP_sw0_b1_0_), .ZN(DP_add_1_root_add_0_root_add_107_carry_1_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_1 ( .A(DP_sw1_b2_1_), .B(
        DP_sw0_b1_1_), .CI(DP_add_1_root_add_0_root_add_107_carry_1_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_2_), .S(DP_ff_1_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_2 ( .A(DP_sw1_b2_2_), .B(
        DP_sw0_b1_2_), .CI(DP_add_1_root_add_0_root_add_107_carry_2_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_3_), .S(DP_ff_2_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_3 ( .A(DP_sw1_b2_3_), .B(
        DP_sw0_b1_3_), .CI(DP_add_1_root_add_0_root_add_107_carry_3_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_4_), .S(DP_ff_3_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_4 ( .A(DP_sw1_b2_4_), .B(
        DP_sw0_b1_4_), .CI(DP_add_1_root_add_0_root_add_107_carry_4_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_5_), .S(DP_ff_4_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_5 ( .A(DP_sw1_b2_5_), .B(
        DP_sw0_b1_5_), .CI(DP_add_1_root_add_0_root_add_107_carry_5_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_6_), .S(DP_ff_5_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_6 ( .A(DP_sw1_b2_6_), .B(
        DP_sw0_b1_6_), .CI(DP_add_1_root_add_0_root_add_107_carry_6_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_7_), .S(DP_ff_6_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_7 ( .A(DP_sw1_b2_7_), .B(
        DP_sw0_b1_7_), .CI(DP_add_1_root_add_0_root_add_107_carry_7_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_8_), .S(DP_ff_7_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_8 ( .A(DP_sw1_b2_8_), .B(
        DP_sw0_b1_8_), .CI(DP_add_1_root_add_0_root_add_107_carry_8_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_9_), .S(DP_ff_8_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_9 ( .A(DP_sw1_b2_9_), .B(
        DP_sw0_b1_9_), .CI(DP_add_1_root_add_0_root_add_107_carry_9_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_10_), .S(DP_ff_9_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_10 ( .A(DP_sw1_b2_10_), .B(
        DP_sw0_b1_10_), .CI(DP_add_1_root_add_0_root_add_107_carry_10_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_11_), .S(DP_ff_10_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_11 ( .A(DP_sw1_b2_11_), .B(
        DP_sw0_b1_11_), .CI(DP_add_1_root_add_0_root_add_107_carry_11_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_12_), .S(DP_ff_11_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_12 ( .A(DP_sw1_b2_11_), .B(
        DP_sw0_b1_11_), .CI(DP_add_1_root_add_0_root_add_107_carry_12_), .S(
        DP_ff_12_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U2 ( .A(DP_w_b0_0_), .B(DP_ff_0_), 
        .Z(DP_y[0]) );
  AND2_X1 DP_add_0_root_add_0_root_add_107_U1 ( .A1(DP_ff_0_), .A2(DP_w_b0_0_), 
        .ZN(DP_add_0_root_add_0_root_add_107_carry_1_) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_1 ( .A(DP_ff_1_), .B(DP_w_b0_1_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_1_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_2_), .S(DP_y[1]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_2 ( .A(DP_ff_2_), .B(DP_w_b0_2_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_2_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_3_), .S(DP_y[2]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_3 ( .A(DP_ff_3_), .B(DP_w_b0_3_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_3_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_4_), .S(DP_y[3]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_4 ( .A(DP_ff_4_), .B(DP_w_b0_4_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_4_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_5_), .S(DP_y[4]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_5 ( .A(DP_ff_5_), .B(DP_w_b0_5_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_5_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_6_), .S(DP_y[5]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_6 ( .A(DP_ff_6_), .B(DP_w_b0_6_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_6_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_7_), .S(DP_y[6]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_7 ( .A(DP_ff_7_), .B(DP_w_b0_7_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_7_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_8_), .S(DP_y[7]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_8 ( .A(DP_ff_8_), .B(DP_w_b0_8_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_8_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_9_), .S(DP_y[8]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_9 ( .A(DP_ff_9_), .B(DP_w_b0_9_), 
        .CI(DP_add_0_root_add_0_root_add_107_carry_9_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_10_), .S(DP_y[9]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_10 ( .A(DP_ff_10_), .B(DP_w_b0_10_), .CI(DP_add_0_root_add_0_root_add_107_carry_10_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_11_), .S(DP_y[10]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_11 ( .A(DP_ff_11_), .B(DP_w_b0_11_), .CI(DP_add_0_root_add_0_root_add_107_carry_11_), .CO(
        DP_add_0_root_add_0_root_add_107_carry_12_), .S(DP_y[11]) );
  FA_X1 DP_add_0_root_add_0_root_add_107_U1_12 ( .A(DP_ff_12_), .B(DP_w_b0_11_), .CI(DP_add_0_root_add_0_root_add_107_carry_12_), .S(DP_y_out_11_) );
  XOR2_X1 DP_mult_105_U563 ( .A(DP_b_int[9]), .B(DP_b_int[10]), .Z(
        DP_mult_105_n653) );
  INV_X1 DP_mult_105_U562 ( .A(DP_b_int[10]), .ZN(DP_mult_105_n543) );
  NOR2_X1 DP_mult_105_U561 ( .A1(DP_mult_105_n543), .A2(DP_w_1_), .ZN(
        DP_mult_105_n658) );
  INV_X1 DP_mult_105_U560 ( .A(DP_mult_105_n658), .ZN(DP_mult_105_n660) );
  NAND2_X1 DP_mult_105_U559 ( .A1(DP_b_int[10]), .A2(DP_mult_105_n532), .ZN(
        DP_mult_105_n530) );
  XNOR2_X1 DP_mult_105_U558 ( .A(DP_w_2_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n529) );
  OAI22_X1 DP_mult_105_U557 ( .A1(DP_mult_105_n660), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n529), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n659) );
  NAND2_X1 DP_mult_105_U556 ( .A1(DP_mult_105_n653), .A2(DP_mult_105_n659), 
        .ZN(DP_mult_105_n656) );
  NAND2_X1 DP_mult_105_U555 ( .A1(DP_mult_105_n658), .A2(DP_mult_105_n659), 
        .ZN(DP_mult_105_n657) );
  INV_X1 DP_mult_105_U554 ( .A(DP_w_0_), .ZN(DP_mult_105_n560) );
  MUX2_X1 DP_mult_105_U553 ( .A(DP_mult_105_n656), .B(DP_mult_105_n657), .S(
        DP_mult_105_n560), .Z(DP_mult_105_n655) );
  INV_X1 DP_mult_105_U552 ( .A(DP_mult_105_n655), .ZN(DP_mult_105_n650) );
  INV_X1 DP_mult_105_U551 ( .A(DP_b_int[8]), .ZN(DP_mult_105_n632) );
  XNOR2_X1 DP_mult_105_U550 ( .A(DP_mult_105_n632), .B(DP_b_int[9]), .ZN(
        DP_mult_105_n654) );
  NAND2_X1 DP_mult_105_U549 ( .A1(DP_mult_105_n546), .A2(DP_mult_105_n654), 
        .ZN(DP_mult_105_n545) );
  NAND3_X1 DP_mult_105_U548 ( .A1(DP_mult_105_n653), .A2(DP_mult_105_n560), 
        .A3(DP_b_int[8]), .ZN(DP_mult_105_n652) );
  OAI21_X1 DP_mult_105_U547 ( .B1(DP_mult_105_n632), .B2(DP_mult_105_n545), 
        .A(DP_mult_105_n652), .ZN(DP_mult_105_n651) );
  AOI222_X1 DP_mult_105_U546 ( .A1(DP_mult_105_n650), .A2(DP_mult_105_n255), 
        .B1(DP_mult_105_n651), .B2(DP_mult_105_n650), .C1(DP_mult_105_n651), 
        .C2(DP_mult_105_n255), .ZN(DP_mult_105_n649) );
  INV_X1 DP_mult_105_U545 ( .A(DP_mult_105_n649), .ZN(DP_mult_105_n648) );
  AOI222_X1 DP_mult_105_U544 ( .A1(DP_mult_105_n648), .A2(DP_mult_105_n253), 
        .B1(DP_mult_105_n648), .B2(DP_mult_105_n254), .C1(DP_mult_105_n254), 
        .C2(DP_mult_105_n253), .ZN(DP_mult_105_n647) );
  INV_X1 DP_mult_105_U543 ( .A(DP_mult_105_n647), .ZN(DP_mult_105_n646) );
  AOI222_X1 DP_mult_105_U542 ( .A1(DP_mult_105_n646), .A2(DP_mult_105_n249), 
        .B1(DP_mult_105_n646), .B2(DP_mult_105_n252), .C1(DP_mult_105_n252), 
        .C2(DP_mult_105_n249), .ZN(DP_mult_105_n645) );
  INV_X1 DP_mult_105_U541 ( .A(DP_mult_105_n645), .ZN(DP_mult_105_n644) );
  AOI222_X1 DP_mult_105_U540 ( .A1(DP_mult_105_n644), .A2(DP_mult_105_n245), 
        .B1(DP_mult_105_n644), .B2(DP_mult_105_n248), .C1(DP_mult_105_n248), 
        .C2(DP_mult_105_n245), .ZN(DP_mult_105_n643) );
  INV_X1 DP_mult_105_U539 ( .A(DP_mult_105_n643), .ZN(DP_mult_105_n642) );
  AOI222_X1 DP_mult_105_U538 ( .A1(DP_mult_105_n642), .A2(DP_mult_105_n239), 
        .B1(DP_mult_105_n642), .B2(DP_mult_105_n244), .C1(DP_mult_105_n244), 
        .C2(DP_mult_105_n239), .ZN(DP_mult_105_n639) );
  INV_X1 DP_mult_105_U537 ( .A(DP_mult_105_n233), .ZN(DP_mult_105_n640) );
  INV_X1 DP_mult_105_U536 ( .A(DP_mult_105_n238), .ZN(DP_mult_105_n641) );
  OAI222_X1 DP_mult_105_U535 ( .A1(DP_mult_105_n639), .A2(DP_mult_105_n640), 
        .B1(DP_mult_105_n639), .B2(DP_mult_105_n641), .C1(DP_mult_105_n641), 
        .C2(DP_mult_105_n640), .ZN(DP_mult_105_n638) );
  AOI222_X1 DP_mult_105_U534 ( .A1(DP_mult_105_n638), .A2(DP_mult_105_n225), 
        .B1(DP_mult_105_n638), .B2(DP_mult_105_n232), .C1(DP_mult_105_n232), 
        .C2(DP_mult_105_n225), .ZN(DP_mult_105_n635) );
  INV_X1 DP_mult_105_U533 ( .A(DP_mult_105_n217), .ZN(DP_mult_105_n636) );
  INV_X1 DP_mult_105_U532 ( .A(DP_mult_105_n224), .ZN(DP_mult_105_n637) );
  OAI222_X1 DP_mult_105_U531 ( .A1(DP_mult_105_n635), .A2(DP_mult_105_n636), 
        .B1(DP_mult_105_n635), .B2(DP_mult_105_n637), .C1(DP_mult_105_n637), 
        .C2(DP_mult_105_n636), .ZN(DP_mult_105_n126) );
  XNOR2_X1 DP_mult_105_U530 ( .A(DP_w_11_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n606) );
  INV_X1 DP_mult_105_U529 ( .A(DP_b_int[4]), .ZN(DP_mult_105_n622) );
  INV_X1 DP_mult_105_U528 ( .A(DP_b_int[2]), .ZN(DP_mult_105_n624) );
  XNOR2_X1 DP_mult_105_U527 ( .A(DP_mult_105_n624), .B(DP_b_int[3]), .ZN(
        DP_mult_105_n634) );
  NAND2_X1 DP_mult_105_U526 ( .A1(DP_mult_105_n593), .A2(DP_mult_105_n634), 
        .ZN(DP_mult_105_n595) );
  XNOR2_X1 DP_mult_105_U525 ( .A(DP_w_12_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n608) );
  OAI22_X1 DP_mult_105_U524 ( .A1(DP_mult_105_n606), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n608), .ZN(DP_mult_105_n142) );
  INV_X1 DP_mult_105_U523 ( .A(DP_mult_105_n142), .ZN(DP_mult_105_n143) );
  XNOR2_X1 DP_mult_105_U522 ( .A(DP_w_11_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n590) );
  INV_X1 DP_mult_105_U521 ( .A(DP_b_int[6]), .ZN(DP_mult_105_n620) );
  XNOR2_X1 DP_mult_105_U520 ( .A(DP_mult_105_n622), .B(DP_b_int[5]), .ZN(
        DP_mult_105_n633) );
  NAND2_X1 DP_mult_105_U519 ( .A1(DP_mult_105_n577), .A2(DP_mult_105_n633), 
        .ZN(DP_mult_105_n579) );
  XNOR2_X1 DP_mult_105_U518 ( .A(DP_w_12_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n592) );
  OAI22_X1 DP_mult_105_U517 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n592), .ZN(DP_mult_105_n152) );
  INV_X1 DP_mult_105_U516 ( .A(DP_mult_105_n152), .ZN(DP_mult_105_n153) );
  XNOR2_X1 DP_mult_105_U515 ( .A(DP_w_11_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n574) );
  XNOR2_X1 DP_mult_105_U514 ( .A(DP_mult_105_n620), .B(DP_b_int[7]), .ZN(
        DP_mult_105_n631) );
  NAND2_X1 DP_mult_105_U513 ( .A1(DP_mult_105_n561), .A2(DP_mult_105_n631), 
        .ZN(DP_mult_105_n563) );
  XNOR2_X1 DP_mult_105_U512 ( .A(DP_w_12_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n576) );
  OAI22_X1 DP_mult_105_U511 ( .A1(DP_mult_105_n574), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n576), .ZN(DP_mult_105_n166) );
  INV_X1 DP_mult_105_U510 ( .A(DP_mult_105_n166), .ZN(DP_mult_105_n167) );
  XNOR2_X1 DP_mult_105_U509 ( .A(DP_w_11_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n557) );
  XNOR2_X1 DP_mult_105_U508 ( .A(DP_w_12_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n559) );
  OAI22_X1 DP_mult_105_U507 ( .A1(DP_mult_105_n557), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n559), .ZN(DP_mult_105_n184) );
  INV_X1 DP_mult_105_U506 ( .A(DP_mult_105_n184), .ZN(DP_mult_105_n185) );
  XNOR2_X1 DP_mult_105_U505 ( .A(DP_w_4_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n599) );
  XNOR2_X1 DP_mult_105_U504 ( .A(DP_w_5_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n600) );
  OAI22_X1 DP_mult_105_U503 ( .A1(DP_mult_105_n599), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n600), .ZN(DP_mult_105_n629) );
  XNOR2_X1 DP_mult_105_U502 ( .A(DP_w_8_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n571) );
  XNOR2_X1 DP_mult_105_U501 ( .A(DP_w_9_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n572) );
  OAI22_X1 DP_mult_105_U500 ( .A1(DP_mult_105_n571), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n572), .ZN(DP_mult_105_n630) );
  OR2_X1 DP_mult_105_U499 ( .A1(DP_mult_105_n629), .A2(DP_mult_105_n630), .ZN(
        DP_mult_105_n194) );
  XNOR2_X1 DP_mult_105_U498 ( .A(DP_mult_105_n629), .B(DP_mult_105_n630), .ZN(
        DP_mult_105_n195) );
  INV_X1 DP_mult_105_U497 ( .A(DP_b_int[0]), .ZN(DP_mult_105_n626) );
  XNOR2_X1 DP_mult_105_U496 ( .A(DP_mult_105_n626), .B(DP_b_int[1]), .ZN(
        DP_mult_105_n628) );
  NAND2_X1 DP_mult_105_U495 ( .A1(DP_mult_105_n526), .A2(DP_mult_105_n628), 
        .ZN(DP_mult_105_n525) );
  OR3_X1 DP_mult_105_U494 ( .A1(DP_mult_105_n526), .A2(DP_w_0_), .A3(
        DP_mult_105_n626), .ZN(DP_mult_105_n627) );
  OAI21_X1 DP_mult_105_U493 ( .B1(DP_mult_105_n626), .B2(DP_mult_105_n525), 
        .A(DP_mult_105_n627), .ZN(DP_mult_105_n256) );
  OR3_X1 DP_mult_105_U492 ( .A1(DP_mult_105_n593), .A2(DP_w_0_), .A3(
        DP_mult_105_n624), .ZN(DP_mult_105_n625) );
  OAI21_X1 DP_mult_105_U491 ( .B1(DP_mult_105_n624), .B2(DP_mult_105_n595), 
        .A(DP_mult_105_n625), .ZN(DP_mult_105_n257) );
  OR3_X1 DP_mult_105_U490 ( .A1(DP_mult_105_n577), .A2(DP_w_0_), .A3(
        DP_mult_105_n622), .ZN(DP_mult_105_n623) );
  OAI21_X1 DP_mult_105_U489 ( .B1(DP_mult_105_n622), .B2(DP_mult_105_n579), 
        .A(DP_mult_105_n623), .ZN(DP_mult_105_n258) );
  OR3_X1 DP_mult_105_U488 ( .A1(DP_mult_105_n561), .A2(DP_w_0_), .A3(
        DP_mult_105_n620), .ZN(DP_mult_105_n621) );
  OAI21_X1 DP_mult_105_U487 ( .B1(DP_mult_105_n620), .B2(DP_mult_105_n563), 
        .A(DP_mult_105_n621), .ZN(DP_mult_105_n259) );
  XNOR2_X1 DP_mult_105_U486 ( .A(DP_w_10_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n619) );
  XNOR2_X1 DP_mult_105_U485 ( .A(DP_w_11_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n528) );
  OAI22_X1 DP_mult_105_U484 ( .A1(DP_mult_105_n619), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n528), .ZN(DP_mult_105_n263) );
  XNOR2_X1 DP_mult_105_U483 ( .A(DP_w_9_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n618) );
  OAI22_X1 DP_mult_105_U482 ( .A1(DP_mult_105_n618), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n619), .ZN(DP_mult_105_n264) );
  XNOR2_X1 DP_mult_105_U481 ( .A(DP_w_8_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n617) );
  OAI22_X1 DP_mult_105_U480 ( .A1(DP_mult_105_n617), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n618), .ZN(DP_mult_105_n265) );
  XNOR2_X1 DP_mult_105_U479 ( .A(DP_w_7_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n616) );
  OAI22_X1 DP_mult_105_U478 ( .A1(DP_mult_105_n616), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n617), .ZN(DP_mult_105_n266) );
  XNOR2_X1 DP_mult_105_U477 ( .A(DP_w_6_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n615) );
  OAI22_X1 DP_mult_105_U476 ( .A1(DP_mult_105_n615), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n616), .ZN(DP_mult_105_n267) );
  XNOR2_X1 DP_mult_105_U475 ( .A(DP_w_5_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n614) );
  OAI22_X1 DP_mult_105_U474 ( .A1(DP_mult_105_n614), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n615), .ZN(DP_mult_105_n268) );
  XNOR2_X1 DP_mult_105_U473 ( .A(DP_w_4_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n613) );
  OAI22_X1 DP_mult_105_U472 ( .A1(DP_mult_105_n613), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n614), .ZN(DP_mult_105_n269) );
  XNOR2_X1 DP_mult_105_U471 ( .A(DP_w_3_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n612) );
  OAI22_X1 DP_mult_105_U470 ( .A1(DP_mult_105_n612), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n613), .ZN(DP_mult_105_n270) );
  XNOR2_X1 DP_mult_105_U469 ( .A(DP_w_2_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n611) );
  OAI22_X1 DP_mult_105_U468 ( .A1(DP_mult_105_n611), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n612), .ZN(DP_mult_105_n271) );
  XNOR2_X1 DP_mult_105_U467 ( .A(DP_w_1_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n610) );
  OAI22_X1 DP_mult_105_U466 ( .A1(DP_mult_105_n610), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n611), .ZN(DP_mult_105_n272) );
  XNOR2_X1 DP_mult_105_U465 ( .A(DP_w_0_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n609) );
  OAI22_X1 DP_mult_105_U464 ( .A1(DP_mult_105_n609), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n610), .ZN(DP_mult_105_n273) );
  NOR2_X1 DP_mult_105_U463 ( .A1(DP_mult_105_n560), .A2(DP_mult_105_n526), 
        .ZN(DP_mult_105_n274) );
  AOI21_X1 DP_mult_105_U462 ( .B1(DP_mult_105_n595), .B2(DP_mult_105_n593), 
        .A(DP_mult_105_n608), .ZN(DP_mult_105_n607) );
  INV_X1 DP_mult_105_U461 ( .A(DP_mult_105_n607), .ZN(DP_mult_105_n275) );
  XNOR2_X1 DP_mult_105_U460 ( .A(DP_w_10_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n605) );
  OAI22_X1 DP_mult_105_U459 ( .A1(DP_mult_105_n605), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n606), .ZN(DP_mult_105_n276) );
  XNOR2_X1 DP_mult_105_U458 ( .A(DP_w_9_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n604) );
  OAI22_X1 DP_mult_105_U457 ( .A1(DP_mult_105_n604), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n605), .ZN(DP_mult_105_n277) );
  XNOR2_X1 DP_mult_105_U456 ( .A(DP_w_8_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n603) );
  OAI22_X1 DP_mult_105_U455 ( .A1(DP_mult_105_n603), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n604), .ZN(DP_mult_105_n278) );
  XNOR2_X1 DP_mult_105_U454 ( .A(DP_w_7_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n602) );
  OAI22_X1 DP_mult_105_U453 ( .A1(DP_mult_105_n602), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n603), .ZN(DP_mult_105_n279) );
  XNOR2_X1 DP_mult_105_U452 ( .A(DP_w_6_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n601) );
  OAI22_X1 DP_mult_105_U451 ( .A1(DP_mult_105_n601), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n602), .ZN(DP_mult_105_n280) );
  OAI22_X1 DP_mult_105_U450 ( .A1(DP_mult_105_n600), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n601), .ZN(DP_mult_105_n281) );
  XNOR2_X1 DP_mult_105_U449 ( .A(DP_w_3_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n598) );
  OAI22_X1 DP_mult_105_U448 ( .A1(DP_mult_105_n598), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n599), .ZN(DP_mult_105_n283) );
  XNOR2_X1 DP_mult_105_U447 ( .A(DP_w_2_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n597) );
  OAI22_X1 DP_mult_105_U446 ( .A1(DP_mult_105_n597), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n598), .ZN(DP_mult_105_n284) );
  XNOR2_X1 DP_mult_105_U445 ( .A(DP_w_1_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n596) );
  OAI22_X1 DP_mult_105_U444 ( .A1(DP_mult_105_n596), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n597), .ZN(DP_mult_105_n285) );
  XNOR2_X1 DP_mult_105_U443 ( .A(DP_w_0_), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n594) );
  OAI22_X1 DP_mult_105_U442 ( .A1(DP_mult_105_n594), .A2(DP_mult_105_n595), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n286) );
  NOR2_X1 DP_mult_105_U441 ( .A1(DP_mult_105_n560), .A2(DP_mult_105_n593), 
        .ZN(DP_mult_105_n287) );
  AOI21_X1 DP_mult_105_U440 ( .B1(DP_mult_105_n579), .B2(DP_mult_105_n577), 
        .A(DP_mult_105_n592), .ZN(DP_mult_105_n591) );
  INV_X1 DP_mult_105_U439 ( .A(DP_mult_105_n591), .ZN(DP_mult_105_n288) );
  XNOR2_X1 DP_mult_105_U438 ( .A(DP_w_10_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n589) );
  OAI22_X1 DP_mult_105_U437 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n590), .ZN(DP_mult_105_n289) );
  XNOR2_X1 DP_mult_105_U436 ( .A(DP_w_9_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n588) );
  OAI22_X1 DP_mult_105_U435 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n589), .ZN(DP_mult_105_n290) );
  XNOR2_X1 DP_mult_105_U434 ( .A(DP_w_8_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n587) );
  OAI22_X1 DP_mult_105_U433 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n588), .ZN(DP_mult_105_n291) );
  XNOR2_X1 DP_mult_105_U432 ( .A(DP_w_7_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n586) );
  OAI22_X1 DP_mult_105_U431 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n587), .ZN(DP_mult_105_n292) );
  XNOR2_X1 DP_mult_105_U430 ( .A(DP_w_6_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n585) );
  OAI22_X1 DP_mult_105_U429 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n586), .ZN(DP_mult_105_n293) );
  XNOR2_X1 DP_mult_105_U428 ( .A(DP_w_5_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n584) );
  OAI22_X1 DP_mult_105_U427 ( .A1(DP_mult_105_n584), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n585), .ZN(DP_mult_105_n294) );
  XNOR2_X1 DP_mult_105_U426 ( .A(DP_w_4_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n583) );
  OAI22_X1 DP_mult_105_U425 ( .A1(DP_mult_105_n583), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n584), .ZN(DP_mult_105_n295) );
  XNOR2_X1 DP_mult_105_U424 ( .A(DP_w_3_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n582) );
  OAI22_X1 DP_mult_105_U423 ( .A1(DP_mult_105_n582), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n583), .ZN(DP_mult_105_n296) );
  XNOR2_X1 DP_mult_105_U422 ( .A(DP_w_2_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n581) );
  OAI22_X1 DP_mult_105_U421 ( .A1(DP_mult_105_n581), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n582), .ZN(DP_mult_105_n297) );
  XNOR2_X1 DP_mult_105_U420 ( .A(DP_w_1_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n580) );
  OAI22_X1 DP_mult_105_U419 ( .A1(DP_mult_105_n580), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n581), .ZN(DP_mult_105_n298) );
  XNOR2_X1 DP_mult_105_U418 ( .A(DP_w_0_), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n578) );
  OAI22_X1 DP_mult_105_U417 ( .A1(DP_mult_105_n578), .A2(DP_mult_105_n579), 
        .B1(DP_mult_105_n577), .B2(DP_mult_105_n580), .ZN(DP_mult_105_n299) );
  NOR2_X1 DP_mult_105_U416 ( .A1(DP_mult_105_n560), .A2(DP_mult_105_n577), 
        .ZN(DP_mult_105_n300) );
  AOI21_X1 DP_mult_105_U415 ( .B1(DP_mult_105_n563), .B2(DP_mult_105_n561), 
        .A(DP_mult_105_n576), .ZN(DP_mult_105_n575) );
  INV_X1 DP_mult_105_U414 ( .A(DP_mult_105_n575), .ZN(DP_mult_105_n301) );
  XNOR2_X1 DP_mult_105_U413 ( .A(DP_w_10_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n573) );
  OAI22_X1 DP_mult_105_U412 ( .A1(DP_mult_105_n573), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n574), .ZN(DP_mult_105_n302) );
  OAI22_X1 DP_mult_105_U411 ( .A1(DP_mult_105_n572), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n573), .ZN(DP_mult_105_n303) );
  XNOR2_X1 DP_mult_105_U410 ( .A(DP_w_7_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n570) );
  OAI22_X1 DP_mult_105_U409 ( .A1(DP_mult_105_n570), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n571), .ZN(DP_mult_105_n305) );
  XNOR2_X1 DP_mult_105_U408 ( .A(DP_w_6_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n569) );
  OAI22_X1 DP_mult_105_U407 ( .A1(DP_mult_105_n569), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n570), .ZN(DP_mult_105_n306) );
  XNOR2_X1 DP_mult_105_U406 ( .A(DP_w_5_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n568) );
  OAI22_X1 DP_mult_105_U405 ( .A1(DP_mult_105_n568), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n569), .ZN(DP_mult_105_n307) );
  XNOR2_X1 DP_mult_105_U404 ( .A(DP_w_4_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n567) );
  OAI22_X1 DP_mult_105_U403 ( .A1(DP_mult_105_n567), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n568), .ZN(DP_mult_105_n308) );
  XNOR2_X1 DP_mult_105_U402 ( .A(DP_w_3_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n566) );
  OAI22_X1 DP_mult_105_U401 ( .A1(DP_mult_105_n566), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n567), .ZN(DP_mult_105_n309) );
  XNOR2_X1 DP_mult_105_U400 ( .A(DP_w_2_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n565) );
  OAI22_X1 DP_mult_105_U399 ( .A1(DP_mult_105_n565), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n566), .ZN(DP_mult_105_n310) );
  XNOR2_X1 DP_mult_105_U398 ( .A(DP_w_1_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n564) );
  OAI22_X1 DP_mult_105_U397 ( .A1(DP_mult_105_n564), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n565), .ZN(DP_mult_105_n311) );
  XNOR2_X1 DP_mult_105_U396 ( .A(DP_w_0_), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n562) );
  OAI22_X1 DP_mult_105_U395 ( .A1(DP_mult_105_n562), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n564), .ZN(DP_mult_105_n312) );
  NOR2_X1 DP_mult_105_U394 ( .A1(DP_mult_105_n560), .A2(DP_mult_105_n561), 
        .ZN(DP_mult_105_n313) );
  AOI21_X1 DP_mult_105_U393 ( .B1(DP_mult_105_n545), .B2(DP_mult_105_n546), 
        .A(DP_mult_105_n559), .ZN(DP_mult_105_n558) );
  INV_X1 DP_mult_105_U392 ( .A(DP_mult_105_n558), .ZN(DP_mult_105_n314) );
  XNOR2_X1 DP_mult_105_U391 ( .A(DP_w_10_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n556) );
  OAI22_X1 DP_mult_105_U390 ( .A1(DP_mult_105_n556), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n557), .ZN(DP_mult_105_n315) );
  XNOR2_X1 DP_mult_105_U389 ( .A(DP_w_9_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n555) );
  OAI22_X1 DP_mult_105_U388 ( .A1(DP_mult_105_n555), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n556), .ZN(DP_mult_105_n316) );
  XNOR2_X1 DP_mult_105_U387 ( .A(DP_w_8_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n554) );
  OAI22_X1 DP_mult_105_U386 ( .A1(DP_mult_105_n554), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n555), .ZN(DP_mult_105_n317) );
  XNOR2_X1 DP_mult_105_U385 ( .A(DP_w_7_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n553) );
  OAI22_X1 DP_mult_105_U384 ( .A1(DP_mult_105_n553), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n554), .ZN(DP_mult_105_n318) );
  XNOR2_X1 DP_mult_105_U383 ( .A(DP_w_6_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n552) );
  OAI22_X1 DP_mult_105_U382 ( .A1(DP_mult_105_n552), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n553), .ZN(DP_mult_105_n319) );
  XNOR2_X1 DP_mult_105_U381 ( .A(DP_w_5_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n551) );
  OAI22_X1 DP_mult_105_U380 ( .A1(DP_mult_105_n551), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n552), .ZN(DP_mult_105_n320) );
  XNOR2_X1 DP_mult_105_U379 ( .A(DP_w_4_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n550) );
  OAI22_X1 DP_mult_105_U378 ( .A1(DP_mult_105_n550), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n551), .ZN(DP_mult_105_n321) );
  XNOR2_X1 DP_mult_105_U377 ( .A(DP_w_3_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n549) );
  OAI22_X1 DP_mult_105_U376 ( .A1(DP_mult_105_n549), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n550), .ZN(DP_mult_105_n322) );
  XNOR2_X1 DP_mult_105_U375 ( .A(DP_w_2_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n548) );
  OAI22_X1 DP_mult_105_U374 ( .A1(DP_mult_105_n548), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n549), .ZN(DP_mult_105_n323) );
  XNOR2_X1 DP_mult_105_U373 ( .A(DP_w_1_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n547) );
  OAI22_X1 DP_mult_105_U372 ( .A1(DP_mult_105_n547), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n548), .ZN(DP_mult_105_n324) );
  XNOR2_X1 DP_mult_105_U371 ( .A(DP_w_0_), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n544) );
  OAI22_X1 DP_mult_105_U370 ( .A1(DP_mult_105_n544), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n546), .B2(DP_mult_105_n547), .ZN(DP_mult_105_n325) );
  XOR2_X1 DP_mult_105_U369 ( .A(DP_w_12_), .B(DP_mult_105_n543), .Z(
        DP_mult_105_n541) );
  AOI21_X1 DP_mult_105_U368 ( .B1(DP_mult_105_n530), .B2(DP_mult_105_n532), 
        .A(DP_mult_105_n541), .ZN(DP_mult_105_n542) );
  INV_X1 DP_mult_105_U367 ( .A(DP_mult_105_n542), .ZN(DP_mult_105_n327) );
  XNOR2_X1 DP_mult_105_U366 ( .A(DP_w_11_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n540) );
  OAI22_X1 DP_mult_105_U365 ( .A1(DP_mult_105_n540), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n541), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n328) );
  XNOR2_X1 DP_mult_105_U364 ( .A(DP_w_10_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n539) );
  OAI22_X1 DP_mult_105_U363 ( .A1(DP_mult_105_n539), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n540), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n329) );
  XNOR2_X1 DP_mult_105_U362 ( .A(DP_w_9_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n538) );
  OAI22_X1 DP_mult_105_U361 ( .A1(DP_mult_105_n538), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n539), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n330) );
  XNOR2_X1 DP_mult_105_U360 ( .A(DP_w_8_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n537) );
  OAI22_X1 DP_mult_105_U359 ( .A1(DP_mult_105_n537), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n538), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n331) );
  XNOR2_X1 DP_mult_105_U358 ( .A(DP_w_7_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n536) );
  OAI22_X1 DP_mult_105_U357 ( .A1(DP_mult_105_n536), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n537), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n332) );
  XNOR2_X1 DP_mult_105_U356 ( .A(DP_w_6_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n535) );
  OAI22_X1 DP_mult_105_U355 ( .A1(DP_mult_105_n535), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n536), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n333) );
  XNOR2_X1 DP_mult_105_U354 ( .A(DP_w_5_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n534) );
  OAI22_X1 DP_mult_105_U353 ( .A1(DP_mult_105_n534), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n535), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n334) );
  XNOR2_X1 DP_mult_105_U352 ( .A(DP_w_4_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n533) );
  OAI22_X1 DP_mult_105_U351 ( .A1(DP_mult_105_n533), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n534), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n335) );
  XNOR2_X1 DP_mult_105_U350 ( .A(DP_w_3_), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n531) );
  OAI22_X1 DP_mult_105_U349 ( .A1(DP_mult_105_n531), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n533), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n336) );
  OAI22_X1 DP_mult_105_U348 ( .A1(DP_mult_105_n529), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n531), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n337) );
  XNOR2_X1 DP_mult_105_U347 ( .A(DP_w_12_), .B(DP_b_int[0]), .ZN(
        DP_mult_105_n527) );
  OAI22_X1 DP_mult_105_U346 ( .A1(DP_mult_105_n528), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n526), .B2(DP_mult_105_n527), .ZN(DP_mult_105_n519) );
  AOI21_X1 DP_mult_105_U345 ( .B1(DP_mult_105_n525), .B2(DP_mult_105_n526), 
        .A(DP_mult_105_n527), .ZN(DP_mult_105_n522) );
  INV_X1 DP_mult_105_U344 ( .A(DP_mult_105_n522), .ZN(DP_mult_105_n520) );
  INV_X1 DP_mult_105_U343 ( .A(DP_mult_105_n519), .ZN(DP_mult_105_n524) );
  AOI222_X1 DP_mult_105_U342 ( .A1(DP_mult_105_n115), .A2(DP_mult_105_n138), 
        .B1(DP_mult_105_n524), .B2(DP_mult_105_n115), .C1(DP_mult_105_n524), 
        .C2(DP_mult_105_n138), .ZN(DP_mult_105_n523) );
  OAI22_X1 DP_mult_105_U341 ( .A1(DP_mult_105_n522), .A2(DP_mult_105_n523), 
        .B1(DP_mult_105_n524), .B2(DP_mult_105_n523), .ZN(DP_mult_105_n521) );
  AOI21_X1 DP_mult_105_U340 ( .B1(DP_mult_105_n519), .B2(DP_mult_105_n520), 
        .A(DP_mult_105_n521), .ZN(DP_w_b0_11_) );
  XOR2_X2 DP_mult_105_U339 ( .A(DP_b_int[3]), .B(DP_mult_105_n622), .Z(
        DP_mult_105_n593) );
  XOR2_X2 DP_mult_105_U338 ( .A(DP_b_int[5]), .B(DP_mult_105_n620), .Z(
        DP_mult_105_n577) );
  XOR2_X2 DP_mult_105_U337 ( .A(DP_b_int[7]), .B(DP_mult_105_n632), .Z(
        DP_mult_105_n561) );
  XOR2_X2 DP_mult_105_U336 ( .A(DP_b_int[1]), .B(DP_mult_105_n624), .Z(
        DP_mult_105_n526) );
  INV_X1 DP_mult_105_U335 ( .A(DP_b_int[11]), .ZN(DP_mult_105_n532) );
  INV_X1 DP_mult_105_U334 ( .A(DP_mult_105_n653), .ZN(DP_mult_105_n546) );
  HA_X1 DP_mult_105_U120 ( .A(DP_mult_105_n325), .B(DP_mult_105_n337), .CO(
        DP_mult_105_n254), .S(DP_mult_105_n255) );
  FA_X1 DP_mult_105_U119 ( .A(DP_mult_105_n336), .B(DP_mult_105_n313), .CI(
        DP_mult_105_n324), .CO(DP_mult_105_n252), .S(DP_mult_105_n253) );
  HA_X1 DP_mult_105_U118 ( .A(DP_mult_105_n259), .B(DP_mult_105_n312), .CO(
        DP_mult_105_n250), .S(DP_mult_105_n251) );
  FA_X1 DP_mult_105_U117 ( .A(DP_mult_105_n323), .B(DP_mult_105_n335), .CI(
        DP_mult_105_n251), .CO(DP_mult_105_n248), .S(DP_mult_105_n249) );
  FA_X1 DP_mult_105_U109 ( .A(DP_mult_105_n334), .B(DP_mult_105_n300), .CI(
        DP_mult_105_n322), .CO(DP_mult_105_n246), .S(DP_mult_105_n247) );
  FA_X1 DP_mult_105_U108 ( .A(DP_mult_105_n250), .B(DP_mult_105_n311), .CI(
        DP_mult_105_n247), .CO(DP_mult_105_n244), .S(DP_mult_105_n245) );
  HA_X1 DP_mult_105_U107 ( .A(DP_mult_105_n258), .B(DP_mult_105_n299), .CO(
        DP_mult_105_n242), .S(DP_mult_105_n243) );
  FA_X1 DP_mult_105_U106 ( .A(DP_mult_105_n310), .B(DP_mult_105_n333), .CI(
        DP_mult_105_n321), .CO(DP_mult_105_n240), .S(DP_mult_105_n241) );
  FA_X1 DP_mult_105_U105 ( .A(DP_mult_105_n246), .B(DP_mult_105_n243), .CI(
        DP_mult_105_n241), .CO(DP_mult_105_n238), .S(DP_mult_105_n239) );
  FA_X1 DP_mult_105_U104 ( .A(DP_mult_105_n309), .B(DP_mult_105_n287), .CI(
        DP_mult_105_n332), .CO(DP_mult_105_n236), .S(DP_mult_105_n237) );
  FA_X1 DP_mult_105_U103 ( .A(DP_mult_105_n298), .B(DP_mult_105_n320), .CI(
        DP_mult_105_n242), .CO(DP_mult_105_n234), .S(DP_mult_105_n235) );
  FA_X1 DP_mult_105_U102 ( .A(DP_mult_105_n237), .B(DP_mult_105_n240), .CI(
        DP_mult_105_n235), .CO(DP_mult_105_n232), .S(DP_mult_105_n233) );
  HA_X1 DP_mult_105_U101 ( .A(DP_mult_105_n257), .B(DP_mult_105_n286), .CO(
        DP_mult_105_n230), .S(DP_mult_105_n231) );
  FA_X1 DP_mult_105_U100 ( .A(DP_mult_105_n297), .B(DP_mult_105_n308), .CI(
        DP_mult_105_n319), .CO(DP_mult_105_n228), .S(DP_mult_105_n229) );
  FA_X1 DP_mult_105_U99 ( .A(DP_mult_105_n231), .B(DP_mult_105_n331), .CI(
        DP_mult_105_n236), .CO(DP_mult_105_n226), .S(DP_mult_105_n227) );
  FA_X1 DP_mult_105_U98 ( .A(DP_mult_105_n229), .B(DP_mult_105_n234), .CI(
        DP_mult_105_n227), .CO(DP_mult_105_n224), .S(DP_mult_105_n225) );
  FA_X1 DP_mult_105_U97 ( .A(DP_mult_105_n296), .B(DP_mult_105_n274), .CI(
        DP_mult_105_n330), .CO(DP_mult_105_n222), .S(DP_mult_105_n223) );
  FA_X1 DP_mult_105_U96 ( .A(DP_mult_105_n285), .B(DP_mult_105_n318), .CI(
        DP_mult_105_n307), .CO(DP_mult_105_n220), .S(DP_mult_105_n221) );
  FA_X1 DP_mult_105_U95 ( .A(DP_mult_105_n228), .B(DP_mult_105_n230), .CI(
        DP_mult_105_n223), .CO(DP_mult_105_n218), .S(DP_mult_105_n219) );
  FA_X1 DP_mult_105_U94 ( .A(DP_mult_105_n226), .B(DP_mult_105_n221), .CI(
        DP_mult_105_n219), .CO(DP_mult_105_n216), .S(DP_mult_105_n217) );
  HA_X1 DP_mult_105_U93 ( .A(DP_mult_105_n256), .B(DP_mult_105_n273), .CO(
        DP_mult_105_n214), .S(DP_mult_105_n215) );
  FA_X1 DP_mult_105_U92 ( .A(DP_mult_105_n284), .B(DP_mult_105_n306), .CI(
        DP_mult_105_n329), .CO(DP_mult_105_n212), .S(DP_mult_105_n213) );
  FA_X1 DP_mult_105_U91 ( .A(DP_mult_105_n295), .B(DP_mult_105_n317), .CI(
        DP_mult_105_n215), .CO(DP_mult_105_n210), .S(DP_mult_105_n211) );
  FA_X1 DP_mult_105_U90 ( .A(DP_mult_105_n220), .B(DP_mult_105_n222), .CI(
        DP_mult_105_n213), .CO(DP_mult_105_n208), .S(DP_mult_105_n209) );
  FA_X1 DP_mult_105_U89 ( .A(DP_mult_105_n218), .B(DP_mult_105_n211), .CI(
        DP_mult_105_n209), .CO(DP_mult_105_n206), .S(DP_mult_105_n207) );
  HA_X1 DP_mult_105_U88 ( .A(DP_mult_105_n272), .B(DP_mult_105_n283), .CO(
        DP_mult_105_n204), .S(DP_mult_105_n205) );
  FA_X1 DP_mult_105_U87 ( .A(DP_mult_105_n328), .B(DP_mult_105_n305), .CI(
        DP_mult_105_n294), .CO(DP_mult_105_n202), .S(DP_mult_105_n203) );
  FA_X1 DP_mult_105_U86 ( .A(DP_mult_105_n214), .B(DP_mult_105_n316), .CI(
        DP_mult_105_n205), .CO(DP_mult_105_n200), .S(DP_mult_105_n201) );
  FA_X1 DP_mult_105_U85 ( .A(DP_mult_105_n203), .B(DP_mult_105_n212), .CI(
        DP_mult_105_n210), .CO(DP_mult_105_n198), .S(DP_mult_105_n199) );
  FA_X1 DP_mult_105_U84 ( .A(DP_mult_105_n208), .B(DP_mult_105_n201), .CI(
        DP_mult_105_n199), .CO(DP_mult_105_n196), .S(DP_mult_105_n197) );
  FA_X1 DP_mult_105_U81 ( .A(DP_mult_105_n271), .B(DP_mult_105_n293), .CI(
        DP_mult_105_n327), .CO(DP_mult_105_n192), .S(DP_mult_105_n193) );
  FA_X1 DP_mult_105_U80 ( .A(DP_mult_105_n204), .B(DP_mult_105_n315), .CI(
        DP_mult_105_n195), .CO(DP_mult_105_n190), .S(DP_mult_105_n191) );
  FA_X1 DP_mult_105_U79 ( .A(DP_mult_105_n193), .B(DP_mult_105_n202), .CI(
        DP_mult_105_n200), .CO(DP_mult_105_n188), .S(DP_mult_105_n189) );
  FA_X1 DP_mult_105_U78 ( .A(DP_mult_105_n198), .B(DP_mult_105_n191), .CI(
        DP_mult_105_n189), .CO(DP_mult_105_n186), .S(DP_mult_105_n187) );
  FA_X1 DP_mult_105_U76 ( .A(DP_mult_105_n303), .B(DP_mult_105_n281), .CI(
        DP_mult_105_n185), .CO(DP_mult_105_n182), .S(DP_mult_105_n183) );
  FA_X1 DP_mult_105_U75 ( .A(DP_mult_105_n270), .B(DP_mult_105_n292), .CI(
        DP_mult_105_n194), .CO(DP_mult_105_n180), .S(DP_mult_105_n181) );
  FA_X1 DP_mult_105_U74 ( .A(DP_mult_105_n190), .B(DP_mult_105_n192), .CI(
        DP_mult_105_n183), .CO(DP_mult_105_n178), .S(DP_mult_105_n179) );
  FA_X1 DP_mult_105_U73 ( .A(DP_mult_105_n188), .B(DP_mult_105_n181), .CI(
        DP_mult_105_n179), .CO(DP_mult_105_n176), .S(DP_mult_105_n177) );
  FA_X1 DP_mult_105_U72 ( .A(DP_mult_105_n184), .B(DP_mult_105_n269), .CI(
        DP_mult_105_n314), .CO(DP_mult_105_n174), .S(DP_mult_105_n175) );
  FA_X1 DP_mult_105_U71 ( .A(DP_mult_105_n280), .B(DP_mult_105_n302), .CI(
        DP_mult_105_n291), .CO(DP_mult_105_n172), .S(DP_mult_105_n173) );
  FA_X1 DP_mult_105_U70 ( .A(DP_mult_105_n180), .B(DP_mult_105_n182), .CI(
        DP_mult_105_n173), .CO(DP_mult_105_n170), .S(DP_mult_105_n171) );
  FA_X1 DP_mult_105_U69 ( .A(DP_mult_105_n178), .B(DP_mult_105_n175), .CI(
        DP_mult_105_n171), .CO(DP_mult_105_n168), .S(DP_mult_105_n169) );
  FA_X1 DP_mult_105_U67 ( .A(DP_mult_105_n268), .B(DP_mult_105_n279), .CI(
        DP_mult_105_n167), .CO(DP_mult_105_n164), .S(DP_mult_105_n165) );
  FA_X1 DP_mult_105_U66 ( .A(DP_mult_105_n174), .B(DP_mult_105_n290), .CI(
        DP_mult_105_n172), .CO(DP_mult_105_n162), .S(DP_mult_105_n163) );
  FA_X1 DP_mult_105_U65 ( .A(DP_mult_105_n170), .B(DP_mult_105_n165), .CI(
        DP_mult_105_n163), .CO(DP_mult_105_n160), .S(DP_mult_105_n161) );
  FA_X1 DP_mult_105_U64 ( .A(DP_mult_105_n166), .B(DP_mult_105_n267), .CI(
        DP_mult_105_n301), .CO(DP_mult_105_n158), .S(DP_mult_105_n159) );
  FA_X1 DP_mult_105_U63 ( .A(DP_mult_105_n278), .B(DP_mult_105_n289), .CI(
        DP_mult_105_n164), .CO(DP_mult_105_n156), .S(DP_mult_105_n157) );
  FA_X1 DP_mult_105_U62 ( .A(DP_mult_105_n162), .B(DP_mult_105_n159), .CI(
        DP_mult_105_n157), .CO(DP_mult_105_n154), .S(DP_mult_105_n155) );
  FA_X1 DP_mult_105_U60 ( .A(DP_mult_105_n266), .B(DP_mult_105_n277), .CI(
        DP_mult_105_n153), .CO(DP_mult_105_n150), .S(DP_mult_105_n151) );
  FA_X1 DP_mult_105_U59 ( .A(DP_mult_105_n151), .B(DP_mult_105_n158), .CI(
        DP_mult_105_n156), .CO(DP_mult_105_n148), .S(DP_mult_105_n149) );
  FA_X1 DP_mult_105_U58 ( .A(DP_mult_105_n265), .B(DP_mult_105_n152), .CI(
        DP_mult_105_n288), .CO(DP_mult_105_n146), .S(DP_mult_105_n147) );
  FA_X1 DP_mult_105_U57 ( .A(DP_mult_105_n150), .B(DP_mult_105_n276), .CI(
        DP_mult_105_n147), .CO(DP_mult_105_n144), .S(DP_mult_105_n145) );
  FA_X1 DP_mult_105_U55 ( .A(DP_mult_105_n143), .B(DP_mult_105_n264), .CI(
        DP_mult_105_n146), .CO(DP_mult_105_n140), .S(DP_mult_105_n141) );
  FA_X1 DP_mult_105_U54 ( .A(DP_mult_105_n263), .B(DP_mult_105_n142), .CI(
        DP_mult_105_n275), .CO(DP_mult_105_n138), .S(DP_mult_105_n139) );
  FA_X1 DP_mult_105_U42 ( .A(DP_mult_105_n207), .B(DP_mult_105_n216), .CI(
        DP_mult_105_n126), .CO(DP_mult_105_n125), .S(DP_w_b0_0_) );
  FA_X1 DP_mult_105_U41 ( .A(DP_mult_105_n197), .B(DP_mult_105_n206), .CI(
        DP_mult_105_n125), .CO(DP_mult_105_n124), .S(DP_w_b0_1_) );
  FA_X1 DP_mult_105_U40 ( .A(DP_mult_105_n187), .B(DP_mult_105_n196), .CI(
        DP_mult_105_n124), .CO(DP_mult_105_n123), .S(DP_w_b0_2_) );
  FA_X1 DP_mult_105_U39 ( .A(DP_mult_105_n177), .B(DP_mult_105_n186), .CI(
        DP_mult_105_n123), .CO(DP_mult_105_n122), .S(DP_w_b0_3_) );
  FA_X1 DP_mult_105_U38 ( .A(DP_mult_105_n169), .B(DP_mult_105_n176), .CI(
        DP_mult_105_n122), .CO(DP_mult_105_n121), .S(DP_w_b0_4_) );
  FA_X1 DP_mult_105_U37 ( .A(DP_mult_105_n161), .B(DP_mult_105_n168), .CI(
        DP_mult_105_n121), .CO(DP_mult_105_n120), .S(DP_w_b0_5_) );
  FA_X1 DP_mult_105_U36 ( .A(DP_mult_105_n155), .B(DP_mult_105_n160), .CI(
        DP_mult_105_n120), .CO(DP_mult_105_n119), .S(DP_w_b0_6_) );
  FA_X1 DP_mult_105_U30 ( .A(DP_mult_105_n149), .B(DP_mult_105_n154), .CI(
        DP_mult_105_n119), .CO(DP_mult_105_n118), .S(DP_w_b0_7_) );
  FA_X1 DP_mult_105_U20 ( .A(DP_mult_105_n145), .B(DP_mult_105_n148), .CI(
        DP_mult_105_n118), .CO(DP_mult_105_n117), .S(DP_w_b0_8_) );
  FA_X1 DP_mult_105_U10 ( .A(DP_mult_105_n141), .B(DP_mult_105_n144), .CI(
        DP_mult_105_n117), .CO(DP_mult_105_n116), .S(DP_w_b0_9_) );
  FA_X1 DP_mult_105_U9 ( .A(DP_mult_105_n140), .B(DP_mult_105_n139), .CI(
        DP_mult_105_n116), .CO(DP_mult_105_n115), .S(DP_w_b0_10_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U14 ( .A(DP_sw1_a2_0_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_0_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U13 ( .A(DP_sw1_a2_10_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_10_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U12 ( .A(DP_sw1_a2_11_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_12_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U11 ( .A(DP_sw1_a2_1_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_1_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U10 ( .A(DP_sw1_a2_2_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_2_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U9 ( .A(DP_sw1_a2_3_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_3_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U8 ( .A(DP_sw1_a2_4_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_4_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U7 ( .A(DP_sw1_a2_5_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_5_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U6 ( .A(DP_sw1_a2_6_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_6_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U5 ( .A(DP_sw1_a2_7_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_7_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U4 ( .A(DP_sw1_a2_8_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_8_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U3 ( .A(DP_sw1_a2_9_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_B_not_9_) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U2 ( .A(DP_x_0_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_0_), .ZN(DP_fb_0_) );
  OR2_X1 DP_sub_1_root_sub_0_root_sub_104_U1 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_B_not_0_), .A2(DP_x_0_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_carry_1_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_1 ( .A(DP_x_1_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_1_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_1_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_2_), .S(DP_fb_1_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_2 ( .A(DP_x_2_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_2_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_2_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_3_), .S(DP_fb_2_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_3 ( .A(DP_x_3_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_3_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_3_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_4_), .S(DP_fb_3_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_4 ( .A(DP_x_4_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_4_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_4_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_5_), .S(DP_fb_4_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_5 ( .A(DP_x_5_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_5_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_5_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_6_), .S(DP_fb_5_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_6 ( .A(DP_x_6_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_6_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_6_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_7_), .S(DP_fb_6_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_7 ( .A(DP_x_7_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_7_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_7_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_8_), .S(DP_fb_7_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_8 ( .A(DP_x_8_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_8_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_8_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_9_), .S(DP_fb_8_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_9 ( .A(DP_x_9_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_9_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_9_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_10_), .S(DP_fb_9_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_10 ( .A(DP_x_10_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_10_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_10_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_11_), .S(DP_fb_10_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_11 ( .A(DP_x_11_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_12_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_11_), .CO(
        DP_sub_1_root_sub_0_root_sub_104_carry_12_), .S(DP_fb_11_) );
  FA_X1 DP_sub_1_root_sub_0_root_sub_104_U2_12 ( .A(DP_x_11_), .B(
        DP_sub_1_root_sub_0_root_sub_104_B_not_12_), .CI(
        DP_sub_1_root_sub_0_root_sub_104_carry_12_), .S(DP_fb_12_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U14 ( .A(DP_sw0_a1_0_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_0_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U13 ( .A(DP_sw0_a1_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_10_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U12 ( .A(DP_sw0_a1_11_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_12_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U11 ( .A(DP_sw0_a1_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_1_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U10 ( .A(DP_sw0_a1_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_2_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U9 ( .A(DP_sw0_a1_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_3_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U8 ( .A(DP_sw0_a1_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_4_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U7 ( .A(DP_sw0_a1_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_5_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U6 ( .A(DP_sw0_a1_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_6_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U5 ( .A(DP_sw0_a1_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_7_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U4 ( .A(DP_sw0_a1_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_8_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U3 ( .A(DP_sw0_a1_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_9_) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U2 ( .A(DP_fb_0_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_0_), .ZN(DP_w_0_) );
  OR2_X1 DP_sub_0_root_sub_0_root_sub_104_U1 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_B_not_0_), .A2(DP_fb_0_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_1_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_1 ( .A(DP_fb_1_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_1_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_1_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_2_), .S(DP_w_1_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_2 ( .A(DP_fb_2_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_2_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_2_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_3_), .S(DP_w_2_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_3 ( .A(DP_fb_3_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_3_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_3_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_4_), .S(DP_w_3_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_4 ( .A(DP_fb_4_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_4_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_4_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_5_), .S(DP_w_4_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_5 ( .A(DP_fb_5_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_5_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_5_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_6_), .S(DP_w_5_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_6 ( .A(DP_fb_6_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_6_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_6_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_7_), .S(DP_w_6_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_7 ( .A(DP_fb_7_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_7_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_7_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_8_), .S(DP_w_7_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_8 ( .A(DP_fb_8_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_8_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_8_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_9_), .S(DP_w_8_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_9 ( .A(DP_fb_9_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_9_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_9_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_10_), .S(DP_w_9_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_10 ( .A(DP_fb_10_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_10_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_10_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_11_), .S(DP_w_10_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_11 ( .A(DP_fb_11_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_12_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_11_), .CO(
        DP_sub_0_root_sub_0_root_sub_104_carry_12_), .S(DP_w_11_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_104_U2_12 ( .A(DP_fb_12_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_12_), .CI(
        DP_sub_0_root_sub_0_root_sub_104_carry_12_), .S(DP_w_12_) );
  XOR2_X1 DP_mult_97_U563 ( .A(DP_a_int[21]), .B(DP_a_int[22]), .Z(
        DP_mult_97_n653) );
  INV_X1 DP_mult_97_U562 ( .A(DP_a_int[22]), .ZN(DP_mult_97_n543) );
  NOR2_X1 DP_mult_97_U561 ( .A1(DP_mult_97_n543), .A2(DP_sw1_1_), .ZN(
        DP_mult_97_n658) );
  INV_X1 DP_mult_97_U560 ( .A(DP_mult_97_n658), .ZN(DP_mult_97_n660) );
  NAND2_X1 DP_mult_97_U559 ( .A1(DP_a_int[22]), .A2(DP_mult_97_n532), .ZN(
        DP_mult_97_n530) );
  XNOR2_X1 DP_mult_97_U558 ( .A(DP_sw1_2_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n529) );
  OAI22_X1 DP_mult_97_U557 ( .A1(DP_mult_97_n660), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n529), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n659) );
  NAND2_X1 DP_mult_97_U556 ( .A1(DP_mult_97_n653), .A2(DP_mult_97_n659), .ZN(
        DP_mult_97_n656) );
  NAND2_X1 DP_mult_97_U555 ( .A1(DP_mult_97_n658), .A2(DP_mult_97_n659), .ZN(
        DP_mult_97_n657) );
  INV_X1 DP_mult_97_U554 ( .A(DP_sw1_0_), .ZN(DP_mult_97_n560) );
  MUX2_X1 DP_mult_97_U553 ( .A(DP_mult_97_n656), .B(DP_mult_97_n657), .S(
        DP_mult_97_n560), .Z(DP_mult_97_n655) );
  INV_X1 DP_mult_97_U552 ( .A(DP_mult_97_n655), .ZN(DP_mult_97_n650) );
  INV_X1 DP_mult_97_U551 ( .A(DP_a_int[20]), .ZN(DP_mult_97_n632) );
  XNOR2_X1 DP_mult_97_U550 ( .A(DP_mult_97_n632), .B(DP_a_int[21]), .ZN(
        DP_mult_97_n654) );
  NAND2_X1 DP_mult_97_U549 ( .A1(DP_mult_97_n546), .A2(DP_mult_97_n654), .ZN(
        DP_mult_97_n545) );
  NAND3_X1 DP_mult_97_U548 ( .A1(DP_mult_97_n653), .A2(DP_mult_97_n560), .A3(
        DP_a_int[20]), .ZN(DP_mult_97_n652) );
  OAI21_X1 DP_mult_97_U547 ( .B1(DP_mult_97_n632), .B2(DP_mult_97_n545), .A(
        DP_mult_97_n652), .ZN(DP_mult_97_n651) );
  AOI222_X1 DP_mult_97_U546 ( .A1(DP_mult_97_n650), .A2(DP_mult_97_n255), .B1(
        DP_mult_97_n651), .B2(DP_mult_97_n650), .C1(DP_mult_97_n651), .C2(
        DP_mult_97_n255), .ZN(DP_mult_97_n649) );
  INV_X1 DP_mult_97_U545 ( .A(DP_mult_97_n649), .ZN(DP_mult_97_n648) );
  AOI222_X1 DP_mult_97_U544 ( .A1(DP_mult_97_n648), .A2(DP_mult_97_n253), .B1(
        DP_mult_97_n648), .B2(DP_mult_97_n254), .C1(DP_mult_97_n254), .C2(
        DP_mult_97_n253), .ZN(DP_mult_97_n647) );
  INV_X1 DP_mult_97_U543 ( .A(DP_mult_97_n647), .ZN(DP_mult_97_n646) );
  AOI222_X1 DP_mult_97_U542 ( .A1(DP_mult_97_n646), .A2(DP_mult_97_n249), .B1(
        DP_mult_97_n646), .B2(DP_mult_97_n252), .C1(DP_mult_97_n252), .C2(
        DP_mult_97_n249), .ZN(DP_mult_97_n645) );
  INV_X1 DP_mult_97_U541 ( .A(DP_mult_97_n645), .ZN(DP_mult_97_n644) );
  AOI222_X1 DP_mult_97_U540 ( .A1(DP_mult_97_n644), .A2(DP_mult_97_n245), .B1(
        DP_mult_97_n644), .B2(DP_mult_97_n248), .C1(DP_mult_97_n248), .C2(
        DP_mult_97_n245), .ZN(DP_mult_97_n643) );
  INV_X1 DP_mult_97_U539 ( .A(DP_mult_97_n643), .ZN(DP_mult_97_n642) );
  AOI222_X1 DP_mult_97_U538 ( .A1(DP_mult_97_n642), .A2(DP_mult_97_n239), .B1(
        DP_mult_97_n642), .B2(DP_mult_97_n244), .C1(DP_mult_97_n244), .C2(
        DP_mult_97_n239), .ZN(DP_mult_97_n639) );
  INV_X1 DP_mult_97_U537 ( .A(DP_mult_97_n233), .ZN(DP_mult_97_n640) );
  INV_X1 DP_mult_97_U536 ( .A(DP_mult_97_n238), .ZN(DP_mult_97_n641) );
  OAI222_X1 DP_mult_97_U535 ( .A1(DP_mult_97_n639), .A2(DP_mult_97_n640), .B1(
        DP_mult_97_n639), .B2(DP_mult_97_n641), .C1(DP_mult_97_n641), .C2(
        DP_mult_97_n640), .ZN(DP_mult_97_n638) );
  AOI222_X1 DP_mult_97_U534 ( .A1(DP_mult_97_n638), .A2(DP_mult_97_n225), .B1(
        DP_mult_97_n638), .B2(DP_mult_97_n232), .C1(DP_mult_97_n232), .C2(
        DP_mult_97_n225), .ZN(DP_mult_97_n635) );
  INV_X1 DP_mult_97_U533 ( .A(DP_mult_97_n217), .ZN(DP_mult_97_n636) );
  INV_X1 DP_mult_97_U532 ( .A(DP_mult_97_n224), .ZN(DP_mult_97_n637) );
  OAI222_X1 DP_mult_97_U531 ( .A1(DP_mult_97_n635), .A2(DP_mult_97_n636), .B1(
        DP_mult_97_n635), .B2(DP_mult_97_n637), .C1(DP_mult_97_n637), .C2(
        DP_mult_97_n636), .ZN(DP_mult_97_n126) );
  XNOR2_X1 DP_mult_97_U530 ( .A(DP_sw1_11_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n606) );
  INV_X1 DP_mult_97_U529 ( .A(DP_a_int[16]), .ZN(DP_mult_97_n622) );
  INV_X1 DP_mult_97_U528 ( .A(DP_a_int[14]), .ZN(DP_mult_97_n624) );
  XNOR2_X1 DP_mult_97_U527 ( .A(DP_mult_97_n624), .B(DP_a_int[15]), .ZN(
        DP_mult_97_n634) );
  NAND2_X1 DP_mult_97_U526 ( .A1(DP_mult_97_n593), .A2(DP_mult_97_n634), .ZN(
        DP_mult_97_n595) );
  XNOR2_X1 DP_mult_97_U525 ( .A(DP_sw1_12_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n608) );
  OAI22_X1 DP_mult_97_U524 ( .A1(DP_mult_97_n606), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n608), .ZN(DP_mult_97_n142) );
  INV_X1 DP_mult_97_U523 ( .A(DP_mult_97_n142), .ZN(DP_mult_97_n143) );
  XNOR2_X1 DP_mult_97_U522 ( .A(DP_sw1_11_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n590) );
  INV_X1 DP_mult_97_U521 ( .A(DP_a_int[18]), .ZN(DP_mult_97_n620) );
  XNOR2_X1 DP_mult_97_U520 ( .A(DP_mult_97_n622), .B(DP_a_int[17]), .ZN(
        DP_mult_97_n633) );
  NAND2_X1 DP_mult_97_U519 ( .A1(DP_mult_97_n577), .A2(DP_mult_97_n633), .ZN(
        DP_mult_97_n579) );
  XNOR2_X1 DP_mult_97_U518 ( .A(DP_sw1_12_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n592) );
  OAI22_X1 DP_mult_97_U517 ( .A1(DP_mult_97_n590), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n592), .ZN(DP_mult_97_n152) );
  INV_X1 DP_mult_97_U516 ( .A(DP_mult_97_n152), .ZN(DP_mult_97_n153) );
  XNOR2_X1 DP_mult_97_U515 ( .A(DP_sw1_11_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n574) );
  XNOR2_X1 DP_mult_97_U514 ( .A(DP_mult_97_n620), .B(DP_a_int[19]), .ZN(
        DP_mult_97_n631) );
  NAND2_X1 DP_mult_97_U513 ( .A1(DP_mult_97_n561), .A2(DP_mult_97_n631), .ZN(
        DP_mult_97_n563) );
  XNOR2_X1 DP_mult_97_U512 ( .A(DP_sw1_12_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n576) );
  OAI22_X1 DP_mult_97_U511 ( .A1(DP_mult_97_n574), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n576), .ZN(DP_mult_97_n166) );
  INV_X1 DP_mult_97_U510 ( .A(DP_mult_97_n166), .ZN(DP_mult_97_n167) );
  XNOR2_X1 DP_mult_97_U509 ( .A(DP_sw1_11_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n557) );
  XNOR2_X1 DP_mult_97_U508 ( .A(DP_sw1_12_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n559) );
  OAI22_X1 DP_mult_97_U507 ( .A1(DP_mult_97_n557), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n559), .ZN(DP_mult_97_n184) );
  INV_X1 DP_mult_97_U506 ( .A(DP_mult_97_n184), .ZN(DP_mult_97_n185) );
  XNOR2_X1 DP_mult_97_U505 ( .A(DP_sw1_4_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n599) );
  XNOR2_X1 DP_mult_97_U504 ( .A(DP_sw1_5_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n600) );
  OAI22_X1 DP_mult_97_U503 ( .A1(DP_mult_97_n599), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n600), .ZN(DP_mult_97_n629) );
  XNOR2_X1 DP_mult_97_U502 ( .A(DP_sw1_8_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n571) );
  XNOR2_X1 DP_mult_97_U501 ( .A(DP_sw1_9_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n572) );
  OAI22_X1 DP_mult_97_U500 ( .A1(DP_mult_97_n571), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n572), .ZN(DP_mult_97_n630) );
  OR2_X1 DP_mult_97_U499 ( .A1(DP_mult_97_n629), .A2(DP_mult_97_n630), .ZN(
        DP_mult_97_n194) );
  XNOR2_X1 DP_mult_97_U498 ( .A(DP_mult_97_n629), .B(DP_mult_97_n630), .ZN(
        DP_mult_97_n195) );
  INV_X1 DP_mult_97_U497 ( .A(DP_a_int[12]), .ZN(DP_mult_97_n626) );
  XNOR2_X1 DP_mult_97_U496 ( .A(DP_mult_97_n626), .B(DP_a_int[13]), .ZN(
        DP_mult_97_n628) );
  NAND2_X1 DP_mult_97_U495 ( .A1(DP_mult_97_n526), .A2(DP_mult_97_n628), .ZN(
        DP_mult_97_n525) );
  OR3_X1 DP_mult_97_U494 ( .A1(DP_mult_97_n526), .A2(DP_sw1_0_), .A3(
        DP_mult_97_n626), .ZN(DP_mult_97_n627) );
  OAI21_X1 DP_mult_97_U493 ( .B1(DP_mult_97_n626), .B2(DP_mult_97_n525), .A(
        DP_mult_97_n627), .ZN(DP_mult_97_n256) );
  OR3_X1 DP_mult_97_U492 ( .A1(DP_mult_97_n593), .A2(DP_sw1_0_), .A3(
        DP_mult_97_n624), .ZN(DP_mult_97_n625) );
  OAI21_X1 DP_mult_97_U491 ( .B1(DP_mult_97_n624), .B2(DP_mult_97_n595), .A(
        DP_mult_97_n625), .ZN(DP_mult_97_n257) );
  OR3_X1 DP_mult_97_U490 ( .A1(DP_mult_97_n577), .A2(DP_sw1_0_), .A3(
        DP_mult_97_n622), .ZN(DP_mult_97_n623) );
  OAI21_X1 DP_mult_97_U489 ( .B1(DP_mult_97_n622), .B2(DP_mult_97_n579), .A(
        DP_mult_97_n623), .ZN(DP_mult_97_n258) );
  OR3_X1 DP_mult_97_U488 ( .A1(DP_mult_97_n561), .A2(DP_sw1_0_), .A3(
        DP_mult_97_n620), .ZN(DP_mult_97_n621) );
  OAI21_X1 DP_mult_97_U487 ( .B1(DP_mult_97_n620), .B2(DP_mult_97_n563), .A(
        DP_mult_97_n621), .ZN(DP_mult_97_n259) );
  XNOR2_X1 DP_mult_97_U486 ( .A(DP_sw1_10_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n619) );
  XNOR2_X1 DP_mult_97_U485 ( .A(DP_sw1_11_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n528) );
  OAI22_X1 DP_mult_97_U484 ( .A1(DP_mult_97_n619), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n528), .ZN(DP_mult_97_n263) );
  XNOR2_X1 DP_mult_97_U483 ( .A(DP_sw1_9_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n618) );
  OAI22_X1 DP_mult_97_U482 ( .A1(DP_mult_97_n618), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n619), .ZN(DP_mult_97_n264) );
  XNOR2_X1 DP_mult_97_U481 ( .A(DP_sw1_8_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n617) );
  OAI22_X1 DP_mult_97_U480 ( .A1(DP_mult_97_n617), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n618), .ZN(DP_mult_97_n265) );
  XNOR2_X1 DP_mult_97_U479 ( .A(DP_sw1_7_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n616) );
  OAI22_X1 DP_mult_97_U478 ( .A1(DP_mult_97_n616), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n617), .ZN(DP_mult_97_n266) );
  XNOR2_X1 DP_mult_97_U477 ( .A(DP_sw1_6_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n615) );
  OAI22_X1 DP_mult_97_U476 ( .A1(DP_mult_97_n615), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n616), .ZN(DP_mult_97_n267) );
  XNOR2_X1 DP_mult_97_U475 ( .A(DP_sw1_5_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n614) );
  OAI22_X1 DP_mult_97_U474 ( .A1(DP_mult_97_n614), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n615), .ZN(DP_mult_97_n268) );
  XNOR2_X1 DP_mult_97_U473 ( .A(DP_sw1_4_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n613) );
  OAI22_X1 DP_mult_97_U472 ( .A1(DP_mult_97_n613), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n614), .ZN(DP_mult_97_n269) );
  XNOR2_X1 DP_mult_97_U471 ( .A(DP_sw1_3_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n612) );
  OAI22_X1 DP_mult_97_U470 ( .A1(DP_mult_97_n612), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n613), .ZN(DP_mult_97_n270) );
  XNOR2_X1 DP_mult_97_U469 ( .A(DP_sw1_2_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n611) );
  OAI22_X1 DP_mult_97_U468 ( .A1(DP_mult_97_n611), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n612), .ZN(DP_mult_97_n271) );
  XNOR2_X1 DP_mult_97_U467 ( .A(DP_sw1_1_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n610) );
  OAI22_X1 DP_mult_97_U466 ( .A1(DP_mult_97_n610), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n611), .ZN(DP_mult_97_n272) );
  XNOR2_X1 DP_mult_97_U465 ( .A(DP_sw1_0_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n609) );
  OAI22_X1 DP_mult_97_U464 ( .A1(DP_mult_97_n609), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n610), .ZN(DP_mult_97_n273) );
  NOR2_X1 DP_mult_97_U463 ( .A1(DP_mult_97_n560), .A2(DP_mult_97_n526), .ZN(
        DP_mult_97_n274) );
  AOI21_X1 DP_mult_97_U462 ( .B1(DP_mult_97_n595), .B2(DP_mult_97_n593), .A(
        DP_mult_97_n608), .ZN(DP_mult_97_n607) );
  INV_X1 DP_mult_97_U461 ( .A(DP_mult_97_n607), .ZN(DP_mult_97_n275) );
  XNOR2_X1 DP_mult_97_U460 ( .A(DP_sw1_10_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n605) );
  OAI22_X1 DP_mult_97_U459 ( .A1(DP_mult_97_n605), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n606), .ZN(DP_mult_97_n276) );
  XNOR2_X1 DP_mult_97_U458 ( .A(DP_sw1_9_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n604) );
  OAI22_X1 DP_mult_97_U457 ( .A1(DP_mult_97_n604), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n605), .ZN(DP_mult_97_n277) );
  XNOR2_X1 DP_mult_97_U456 ( .A(DP_sw1_8_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n603) );
  OAI22_X1 DP_mult_97_U455 ( .A1(DP_mult_97_n603), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n604), .ZN(DP_mult_97_n278) );
  XNOR2_X1 DP_mult_97_U454 ( .A(DP_sw1_7_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n602) );
  OAI22_X1 DP_mult_97_U453 ( .A1(DP_mult_97_n602), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n603), .ZN(DP_mult_97_n279) );
  XNOR2_X1 DP_mult_97_U452 ( .A(DP_sw1_6_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n601) );
  OAI22_X1 DP_mult_97_U451 ( .A1(DP_mult_97_n601), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n602), .ZN(DP_mult_97_n280) );
  OAI22_X1 DP_mult_97_U450 ( .A1(DP_mult_97_n600), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n601), .ZN(DP_mult_97_n281) );
  XNOR2_X1 DP_mult_97_U449 ( .A(DP_sw1_3_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n598) );
  OAI22_X1 DP_mult_97_U448 ( .A1(DP_mult_97_n598), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n599), .ZN(DP_mult_97_n283) );
  XNOR2_X1 DP_mult_97_U447 ( .A(DP_sw1_2_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n597) );
  OAI22_X1 DP_mult_97_U446 ( .A1(DP_mult_97_n597), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n598), .ZN(DP_mult_97_n284) );
  XNOR2_X1 DP_mult_97_U445 ( .A(DP_sw1_1_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n596) );
  OAI22_X1 DP_mult_97_U444 ( .A1(DP_mult_97_n596), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n597), .ZN(DP_mult_97_n285) );
  XNOR2_X1 DP_mult_97_U443 ( .A(DP_sw1_0_), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n594) );
  OAI22_X1 DP_mult_97_U442 ( .A1(DP_mult_97_n594), .A2(DP_mult_97_n595), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n286) );
  NOR2_X1 DP_mult_97_U441 ( .A1(DP_mult_97_n560), .A2(DP_mult_97_n593), .ZN(
        DP_mult_97_n287) );
  AOI21_X1 DP_mult_97_U440 ( .B1(DP_mult_97_n579), .B2(DP_mult_97_n577), .A(
        DP_mult_97_n592), .ZN(DP_mult_97_n591) );
  INV_X1 DP_mult_97_U439 ( .A(DP_mult_97_n591), .ZN(DP_mult_97_n288) );
  XNOR2_X1 DP_mult_97_U438 ( .A(DP_sw1_10_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n589) );
  OAI22_X1 DP_mult_97_U437 ( .A1(DP_mult_97_n589), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n590), .ZN(DP_mult_97_n289) );
  XNOR2_X1 DP_mult_97_U436 ( .A(DP_sw1_9_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n588) );
  OAI22_X1 DP_mult_97_U435 ( .A1(DP_mult_97_n588), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n589), .ZN(DP_mult_97_n290) );
  XNOR2_X1 DP_mult_97_U434 ( .A(DP_sw1_8_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n587) );
  OAI22_X1 DP_mult_97_U433 ( .A1(DP_mult_97_n587), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n588), .ZN(DP_mult_97_n291) );
  XNOR2_X1 DP_mult_97_U432 ( .A(DP_sw1_7_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n586) );
  OAI22_X1 DP_mult_97_U431 ( .A1(DP_mult_97_n586), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n587), .ZN(DP_mult_97_n292) );
  XNOR2_X1 DP_mult_97_U430 ( .A(DP_sw1_6_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n585) );
  OAI22_X1 DP_mult_97_U429 ( .A1(DP_mult_97_n585), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n586), .ZN(DP_mult_97_n293) );
  XNOR2_X1 DP_mult_97_U428 ( .A(DP_sw1_5_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n584) );
  OAI22_X1 DP_mult_97_U427 ( .A1(DP_mult_97_n584), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n585), .ZN(DP_mult_97_n294) );
  XNOR2_X1 DP_mult_97_U426 ( .A(DP_sw1_4_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n583) );
  OAI22_X1 DP_mult_97_U425 ( .A1(DP_mult_97_n583), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n584), .ZN(DP_mult_97_n295) );
  XNOR2_X1 DP_mult_97_U424 ( .A(DP_sw1_3_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n582) );
  OAI22_X1 DP_mult_97_U423 ( .A1(DP_mult_97_n582), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n583), .ZN(DP_mult_97_n296) );
  XNOR2_X1 DP_mult_97_U422 ( .A(DP_sw1_2_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n581) );
  OAI22_X1 DP_mult_97_U421 ( .A1(DP_mult_97_n581), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n582), .ZN(DP_mult_97_n297) );
  XNOR2_X1 DP_mult_97_U420 ( .A(DP_sw1_1_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n580) );
  OAI22_X1 DP_mult_97_U419 ( .A1(DP_mult_97_n580), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n581), .ZN(DP_mult_97_n298) );
  XNOR2_X1 DP_mult_97_U418 ( .A(DP_sw1_0_), .B(DP_a_int[16]), .ZN(
        DP_mult_97_n578) );
  OAI22_X1 DP_mult_97_U417 ( .A1(DP_mult_97_n578), .A2(DP_mult_97_n579), .B1(
        DP_mult_97_n577), .B2(DP_mult_97_n580), .ZN(DP_mult_97_n299) );
  NOR2_X1 DP_mult_97_U416 ( .A1(DP_mult_97_n560), .A2(DP_mult_97_n577), .ZN(
        DP_mult_97_n300) );
  AOI21_X1 DP_mult_97_U415 ( .B1(DP_mult_97_n563), .B2(DP_mult_97_n561), .A(
        DP_mult_97_n576), .ZN(DP_mult_97_n575) );
  INV_X1 DP_mult_97_U414 ( .A(DP_mult_97_n575), .ZN(DP_mult_97_n301) );
  XNOR2_X1 DP_mult_97_U413 ( .A(DP_sw1_10_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n573) );
  OAI22_X1 DP_mult_97_U412 ( .A1(DP_mult_97_n573), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n574), .ZN(DP_mult_97_n302) );
  OAI22_X1 DP_mult_97_U411 ( .A1(DP_mult_97_n572), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n573), .ZN(DP_mult_97_n303) );
  XNOR2_X1 DP_mult_97_U410 ( .A(DP_sw1_7_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n570) );
  OAI22_X1 DP_mult_97_U409 ( .A1(DP_mult_97_n570), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n571), .ZN(DP_mult_97_n305) );
  XNOR2_X1 DP_mult_97_U408 ( .A(DP_sw1_6_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n569) );
  OAI22_X1 DP_mult_97_U407 ( .A1(DP_mult_97_n569), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n570), .ZN(DP_mult_97_n306) );
  XNOR2_X1 DP_mult_97_U406 ( .A(DP_sw1_5_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n568) );
  OAI22_X1 DP_mult_97_U405 ( .A1(DP_mult_97_n568), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n569), .ZN(DP_mult_97_n307) );
  XNOR2_X1 DP_mult_97_U404 ( .A(DP_sw1_4_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n567) );
  OAI22_X1 DP_mult_97_U403 ( .A1(DP_mult_97_n567), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n568), .ZN(DP_mult_97_n308) );
  XNOR2_X1 DP_mult_97_U402 ( .A(DP_sw1_3_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n566) );
  OAI22_X1 DP_mult_97_U401 ( .A1(DP_mult_97_n566), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n567), .ZN(DP_mult_97_n309) );
  XNOR2_X1 DP_mult_97_U400 ( .A(DP_sw1_2_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n565) );
  OAI22_X1 DP_mult_97_U399 ( .A1(DP_mult_97_n565), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n566), .ZN(DP_mult_97_n310) );
  XNOR2_X1 DP_mult_97_U398 ( .A(DP_sw1_1_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n564) );
  OAI22_X1 DP_mult_97_U397 ( .A1(DP_mult_97_n564), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n565), .ZN(DP_mult_97_n311) );
  XNOR2_X1 DP_mult_97_U396 ( .A(DP_sw1_0_), .B(DP_a_int[18]), .ZN(
        DP_mult_97_n562) );
  OAI22_X1 DP_mult_97_U395 ( .A1(DP_mult_97_n562), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n564), .ZN(DP_mult_97_n312) );
  NOR2_X1 DP_mult_97_U394 ( .A1(DP_mult_97_n560), .A2(DP_mult_97_n561), .ZN(
        DP_mult_97_n313) );
  AOI21_X1 DP_mult_97_U393 ( .B1(DP_mult_97_n545), .B2(DP_mult_97_n546), .A(
        DP_mult_97_n559), .ZN(DP_mult_97_n558) );
  INV_X1 DP_mult_97_U392 ( .A(DP_mult_97_n558), .ZN(DP_mult_97_n314) );
  XNOR2_X1 DP_mult_97_U391 ( .A(DP_sw1_10_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n556) );
  OAI22_X1 DP_mult_97_U390 ( .A1(DP_mult_97_n556), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n557), .ZN(DP_mult_97_n315) );
  XNOR2_X1 DP_mult_97_U389 ( .A(DP_sw1_9_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n555) );
  OAI22_X1 DP_mult_97_U388 ( .A1(DP_mult_97_n555), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n556), .ZN(DP_mult_97_n316) );
  XNOR2_X1 DP_mult_97_U387 ( .A(DP_sw1_8_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n554) );
  OAI22_X1 DP_mult_97_U386 ( .A1(DP_mult_97_n554), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n555), .ZN(DP_mult_97_n317) );
  XNOR2_X1 DP_mult_97_U385 ( .A(DP_sw1_7_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n553) );
  OAI22_X1 DP_mult_97_U384 ( .A1(DP_mult_97_n553), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n554), .ZN(DP_mult_97_n318) );
  XNOR2_X1 DP_mult_97_U383 ( .A(DP_sw1_6_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n552) );
  OAI22_X1 DP_mult_97_U382 ( .A1(DP_mult_97_n552), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n553), .ZN(DP_mult_97_n319) );
  XNOR2_X1 DP_mult_97_U381 ( .A(DP_sw1_5_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n551) );
  OAI22_X1 DP_mult_97_U380 ( .A1(DP_mult_97_n551), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n552), .ZN(DP_mult_97_n320) );
  XNOR2_X1 DP_mult_97_U379 ( .A(DP_sw1_4_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n550) );
  OAI22_X1 DP_mult_97_U378 ( .A1(DP_mult_97_n550), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n551), .ZN(DP_mult_97_n321) );
  XNOR2_X1 DP_mult_97_U377 ( .A(DP_sw1_3_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n549) );
  OAI22_X1 DP_mult_97_U376 ( .A1(DP_mult_97_n549), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n550), .ZN(DP_mult_97_n322) );
  XNOR2_X1 DP_mult_97_U375 ( .A(DP_sw1_2_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n548) );
  OAI22_X1 DP_mult_97_U374 ( .A1(DP_mult_97_n548), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n549), .ZN(DP_mult_97_n323) );
  XNOR2_X1 DP_mult_97_U373 ( .A(DP_sw1_1_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n547) );
  OAI22_X1 DP_mult_97_U372 ( .A1(DP_mult_97_n547), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n548), .ZN(DP_mult_97_n324) );
  XNOR2_X1 DP_mult_97_U371 ( .A(DP_sw1_0_), .B(DP_a_int[20]), .ZN(
        DP_mult_97_n544) );
  OAI22_X1 DP_mult_97_U370 ( .A1(DP_mult_97_n544), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n546), .B2(DP_mult_97_n547), .ZN(DP_mult_97_n325) );
  XOR2_X1 DP_mult_97_U369 ( .A(DP_sw1_12_), .B(DP_mult_97_n543), .Z(
        DP_mult_97_n541) );
  AOI21_X1 DP_mult_97_U368 ( .B1(DP_mult_97_n530), .B2(DP_mult_97_n532), .A(
        DP_mult_97_n541), .ZN(DP_mult_97_n542) );
  INV_X1 DP_mult_97_U367 ( .A(DP_mult_97_n542), .ZN(DP_mult_97_n327) );
  XNOR2_X1 DP_mult_97_U366 ( .A(DP_sw1_11_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n540) );
  OAI22_X1 DP_mult_97_U365 ( .A1(DP_mult_97_n540), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n541), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n328) );
  XNOR2_X1 DP_mult_97_U364 ( .A(DP_sw1_10_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n539) );
  OAI22_X1 DP_mult_97_U363 ( .A1(DP_mult_97_n539), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n540), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n329) );
  XNOR2_X1 DP_mult_97_U362 ( .A(DP_sw1_9_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n538) );
  OAI22_X1 DP_mult_97_U361 ( .A1(DP_mult_97_n538), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n539), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n330) );
  XNOR2_X1 DP_mult_97_U360 ( .A(DP_sw1_8_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n537) );
  OAI22_X1 DP_mult_97_U359 ( .A1(DP_mult_97_n537), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n538), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n331) );
  XNOR2_X1 DP_mult_97_U358 ( .A(DP_sw1_7_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n536) );
  OAI22_X1 DP_mult_97_U357 ( .A1(DP_mult_97_n536), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n537), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n332) );
  XNOR2_X1 DP_mult_97_U356 ( .A(DP_sw1_6_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n535) );
  OAI22_X1 DP_mult_97_U355 ( .A1(DP_mult_97_n535), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n536), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n333) );
  XNOR2_X1 DP_mult_97_U354 ( .A(DP_sw1_5_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n534) );
  OAI22_X1 DP_mult_97_U353 ( .A1(DP_mult_97_n534), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n535), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n334) );
  XNOR2_X1 DP_mult_97_U352 ( .A(DP_sw1_4_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n533) );
  OAI22_X1 DP_mult_97_U351 ( .A1(DP_mult_97_n533), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n534), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n335) );
  XNOR2_X1 DP_mult_97_U350 ( .A(DP_sw1_3_), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n531) );
  OAI22_X1 DP_mult_97_U349 ( .A1(DP_mult_97_n531), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n533), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n336) );
  OAI22_X1 DP_mult_97_U348 ( .A1(DP_mult_97_n529), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n531), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n337) );
  XNOR2_X1 DP_mult_97_U347 ( .A(DP_sw1_12_), .B(DP_a_int[12]), .ZN(
        DP_mult_97_n527) );
  OAI22_X1 DP_mult_97_U346 ( .A1(DP_mult_97_n528), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n526), .B2(DP_mult_97_n527), .ZN(DP_mult_97_n519) );
  AOI21_X1 DP_mult_97_U345 ( .B1(DP_mult_97_n525), .B2(DP_mult_97_n526), .A(
        DP_mult_97_n527), .ZN(DP_mult_97_n522) );
  INV_X1 DP_mult_97_U344 ( .A(DP_mult_97_n522), .ZN(DP_mult_97_n520) );
  INV_X1 DP_mult_97_U343 ( .A(DP_mult_97_n519), .ZN(DP_mult_97_n524) );
  AOI222_X1 DP_mult_97_U342 ( .A1(DP_mult_97_n115), .A2(DP_mult_97_n138), .B1(
        DP_mult_97_n524), .B2(DP_mult_97_n115), .C1(DP_mult_97_n524), .C2(
        DP_mult_97_n138), .ZN(DP_mult_97_n523) );
  OAI22_X1 DP_mult_97_U341 ( .A1(DP_mult_97_n522), .A2(DP_mult_97_n523), .B1(
        DP_mult_97_n524), .B2(DP_mult_97_n523), .ZN(DP_mult_97_n521) );
  AOI21_X1 DP_mult_97_U340 ( .B1(DP_mult_97_n519), .B2(DP_mult_97_n520), .A(
        DP_mult_97_n521), .ZN(DP_sw1_a2_11_) );
  XOR2_X2 DP_mult_97_U339 ( .A(DP_a_int[15]), .B(DP_mult_97_n622), .Z(
        DP_mult_97_n593) );
  XOR2_X2 DP_mult_97_U338 ( .A(DP_a_int[17]), .B(DP_mult_97_n620), .Z(
        DP_mult_97_n577) );
  XOR2_X2 DP_mult_97_U337 ( .A(DP_a_int[19]), .B(DP_mult_97_n632), .Z(
        DP_mult_97_n561) );
  XOR2_X2 DP_mult_97_U336 ( .A(DP_a_int[13]), .B(DP_mult_97_n624), .Z(
        DP_mult_97_n526) );
  INV_X1 DP_mult_97_U335 ( .A(DP_a_int[23]), .ZN(DP_mult_97_n532) );
  INV_X1 DP_mult_97_U334 ( .A(DP_mult_97_n653), .ZN(DP_mult_97_n546) );
  HA_X1 DP_mult_97_U120 ( .A(DP_mult_97_n325), .B(DP_mult_97_n337), .CO(
        DP_mult_97_n254), .S(DP_mult_97_n255) );
  FA_X1 DP_mult_97_U119 ( .A(DP_mult_97_n336), .B(DP_mult_97_n313), .CI(
        DP_mult_97_n324), .CO(DP_mult_97_n252), .S(DP_mult_97_n253) );
  HA_X1 DP_mult_97_U118 ( .A(DP_mult_97_n259), .B(DP_mult_97_n312), .CO(
        DP_mult_97_n250), .S(DP_mult_97_n251) );
  FA_X1 DP_mult_97_U117 ( .A(DP_mult_97_n323), .B(DP_mult_97_n335), .CI(
        DP_mult_97_n251), .CO(DP_mult_97_n248), .S(DP_mult_97_n249) );
  FA_X1 DP_mult_97_U109 ( .A(DP_mult_97_n334), .B(DP_mult_97_n300), .CI(
        DP_mult_97_n322), .CO(DP_mult_97_n246), .S(DP_mult_97_n247) );
  FA_X1 DP_mult_97_U108 ( .A(DP_mult_97_n250), .B(DP_mult_97_n311), .CI(
        DP_mult_97_n247), .CO(DP_mult_97_n244), .S(DP_mult_97_n245) );
  HA_X1 DP_mult_97_U107 ( .A(DP_mult_97_n258), .B(DP_mult_97_n299), .CO(
        DP_mult_97_n242), .S(DP_mult_97_n243) );
  FA_X1 DP_mult_97_U106 ( .A(DP_mult_97_n310), .B(DP_mult_97_n333), .CI(
        DP_mult_97_n321), .CO(DP_mult_97_n240), .S(DP_mult_97_n241) );
  FA_X1 DP_mult_97_U105 ( .A(DP_mult_97_n246), .B(DP_mult_97_n243), .CI(
        DP_mult_97_n241), .CO(DP_mult_97_n238), .S(DP_mult_97_n239) );
  FA_X1 DP_mult_97_U104 ( .A(DP_mult_97_n309), .B(DP_mult_97_n287), .CI(
        DP_mult_97_n332), .CO(DP_mult_97_n236), .S(DP_mult_97_n237) );
  FA_X1 DP_mult_97_U103 ( .A(DP_mult_97_n298), .B(DP_mult_97_n320), .CI(
        DP_mult_97_n242), .CO(DP_mult_97_n234), .S(DP_mult_97_n235) );
  FA_X1 DP_mult_97_U102 ( .A(DP_mult_97_n237), .B(DP_mult_97_n240), .CI(
        DP_mult_97_n235), .CO(DP_mult_97_n232), .S(DP_mult_97_n233) );
  HA_X1 DP_mult_97_U101 ( .A(DP_mult_97_n257), .B(DP_mult_97_n286), .CO(
        DP_mult_97_n230), .S(DP_mult_97_n231) );
  FA_X1 DP_mult_97_U100 ( .A(DP_mult_97_n297), .B(DP_mult_97_n308), .CI(
        DP_mult_97_n319), .CO(DP_mult_97_n228), .S(DP_mult_97_n229) );
  FA_X1 DP_mult_97_U99 ( .A(DP_mult_97_n231), .B(DP_mult_97_n331), .CI(
        DP_mult_97_n236), .CO(DP_mult_97_n226), .S(DP_mult_97_n227) );
  FA_X1 DP_mult_97_U98 ( .A(DP_mult_97_n229), .B(DP_mult_97_n234), .CI(
        DP_mult_97_n227), .CO(DP_mult_97_n224), .S(DP_mult_97_n225) );
  FA_X1 DP_mult_97_U97 ( .A(DP_mult_97_n296), .B(DP_mult_97_n274), .CI(
        DP_mult_97_n330), .CO(DP_mult_97_n222), .S(DP_mult_97_n223) );
  FA_X1 DP_mult_97_U96 ( .A(DP_mult_97_n285), .B(DP_mult_97_n318), .CI(
        DP_mult_97_n307), .CO(DP_mult_97_n220), .S(DP_mult_97_n221) );
  FA_X1 DP_mult_97_U95 ( .A(DP_mult_97_n228), .B(DP_mult_97_n230), .CI(
        DP_mult_97_n223), .CO(DP_mult_97_n218), .S(DP_mult_97_n219) );
  FA_X1 DP_mult_97_U94 ( .A(DP_mult_97_n226), .B(DP_mult_97_n221), .CI(
        DP_mult_97_n219), .CO(DP_mult_97_n216), .S(DP_mult_97_n217) );
  HA_X1 DP_mult_97_U93 ( .A(DP_mult_97_n256), .B(DP_mult_97_n273), .CO(
        DP_mult_97_n214), .S(DP_mult_97_n215) );
  FA_X1 DP_mult_97_U92 ( .A(DP_mult_97_n284), .B(DP_mult_97_n306), .CI(
        DP_mult_97_n329), .CO(DP_mult_97_n212), .S(DP_mult_97_n213) );
  FA_X1 DP_mult_97_U91 ( .A(DP_mult_97_n295), .B(DP_mult_97_n317), .CI(
        DP_mult_97_n215), .CO(DP_mult_97_n210), .S(DP_mult_97_n211) );
  FA_X1 DP_mult_97_U90 ( .A(DP_mult_97_n220), .B(DP_mult_97_n222), .CI(
        DP_mult_97_n213), .CO(DP_mult_97_n208), .S(DP_mult_97_n209) );
  FA_X1 DP_mult_97_U89 ( .A(DP_mult_97_n218), .B(DP_mult_97_n211), .CI(
        DP_mult_97_n209), .CO(DP_mult_97_n206), .S(DP_mult_97_n207) );
  HA_X1 DP_mult_97_U88 ( .A(DP_mult_97_n272), .B(DP_mult_97_n283), .CO(
        DP_mult_97_n204), .S(DP_mult_97_n205) );
  FA_X1 DP_mult_97_U87 ( .A(DP_mult_97_n328), .B(DP_mult_97_n305), .CI(
        DP_mult_97_n294), .CO(DP_mult_97_n202), .S(DP_mult_97_n203) );
  FA_X1 DP_mult_97_U86 ( .A(DP_mult_97_n214), .B(DP_mult_97_n316), .CI(
        DP_mult_97_n205), .CO(DP_mult_97_n200), .S(DP_mult_97_n201) );
  FA_X1 DP_mult_97_U85 ( .A(DP_mult_97_n203), .B(DP_mult_97_n212), .CI(
        DP_mult_97_n210), .CO(DP_mult_97_n198), .S(DP_mult_97_n199) );
  FA_X1 DP_mult_97_U84 ( .A(DP_mult_97_n208), .B(DP_mult_97_n201), .CI(
        DP_mult_97_n199), .CO(DP_mult_97_n196), .S(DP_mult_97_n197) );
  FA_X1 DP_mult_97_U81 ( .A(DP_mult_97_n271), .B(DP_mult_97_n293), .CI(
        DP_mult_97_n327), .CO(DP_mult_97_n192), .S(DP_mult_97_n193) );
  FA_X1 DP_mult_97_U80 ( .A(DP_mult_97_n204), .B(DP_mult_97_n315), .CI(
        DP_mult_97_n195), .CO(DP_mult_97_n190), .S(DP_mult_97_n191) );
  FA_X1 DP_mult_97_U79 ( .A(DP_mult_97_n193), .B(DP_mult_97_n202), .CI(
        DP_mult_97_n200), .CO(DP_mult_97_n188), .S(DP_mult_97_n189) );
  FA_X1 DP_mult_97_U78 ( .A(DP_mult_97_n198), .B(DP_mult_97_n191), .CI(
        DP_mult_97_n189), .CO(DP_mult_97_n186), .S(DP_mult_97_n187) );
  FA_X1 DP_mult_97_U76 ( .A(DP_mult_97_n303), .B(DP_mult_97_n281), .CI(
        DP_mult_97_n185), .CO(DP_mult_97_n182), .S(DP_mult_97_n183) );
  FA_X1 DP_mult_97_U75 ( .A(DP_mult_97_n270), .B(DP_mult_97_n292), .CI(
        DP_mult_97_n194), .CO(DP_mult_97_n180), .S(DP_mult_97_n181) );
  FA_X1 DP_mult_97_U74 ( .A(DP_mult_97_n190), .B(DP_mult_97_n192), .CI(
        DP_mult_97_n183), .CO(DP_mult_97_n178), .S(DP_mult_97_n179) );
  FA_X1 DP_mult_97_U73 ( .A(DP_mult_97_n188), .B(DP_mult_97_n181), .CI(
        DP_mult_97_n179), .CO(DP_mult_97_n176), .S(DP_mult_97_n177) );
  FA_X1 DP_mult_97_U72 ( .A(DP_mult_97_n184), .B(DP_mult_97_n269), .CI(
        DP_mult_97_n314), .CO(DP_mult_97_n174), .S(DP_mult_97_n175) );
  FA_X1 DP_mult_97_U71 ( .A(DP_mult_97_n280), .B(DP_mult_97_n302), .CI(
        DP_mult_97_n291), .CO(DP_mult_97_n172), .S(DP_mult_97_n173) );
  FA_X1 DP_mult_97_U70 ( .A(DP_mult_97_n180), .B(DP_mult_97_n182), .CI(
        DP_mult_97_n173), .CO(DP_mult_97_n170), .S(DP_mult_97_n171) );
  FA_X1 DP_mult_97_U69 ( .A(DP_mult_97_n178), .B(DP_mult_97_n175), .CI(
        DP_mult_97_n171), .CO(DP_mult_97_n168), .S(DP_mult_97_n169) );
  FA_X1 DP_mult_97_U67 ( .A(DP_mult_97_n268), .B(DP_mult_97_n279), .CI(
        DP_mult_97_n167), .CO(DP_mult_97_n164), .S(DP_mult_97_n165) );
  FA_X1 DP_mult_97_U66 ( .A(DP_mult_97_n174), .B(DP_mult_97_n290), .CI(
        DP_mult_97_n172), .CO(DP_mult_97_n162), .S(DP_mult_97_n163) );
  FA_X1 DP_mult_97_U65 ( .A(DP_mult_97_n170), .B(DP_mult_97_n165), .CI(
        DP_mult_97_n163), .CO(DP_mult_97_n160), .S(DP_mult_97_n161) );
  FA_X1 DP_mult_97_U64 ( .A(DP_mult_97_n166), .B(DP_mult_97_n267), .CI(
        DP_mult_97_n301), .CO(DP_mult_97_n158), .S(DP_mult_97_n159) );
  FA_X1 DP_mult_97_U63 ( .A(DP_mult_97_n278), .B(DP_mult_97_n289), .CI(
        DP_mult_97_n164), .CO(DP_mult_97_n156), .S(DP_mult_97_n157) );
  FA_X1 DP_mult_97_U62 ( .A(DP_mult_97_n162), .B(DP_mult_97_n159), .CI(
        DP_mult_97_n157), .CO(DP_mult_97_n154), .S(DP_mult_97_n155) );
  FA_X1 DP_mult_97_U60 ( .A(DP_mult_97_n266), .B(DP_mult_97_n277), .CI(
        DP_mult_97_n153), .CO(DP_mult_97_n150), .S(DP_mult_97_n151) );
  FA_X1 DP_mult_97_U59 ( .A(DP_mult_97_n151), .B(DP_mult_97_n158), .CI(
        DP_mult_97_n156), .CO(DP_mult_97_n148), .S(DP_mult_97_n149) );
  FA_X1 DP_mult_97_U58 ( .A(DP_mult_97_n265), .B(DP_mult_97_n152), .CI(
        DP_mult_97_n288), .CO(DP_mult_97_n146), .S(DP_mult_97_n147) );
  FA_X1 DP_mult_97_U57 ( .A(DP_mult_97_n150), .B(DP_mult_97_n276), .CI(
        DP_mult_97_n147), .CO(DP_mult_97_n144), .S(DP_mult_97_n145) );
  FA_X1 DP_mult_97_U55 ( .A(DP_mult_97_n143), .B(DP_mult_97_n264), .CI(
        DP_mult_97_n146), .CO(DP_mult_97_n140), .S(DP_mult_97_n141) );
  FA_X1 DP_mult_97_U54 ( .A(DP_mult_97_n263), .B(DP_mult_97_n142), .CI(
        DP_mult_97_n275), .CO(DP_mult_97_n138), .S(DP_mult_97_n139) );
  FA_X1 DP_mult_97_U42 ( .A(DP_mult_97_n207), .B(DP_mult_97_n216), .CI(
        DP_mult_97_n126), .CO(DP_mult_97_n125), .S(DP_sw1_a2_0_) );
  FA_X1 DP_mult_97_U41 ( .A(DP_mult_97_n197), .B(DP_mult_97_n206), .CI(
        DP_mult_97_n125), .CO(DP_mult_97_n124), .S(DP_sw1_a2_1_) );
  FA_X1 DP_mult_97_U40 ( .A(DP_mult_97_n187), .B(DP_mult_97_n196), .CI(
        DP_mult_97_n124), .CO(DP_mult_97_n123), .S(DP_sw1_a2_2_) );
  FA_X1 DP_mult_97_U39 ( .A(DP_mult_97_n177), .B(DP_mult_97_n186), .CI(
        DP_mult_97_n123), .CO(DP_mult_97_n122), .S(DP_sw1_a2_3_) );
  FA_X1 DP_mult_97_U38 ( .A(DP_mult_97_n169), .B(DP_mult_97_n176), .CI(
        DP_mult_97_n122), .CO(DP_mult_97_n121), .S(DP_sw1_a2_4_) );
  FA_X1 DP_mult_97_U37 ( .A(DP_mult_97_n161), .B(DP_mult_97_n168), .CI(
        DP_mult_97_n121), .CO(DP_mult_97_n120), .S(DP_sw1_a2_5_) );
  FA_X1 DP_mult_97_U36 ( .A(DP_mult_97_n155), .B(DP_mult_97_n160), .CI(
        DP_mult_97_n120), .CO(DP_mult_97_n119), .S(DP_sw1_a2_6_) );
  FA_X1 DP_mult_97_U30 ( .A(DP_mult_97_n149), .B(DP_mult_97_n154), .CI(
        DP_mult_97_n119), .CO(DP_mult_97_n118), .S(DP_sw1_a2_7_) );
  FA_X1 DP_mult_97_U20 ( .A(DP_mult_97_n145), .B(DP_mult_97_n148), .CI(
        DP_mult_97_n118), .CO(DP_mult_97_n117), .S(DP_sw1_a2_8_) );
  FA_X1 DP_mult_97_U10 ( .A(DP_mult_97_n141), .B(DP_mult_97_n144), .CI(
        DP_mult_97_n117), .CO(DP_mult_97_n116), .S(DP_sw1_a2_9_) );
  FA_X1 DP_mult_97_U9 ( .A(DP_mult_97_n140), .B(DP_mult_97_n139), .CI(
        DP_mult_97_n116), .CO(DP_mult_97_n115), .S(DP_sw1_a2_10_) );
  XOR2_X1 DP_mult_99_U563 ( .A(DP_b_int[33]), .B(DP_b_int[34]), .Z(
        DP_mult_99_n653) );
  INV_X1 DP_mult_99_U562 ( .A(DP_b_int[34]), .ZN(DP_mult_99_n543) );
  NOR2_X1 DP_mult_99_U561 ( .A1(DP_mult_99_n543), .A2(DP_sw1_1_), .ZN(
        DP_mult_99_n658) );
  INV_X1 DP_mult_99_U560 ( .A(DP_mult_99_n658), .ZN(DP_mult_99_n660) );
  NAND2_X1 DP_mult_99_U559 ( .A1(DP_b_int[34]), .A2(DP_mult_99_n532), .ZN(
        DP_mult_99_n530) );
  XNOR2_X1 DP_mult_99_U558 ( .A(DP_sw1_2_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n529) );
  OAI22_X1 DP_mult_99_U557 ( .A1(DP_mult_99_n660), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n529), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n659) );
  NAND2_X1 DP_mult_99_U556 ( .A1(DP_mult_99_n653), .A2(DP_mult_99_n659), .ZN(
        DP_mult_99_n656) );
  NAND2_X1 DP_mult_99_U555 ( .A1(DP_mult_99_n658), .A2(DP_mult_99_n659), .ZN(
        DP_mult_99_n657) );
  INV_X1 DP_mult_99_U554 ( .A(DP_sw1_0_), .ZN(DP_mult_99_n560) );
  MUX2_X1 DP_mult_99_U553 ( .A(DP_mult_99_n656), .B(DP_mult_99_n657), .S(
        DP_mult_99_n560), .Z(DP_mult_99_n655) );
  INV_X1 DP_mult_99_U552 ( .A(DP_mult_99_n655), .ZN(DP_mult_99_n650) );
  INV_X1 DP_mult_99_U551 ( .A(DP_b_int[32]), .ZN(DP_mult_99_n632) );
  XNOR2_X1 DP_mult_99_U550 ( .A(DP_mult_99_n632), .B(DP_b_int[33]), .ZN(
        DP_mult_99_n654) );
  NAND2_X1 DP_mult_99_U549 ( .A1(DP_mult_99_n546), .A2(DP_mult_99_n654), .ZN(
        DP_mult_99_n545) );
  NAND3_X1 DP_mult_99_U548 ( .A1(DP_mult_99_n653), .A2(DP_mult_99_n560), .A3(
        DP_b_int[32]), .ZN(DP_mult_99_n652) );
  OAI21_X1 DP_mult_99_U547 ( .B1(DP_mult_99_n632), .B2(DP_mult_99_n545), .A(
        DP_mult_99_n652), .ZN(DP_mult_99_n651) );
  AOI222_X1 DP_mult_99_U546 ( .A1(DP_mult_99_n650), .A2(DP_mult_99_n255), .B1(
        DP_mult_99_n651), .B2(DP_mult_99_n650), .C1(DP_mult_99_n651), .C2(
        DP_mult_99_n255), .ZN(DP_mult_99_n649) );
  INV_X1 DP_mult_99_U545 ( .A(DP_mult_99_n649), .ZN(DP_mult_99_n648) );
  AOI222_X1 DP_mult_99_U544 ( .A1(DP_mult_99_n648), .A2(DP_mult_99_n253), .B1(
        DP_mult_99_n648), .B2(DP_mult_99_n254), .C1(DP_mult_99_n254), .C2(
        DP_mult_99_n253), .ZN(DP_mult_99_n647) );
  INV_X1 DP_mult_99_U543 ( .A(DP_mult_99_n647), .ZN(DP_mult_99_n646) );
  AOI222_X1 DP_mult_99_U542 ( .A1(DP_mult_99_n646), .A2(DP_mult_99_n249), .B1(
        DP_mult_99_n646), .B2(DP_mult_99_n252), .C1(DP_mult_99_n252), .C2(
        DP_mult_99_n249), .ZN(DP_mult_99_n645) );
  INV_X1 DP_mult_99_U541 ( .A(DP_mult_99_n645), .ZN(DP_mult_99_n644) );
  AOI222_X1 DP_mult_99_U540 ( .A1(DP_mult_99_n644), .A2(DP_mult_99_n245), .B1(
        DP_mult_99_n644), .B2(DP_mult_99_n248), .C1(DP_mult_99_n248), .C2(
        DP_mult_99_n245), .ZN(DP_mult_99_n643) );
  INV_X1 DP_mult_99_U539 ( .A(DP_mult_99_n643), .ZN(DP_mult_99_n642) );
  AOI222_X1 DP_mult_99_U538 ( .A1(DP_mult_99_n642), .A2(DP_mult_99_n239), .B1(
        DP_mult_99_n642), .B2(DP_mult_99_n244), .C1(DP_mult_99_n244), .C2(
        DP_mult_99_n239), .ZN(DP_mult_99_n639) );
  INV_X1 DP_mult_99_U537 ( .A(DP_mult_99_n233), .ZN(DP_mult_99_n640) );
  INV_X1 DP_mult_99_U536 ( .A(DP_mult_99_n238), .ZN(DP_mult_99_n641) );
  OAI222_X1 DP_mult_99_U535 ( .A1(DP_mult_99_n639), .A2(DP_mult_99_n640), .B1(
        DP_mult_99_n639), .B2(DP_mult_99_n641), .C1(DP_mult_99_n641), .C2(
        DP_mult_99_n640), .ZN(DP_mult_99_n638) );
  AOI222_X1 DP_mult_99_U534 ( .A1(DP_mult_99_n638), .A2(DP_mult_99_n225), .B1(
        DP_mult_99_n638), .B2(DP_mult_99_n232), .C1(DP_mult_99_n232), .C2(
        DP_mult_99_n225), .ZN(DP_mult_99_n635) );
  INV_X1 DP_mult_99_U533 ( .A(DP_mult_99_n217), .ZN(DP_mult_99_n636) );
  INV_X1 DP_mult_99_U532 ( .A(DP_mult_99_n224), .ZN(DP_mult_99_n637) );
  OAI222_X1 DP_mult_99_U531 ( .A1(DP_mult_99_n635), .A2(DP_mult_99_n636), .B1(
        DP_mult_99_n635), .B2(DP_mult_99_n637), .C1(DP_mult_99_n637), .C2(
        DP_mult_99_n636), .ZN(DP_mult_99_n126) );
  XNOR2_X1 DP_mult_99_U530 ( .A(DP_sw1_11_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n606) );
  INV_X1 DP_mult_99_U529 ( .A(DP_b_int[28]), .ZN(DP_mult_99_n622) );
  INV_X1 DP_mult_99_U528 ( .A(DP_b_int[26]), .ZN(DP_mult_99_n624) );
  XNOR2_X1 DP_mult_99_U527 ( .A(DP_mult_99_n624), .B(DP_b_int[27]), .ZN(
        DP_mult_99_n634) );
  NAND2_X1 DP_mult_99_U526 ( .A1(DP_mult_99_n593), .A2(DP_mult_99_n634), .ZN(
        DP_mult_99_n595) );
  XNOR2_X1 DP_mult_99_U525 ( .A(DP_sw1_12_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n608) );
  OAI22_X1 DP_mult_99_U524 ( .A1(DP_mult_99_n606), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n608), .ZN(DP_mult_99_n142) );
  INV_X1 DP_mult_99_U523 ( .A(DP_mult_99_n142), .ZN(DP_mult_99_n143) );
  XNOR2_X1 DP_mult_99_U522 ( .A(DP_sw1_11_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n590) );
  INV_X1 DP_mult_99_U521 ( .A(DP_b_int[30]), .ZN(DP_mult_99_n620) );
  XNOR2_X1 DP_mult_99_U520 ( .A(DP_mult_99_n622), .B(DP_b_int[29]), .ZN(
        DP_mult_99_n633) );
  NAND2_X1 DP_mult_99_U519 ( .A1(DP_mult_99_n577), .A2(DP_mult_99_n633), .ZN(
        DP_mult_99_n579) );
  XNOR2_X1 DP_mult_99_U518 ( .A(DP_sw1_12_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n592) );
  OAI22_X1 DP_mult_99_U517 ( .A1(DP_mult_99_n590), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n592), .ZN(DP_mult_99_n152) );
  INV_X1 DP_mult_99_U516 ( .A(DP_mult_99_n152), .ZN(DP_mult_99_n153) );
  XNOR2_X1 DP_mult_99_U515 ( .A(DP_sw1_11_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n574) );
  XNOR2_X1 DP_mult_99_U514 ( .A(DP_mult_99_n620), .B(DP_b_int[31]), .ZN(
        DP_mult_99_n631) );
  NAND2_X1 DP_mult_99_U513 ( .A1(DP_mult_99_n561), .A2(DP_mult_99_n631), .ZN(
        DP_mult_99_n563) );
  XNOR2_X1 DP_mult_99_U512 ( .A(DP_sw1_12_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n576) );
  OAI22_X1 DP_mult_99_U511 ( .A1(DP_mult_99_n574), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n576), .ZN(DP_mult_99_n166) );
  INV_X1 DP_mult_99_U510 ( .A(DP_mult_99_n166), .ZN(DP_mult_99_n167) );
  XNOR2_X1 DP_mult_99_U509 ( .A(DP_sw1_11_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n557) );
  XNOR2_X1 DP_mult_99_U508 ( .A(DP_sw1_12_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n559) );
  OAI22_X1 DP_mult_99_U507 ( .A1(DP_mult_99_n557), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n559), .ZN(DP_mult_99_n184) );
  INV_X1 DP_mult_99_U506 ( .A(DP_mult_99_n184), .ZN(DP_mult_99_n185) );
  XNOR2_X1 DP_mult_99_U505 ( .A(DP_sw1_4_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n599) );
  XNOR2_X1 DP_mult_99_U504 ( .A(DP_sw1_5_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n600) );
  OAI22_X1 DP_mult_99_U503 ( .A1(DP_mult_99_n599), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n600), .ZN(DP_mult_99_n629) );
  XNOR2_X1 DP_mult_99_U502 ( .A(DP_sw1_8_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n571) );
  XNOR2_X1 DP_mult_99_U501 ( .A(DP_sw1_9_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n572) );
  OAI22_X1 DP_mult_99_U500 ( .A1(DP_mult_99_n571), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n572), .ZN(DP_mult_99_n630) );
  OR2_X1 DP_mult_99_U499 ( .A1(DP_mult_99_n629), .A2(DP_mult_99_n630), .ZN(
        DP_mult_99_n194) );
  XNOR2_X1 DP_mult_99_U498 ( .A(DP_mult_99_n629), .B(DP_mult_99_n630), .ZN(
        DP_mult_99_n195) );
  INV_X1 DP_mult_99_U497 ( .A(DP_b_int[24]), .ZN(DP_mult_99_n626) );
  XNOR2_X1 DP_mult_99_U496 ( .A(DP_mult_99_n626), .B(DP_b_int[25]), .ZN(
        DP_mult_99_n628) );
  NAND2_X1 DP_mult_99_U495 ( .A1(DP_mult_99_n526), .A2(DP_mult_99_n628), .ZN(
        DP_mult_99_n525) );
  OR3_X1 DP_mult_99_U494 ( .A1(DP_mult_99_n526), .A2(DP_sw1_0_), .A3(
        DP_mult_99_n626), .ZN(DP_mult_99_n627) );
  OAI21_X1 DP_mult_99_U493 ( .B1(DP_mult_99_n626), .B2(DP_mult_99_n525), .A(
        DP_mult_99_n627), .ZN(DP_mult_99_n256) );
  OR3_X1 DP_mult_99_U492 ( .A1(DP_mult_99_n593), .A2(DP_sw1_0_), .A3(
        DP_mult_99_n624), .ZN(DP_mult_99_n625) );
  OAI21_X1 DP_mult_99_U491 ( .B1(DP_mult_99_n624), .B2(DP_mult_99_n595), .A(
        DP_mult_99_n625), .ZN(DP_mult_99_n257) );
  OR3_X1 DP_mult_99_U490 ( .A1(DP_mult_99_n577), .A2(DP_sw1_0_), .A3(
        DP_mult_99_n622), .ZN(DP_mult_99_n623) );
  OAI21_X1 DP_mult_99_U489 ( .B1(DP_mult_99_n622), .B2(DP_mult_99_n579), .A(
        DP_mult_99_n623), .ZN(DP_mult_99_n258) );
  OR3_X1 DP_mult_99_U488 ( .A1(DP_mult_99_n561), .A2(DP_sw1_0_), .A3(
        DP_mult_99_n620), .ZN(DP_mult_99_n621) );
  OAI21_X1 DP_mult_99_U487 ( .B1(DP_mult_99_n620), .B2(DP_mult_99_n563), .A(
        DP_mult_99_n621), .ZN(DP_mult_99_n259) );
  XNOR2_X1 DP_mult_99_U486 ( .A(DP_sw1_10_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n619) );
  XNOR2_X1 DP_mult_99_U485 ( .A(DP_sw1_11_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n528) );
  OAI22_X1 DP_mult_99_U484 ( .A1(DP_mult_99_n619), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n528), .ZN(DP_mult_99_n263) );
  XNOR2_X1 DP_mult_99_U483 ( .A(DP_sw1_9_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n618) );
  OAI22_X1 DP_mult_99_U482 ( .A1(DP_mult_99_n618), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n619), .ZN(DP_mult_99_n264) );
  XNOR2_X1 DP_mult_99_U481 ( .A(DP_sw1_8_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n617) );
  OAI22_X1 DP_mult_99_U480 ( .A1(DP_mult_99_n617), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n618), .ZN(DP_mult_99_n265) );
  XNOR2_X1 DP_mult_99_U479 ( .A(DP_sw1_7_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n616) );
  OAI22_X1 DP_mult_99_U478 ( .A1(DP_mult_99_n616), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n617), .ZN(DP_mult_99_n266) );
  XNOR2_X1 DP_mult_99_U477 ( .A(DP_sw1_6_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n615) );
  OAI22_X1 DP_mult_99_U476 ( .A1(DP_mult_99_n615), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n616), .ZN(DP_mult_99_n267) );
  XNOR2_X1 DP_mult_99_U475 ( .A(DP_sw1_5_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n614) );
  OAI22_X1 DP_mult_99_U474 ( .A1(DP_mult_99_n614), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n615), .ZN(DP_mult_99_n268) );
  XNOR2_X1 DP_mult_99_U473 ( .A(DP_sw1_4_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n613) );
  OAI22_X1 DP_mult_99_U472 ( .A1(DP_mult_99_n613), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n614), .ZN(DP_mult_99_n269) );
  XNOR2_X1 DP_mult_99_U471 ( .A(DP_sw1_3_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n612) );
  OAI22_X1 DP_mult_99_U470 ( .A1(DP_mult_99_n612), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n613), .ZN(DP_mult_99_n270) );
  XNOR2_X1 DP_mult_99_U469 ( .A(DP_sw1_2_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n611) );
  OAI22_X1 DP_mult_99_U468 ( .A1(DP_mult_99_n611), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n612), .ZN(DP_mult_99_n271) );
  XNOR2_X1 DP_mult_99_U467 ( .A(DP_sw1_1_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n610) );
  OAI22_X1 DP_mult_99_U466 ( .A1(DP_mult_99_n610), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n611), .ZN(DP_mult_99_n272) );
  XNOR2_X1 DP_mult_99_U465 ( .A(DP_sw1_0_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n609) );
  OAI22_X1 DP_mult_99_U464 ( .A1(DP_mult_99_n609), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n610), .ZN(DP_mult_99_n273) );
  NOR2_X1 DP_mult_99_U463 ( .A1(DP_mult_99_n560), .A2(DP_mult_99_n526), .ZN(
        DP_mult_99_n274) );
  AOI21_X1 DP_mult_99_U462 ( .B1(DP_mult_99_n595), .B2(DP_mult_99_n593), .A(
        DP_mult_99_n608), .ZN(DP_mult_99_n607) );
  INV_X1 DP_mult_99_U461 ( .A(DP_mult_99_n607), .ZN(DP_mult_99_n275) );
  XNOR2_X1 DP_mult_99_U460 ( .A(DP_sw1_10_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n605) );
  OAI22_X1 DP_mult_99_U459 ( .A1(DP_mult_99_n605), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n606), .ZN(DP_mult_99_n276) );
  XNOR2_X1 DP_mult_99_U458 ( .A(DP_sw1_9_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n604) );
  OAI22_X1 DP_mult_99_U457 ( .A1(DP_mult_99_n604), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n605), .ZN(DP_mult_99_n277) );
  XNOR2_X1 DP_mult_99_U456 ( .A(DP_sw1_8_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n603) );
  OAI22_X1 DP_mult_99_U455 ( .A1(DP_mult_99_n603), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n604), .ZN(DP_mult_99_n278) );
  XNOR2_X1 DP_mult_99_U454 ( .A(DP_sw1_7_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n602) );
  OAI22_X1 DP_mult_99_U453 ( .A1(DP_mult_99_n602), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n603), .ZN(DP_mult_99_n279) );
  XNOR2_X1 DP_mult_99_U452 ( .A(DP_sw1_6_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n601) );
  OAI22_X1 DP_mult_99_U451 ( .A1(DP_mult_99_n601), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n602), .ZN(DP_mult_99_n280) );
  OAI22_X1 DP_mult_99_U450 ( .A1(DP_mult_99_n600), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n601), .ZN(DP_mult_99_n281) );
  XNOR2_X1 DP_mult_99_U449 ( .A(DP_sw1_3_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n598) );
  OAI22_X1 DP_mult_99_U448 ( .A1(DP_mult_99_n598), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n599), .ZN(DP_mult_99_n283) );
  XNOR2_X1 DP_mult_99_U447 ( .A(DP_sw1_2_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n597) );
  OAI22_X1 DP_mult_99_U446 ( .A1(DP_mult_99_n597), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n598), .ZN(DP_mult_99_n284) );
  XNOR2_X1 DP_mult_99_U445 ( .A(DP_sw1_1_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n596) );
  OAI22_X1 DP_mult_99_U444 ( .A1(DP_mult_99_n596), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n597), .ZN(DP_mult_99_n285) );
  XNOR2_X1 DP_mult_99_U443 ( .A(DP_sw1_0_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n594) );
  OAI22_X1 DP_mult_99_U442 ( .A1(DP_mult_99_n594), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n596), .ZN(DP_mult_99_n286) );
  NOR2_X1 DP_mult_99_U441 ( .A1(DP_mult_99_n560), .A2(DP_mult_99_n593), .ZN(
        DP_mult_99_n287) );
  AOI21_X1 DP_mult_99_U440 ( .B1(DP_mult_99_n579), .B2(DP_mult_99_n577), .A(
        DP_mult_99_n592), .ZN(DP_mult_99_n591) );
  INV_X1 DP_mult_99_U439 ( .A(DP_mult_99_n591), .ZN(DP_mult_99_n288) );
  XNOR2_X1 DP_mult_99_U438 ( .A(DP_sw1_10_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n589) );
  OAI22_X1 DP_mult_99_U437 ( .A1(DP_mult_99_n589), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n590), .ZN(DP_mult_99_n289) );
  XNOR2_X1 DP_mult_99_U436 ( .A(DP_sw1_9_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n588) );
  OAI22_X1 DP_mult_99_U435 ( .A1(DP_mult_99_n588), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n589), .ZN(DP_mult_99_n290) );
  XNOR2_X1 DP_mult_99_U434 ( .A(DP_sw1_8_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n587) );
  OAI22_X1 DP_mult_99_U433 ( .A1(DP_mult_99_n587), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n588), .ZN(DP_mult_99_n291) );
  XNOR2_X1 DP_mult_99_U432 ( .A(DP_sw1_7_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n586) );
  OAI22_X1 DP_mult_99_U431 ( .A1(DP_mult_99_n586), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n587), .ZN(DP_mult_99_n292) );
  XNOR2_X1 DP_mult_99_U430 ( .A(DP_sw1_6_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n585) );
  OAI22_X1 DP_mult_99_U429 ( .A1(DP_mult_99_n585), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n586), .ZN(DP_mult_99_n293) );
  XNOR2_X1 DP_mult_99_U428 ( .A(DP_sw1_5_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n584) );
  OAI22_X1 DP_mult_99_U427 ( .A1(DP_mult_99_n584), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n585), .ZN(DP_mult_99_n294) );
  XNOR2_X1 DP_mult_99_U426 ( .A(DP_sw1_4_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n583) );
  OAI22_X1 DP_mult_99_U425 ( .A1(DP_mult_99_n583), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n584), .ZN(DP_mult_99_n295) );
  XNOR2_X1 DP_mult_99_U424 ( .A(DP_sw1_3_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n582) );
  OAI22_X1 DP_mult_99_U423 ( .A1(DP_mult_99_n582), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n583), .ZN(DP_mult_99_n296) );
  XNOR2_X1 DP_mult_99_U422 ( .A(DP_sw1_2_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n581) );
  OAI22_X1 DP_mult_99_U421 ( .A1(DP_mult_99_n581), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n582), .ZN(DP_mult_99_n297) );
  XNOR2_X1 DP_mult_99_U420 ( .A(DP_sw1_1_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n580) );
  OAI22_X1 DP_mult_99_U419 ( .A1(DP_mult_99_n580), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n581), .ZN(DP_mult_99_n298) );
  XNOR2_X1 DP_mult_99_U418 ( .A(DP_sw1_0_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n578) );
  OAI22_X1 DP_mult_99_U417 ( .A1(DP_mult_99_n578), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n580), .ZN(DP_mult_99_n299) );
  NOR2_X1 DP_mult_99_U416 ( .A1(DP_mult_99_n560), .A2(DP_mult_99_n577), .ZN(
        DP_mult_99_n300) );
  AOI21_X1 DP_mult_99_U415 ( .B1(DP_mult_99_n563), .B2(DP_mult_99_n561), .A(
        DP_mult_99_n576), .ZN(DP_mult_99_n575) );
  INV_X1 DP_mult_99_U414 ( .A(DP_mult_99_n575), .ZN(DP_mult_99_n301) );
  XNOR2_X1 DP_mult_99_U413 ( .A(DP_sw1_10_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n573) );
  OAI22_X1 DP_mult_99_U412 ( .A1(DP_mult_99_n573), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n574), .ZN(DP_mult_99_n302) );
  OAI22_X1 DP_mult_99_U411 ( .A1(DP_mult_99_n572), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n573), .ZN(DP_mult_99_n303) );
  XNOR2_X1 DP_mult_99_U410 ( .A(DP_sw1_7_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n570) );
  OAI22_X1 DP_mult_99_U409 ( .A1(DP_mult_99_n570), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n571), .ZN(DP_mult_99_n305) );
  XNOR2_X1 DP_mult_99_U408 ( .A(DP_sw1_6_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n569) );
  OAI22_X1 DP_mult_99_U407 ( .A1(DP_mult_99_n569), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n570), .ZN(DP_mult_99_n306) );
  XNOR2_X1 DP_mult_99_U406 ( .A(DP_sw1_5_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n568) );
  OAI22_X1 DP_mult_99_U405 ( .A1(DP_mult_99_n568), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n569), .ZN(DP_mult_99_n307) );
  XNOR2_X1 DP_mult_99_U404 ( .A(DP_sw1_4_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n567) );
  OAI22_X1 DP_mult_99_U403 ( .A1(DP_mult_99_n567), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n568), .ZN(DP_mult_99_n308) );
  XNOR2_X1 DP_mult_99_U402 ( .A(DP_sw1_3_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n566) );
  OAI22_X1 DP_mult_99_U401 ( .A1(DP_mult_99_n566), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n567), .ZN(DP_mult_99_n309) );
  XNOR2_X1 DP_mult_99_U400 ( .A(DP_sw1_2_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n565) );
  OAI22_X1 DP_mult_99_U399 ( .A1(DP_mult_99_n565), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n566), .ZN(DP_mult_99_n310) );
  XNOR2_X1 DP_mult_99_U398 ( .A(DP_sw1_1_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n564) );
  OAI22_X1 DP_mult_99_U397 ( .A1(DP_mult_99_n564), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n565), .ZN(DP_mult_99_n311) );
  XNOR2_X1 DP_mult_99_U396 ( .A(DP_sw1_0_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n562) );
  OAI22_X1 DP_mult_99_U395 ( .A1(DP_mult_99_n562), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n564), .ZN(DP_mult_99_n312) );
  NOR2_X1 DP_mult_99_U394 ( .A1(DP_mult_99_n560), .A2(DP_mult_99_n561), .ZN(
        DP_mult_99_n313) );
  AOI21_X1 DP_mult_99_U393 ( .B1(DP_mult_99_n545), .B2(DP_mult_99_n546), .A(
        DP_mult_99_n559), .ZN(DP_mult_99_n558) );
  INV_X1 DP_mult_99_U392 ( .A(DP_mult_99_n558), .ZN(DP_mult_99_n314) );
  XNOR2_X1 DP_mult_99_U391 ( .A(DP_sw1_10_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n556) );
  OAI22_X1 DP_mult_99_U390 ( .A1(DP_mult_99_n556), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n557), .ZN(DP_mult_99_n315) );
  XNOR2_X1 DP_mult_99_U389 ( .A(DP_sw1_9_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n555) );
  OAI22_X1 DP_mult_99_U388 ( .A1(DP_mult_99_n555), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n556), .ZN(DP_mult_99_n316) );
  XNOR2_X1 DP_mult_99_U387 ( .A(DP_sw1_8_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n554) );
  OAI22_X1 DP_mult_99_U386 ( .A1(DP_mult_99_n554), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n555), .ZN(DP_mult_99_n317) );
  XNOR2_X1 DP_mult_99_U385 ( .A(DP_sw1_7_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n553) );
  OAI22_X1 DP_mult_99_U384 ( .A1(DP_mult_99_n553), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n554), .ZN(DP_mult_99_n318) );
  XNOR2_X1 DP_mult_99_U383 ( .A(DP_sw1_6_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n552) );
  OAI22_X1 DP_mult_99_U382 ( .A1(DP_mult_99_n552), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n553), .ZN(DP_mult_99_n319) );
  XNOR2_X1 DP_mult_99_U381 ( .A(DP_sw1_5_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n551) );
  OAI22_X1 DP_mult_99_U380 ( .A1(DP_mult_99_n551), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n552), .ZN(DP_mult_99_n320) );
  XNOR2_X1 DP_mult_99_U379 ( .A(DP_sw1_4_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n550) );
  OAI22_X1 DP_mult_99_U378 ( .A1(DP_mult_99_n550), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n551), .ZN(DP_mult_99_n321) );
  XNOR2_X1 DP_mult_99_U377 ( .A(DP_sw1_3_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n549) );
  OAI22_X1 DP_mult_99_U376 ( .A1(DP_mult_99_n549), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n550), .ZN(DP_mult_99_n322) );
  XNOR2_X1 DP_mult_99_U375 ( .A(DP_sw1_2_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n548) );
  OAI22_X1 DP_mult_99_U374 ( .A1(DP_mult_99_n548), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n549), .ZN(DP_mult_99_n323) );
  XNOR2_X1 DP_mult_99_U373 ( .A(DP_sw1_1_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n547) );
  OAI22_X1 DP_mult_99_U372 ( .A1(DP_mult_99_n547), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n548), .ZN(DP_mult_99_n324) );
  XNOR2_X1 DP_mult_99_U371 ( .A(DP_sw1_0_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n544) );
  OAI22_X1 DP_mult_99_U370 ( .A1(DP_mult_99_n544), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n547), .ZN(DP_mult_99_n325) );
  XOR2_X1 DP_mult_99_U369 ( .A(DP_sw1_12_), .B(DP_mult_99_n543), .Z(
        DP_mult_99_n541) );
  AOI21_X1 DP_mult_99_U368 ( .B1(DP_mult_99_n530), .B2(DP_mult_99_n532), .A(
        DP_mult_99_n541), .ZN(DP_mult_99_n542) );
  INV_X1 DP_mult_99_U367 ( .A(DP_mult_99_n542), .ZN(DP_mult_99_n327) );
  XNOR2_X1 DP_mult_99_U366 ( .A(DP_sw1_11_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n540) );
  OAI22_X1 DP_mult_99_U365 ( .A1(DP_mult_99_n540), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n541), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n328) );
  XNOR2_X1 DP_mult_99_U364 ( .A(DP_sw1_10_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n539) );
  OAI22_X1 DP_mult_99_U363 ( .A1(DP_mult_99_n539), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n540), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n329) );
  XNOR2_X1 DP_mult_99_U362 ( .A(DP_sw1_9_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n538) );
  OAI22_X1 DP_mult_99_U361 ( .A1(DP_mult_99_n538), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n539), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n330) );
  XNOR2_X1 DP_mult_99_U360 ( .A(DP_sw1_8_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n537) );
  OAI22_X1 DP_mult_99_U359 ( .A1(DP_mult_99_n537), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n538), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n331) );
  XNOR2_X1 DP_mult_99_U358 ( .A(DP_sw1_7_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n536) );
  OAI22_X1 DP_mult_99_U357 ( .A1(DP_mult_99_n536), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n537), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n332) );
  XNOR2_X1 DP_mult_99_U356 ( .A(DP_sw1_6_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n535) );
  OAI22_X1 DP_mult_99_U355 ( .A1(DP_mult_99_n535), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n536), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n333) );
  XNOR2_X1 DP_mult_99_U354 ( .A(DP_sw1_5_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n534) );
  OAI22_X1 DP_mult_99_U353 ( .A1(DP_mult_99_n534), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n535), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n334) );
  XNOR2_X1 DP_mult_99_U352 ( .A(DP_sw1_4_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n533) );
  OAI22_X1 DP_mult_99_U351 ( .A1(DP_mult_99_n533), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n534), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n335) );
  XNOR2_X1 DP_mult_99_U350 ( .A(DP_sw1_3_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n531) );
  OAI22_X1 DP_mult_99_U349 ( .A1(DP_mult_99_n531), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n533), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n336) );
  OAI22_X1 DP_mult_99_U348 ( .A1(DP_mult_99_n529), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n531), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n337) );
  XNOR2_X1 DP_mult_99_U347 ( .A(DP_sw1_12_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n527) );
  OAI22_X1 DP_mult_99_U346 ( .A1(DP_mult_99_n528), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n527), .ZN(DP_mult_99_n519) );
  AOI21_X1 DP_mult_99_U345 ( .B1(DP_mult_99_n525), .B2(DP_mult_99_n526), .A(
        DP_mult_99_n527), .ZN(DP_mult_99_n522) );
  INV_X1 DP_mult_99_U344 ( .A(DP_mult_99_n522), .ZN(DP_mult_99_n520) );
  INV_X1 DP_mult_99_U343 ( .A(DP_mult_99_n519), .ZN(DP_mult_99_n524) );
  AOI222_X1 DP_mult_99_U342 ( .A1(DP_mult_99_n115), .A2(DP_mult_99_n138), .B1(
        DP_mult_99_n524), .B2(DP_mult_99_n115), .C1(DP_mult_99_n524), .C2(
        DP_mult_99_n138), .ZN(DP_mult_99_n523) );
  OAI22_X1 DP_mult_99_U341 ( .A1(DP_mult_99_n522), .A2(DP_mult_99_n523), .B1(
        DP_mult_99_n524), .B2(DP_mult_99_n523), .ZN(DP_mult_99_n521) );
  AOI21_X1 DP_mult_99_U340 ( .B1(DP_mult_99_n519), .B2(DP_mult_99_n520), .A(
        DP_mult_99_n521), .ZN(DP_sw1_b2_11_) );
  XOR2_X2 DP_mult_99_U339 ( .A(DP_b_int[27]), .B(DP_mult_99_n622), .Z(
        DP_mult_99_n593) );
  XOR2_X2 DP_mult_99_U338 ( .A(DP_b_int[29]), .B(DP_mult_99_n620), .Z(
        DP_mult_99_n577) );
  XOR2_X2 DP_mult_99_U337 ( .A(DP_b_int[31]), .B(DP_mult_99_n632), .Z(
        DP_mult_99_n561) );
  XOR2_X2 DP_mult_99_U336 ( .A(DP_b_int[25]), .B(DP_mult_99_n624), .Z(
        DP_mult_99_n526) );
  INV_X1 DP_mult_99_U335 ( .A(DP_b_int[35]), .ZN(DP_mult_99_n532) );
  INV_X1 DP_mult_99_U334 ( .A(DP_mult_99_n653), .ZN(DP_mult_99_n546) );
  HA_X1 DP_mult_99_U120 ( .A(DP_mult_99_n325), .B(DP_mult_99_n337), .CO(
        DP_mult_99_n254), .S(DP_mult_99_n255) );
  FA_X1 DP_mult_99_U119 ( .A(DP_mult_99_n336), .B(DP_mult_99_n313), .CI(
        DP_mult_99_n324), .CO(DP_mult_99_n252), .S(DP_mult_99_n253) );
  HA_X1 DP_mult_99_U118 ( .A(DP_mult_99_n259), .B(DP_mult_99_n312), .CO(
        DP_mult_99_n250), .S(DP_mult_99_n251) );
  FA_X1 DP_mult_99_U117 ( .A(DP_mult_99_n323), .B(DP_mult_99_n335), .CI(
        DP_mult_99_n251), .CO(DP_mult_99_n248), .S(DP_mult_99_n249) );
  FA_X1 DP_mult_99_U109 ( .A(DP_mult_99_n334), .B(DP_mult_99_n300), .CI(
        DP_mult_99_n322), .CO(DP_mult_99_n246), .S(DP_mult_99_n247) );
  FA_X1 DP_mult_99_U108 ( .A(DP_mult_99_n250), .B(DP_mult_99_n311), .CI(
        DP_mult_99_n247), .CO(DP_mult_99_n244), .S(DP_mult_99_n245) );
  HA_X1 DP_mult_99_U107 ( .A(DP_mult_99_n258), .B(DP_mult_99_n299), .CO(
        DP_mult_99_n242), .S(DP_mult_99_n243) );
  FA_X1 DP_mult_99_U106 ( .A(DP_mult_99_n310), .B(DP_mult_99_n333), .CI(
        DP_mult_99_n321), .CO(DP_mult_99_n240), .S(DP_mult_99_n241) );
  FA_X1 DP_mult_99_U105 ( .A(DP_mult_99_n246), .B(DP_mult_99_n243), .CI(
        DP_mult_99_n241), .CO(DP_mult_99_n238), .S(DP_mult_99_n239) );
  FA_X1 DP_mult_99_U104 ( .A(DP_mult_99_n309), .B(DP_mult_99_n287), .CI(
        DP_mult_99_n332), .CO(DP_mult_99_n236), .S(DP_mult_99_n237) );
  FA_X1 DP_mult_99_U103 ( .A(DP_mult_99_n298), .B(DP_mult_99_n320), .CI(
        DP_mult_99_n242), .CO(DP_mult_99_n234), .S(DP_mult_99_n235) );
  FA_X1 DP_mult_99_U102 ( .A(DP_mult_99_n237), .B(DP_mult_99_n240), .CI(
        DP_mult_99_n235), .CO(DP_mult_99_n232), .S(DP_mult_99_n233) );
  HA_X1 DP_mult_99_U101 ( .A(DP_mult_99_n257), .B(DP_mult_99_n286), .CO(
        DP_mult_99_n230), .S(DP_mult_99_n231) );
  FA_X1 DP_mult_99_U100 ( .A(DP_mult_99_n297), .B(DP_mult_99_n308), .CI(
        DP_mult_99_n319), .CO(DP_mult_99_n228), .S(DP_mult_99_n229) );
  FA_X1 DP_mult_99_U99 ( .A(DP_mult_99_n231), .B(DP_mult_99_n331), .CI(
        DP_mult_99_n236), .CO(DP_mult_99_n226), .S(DP_mult_99_n227) );
  FA_X1 DP_mult_99_U98 ( .A(DP_mult_99_n229), .B(DP_mult_99_n234), .CI(
        DP_mult_99_n227), .CO(DP_mult_99_n224), .S(DP_mult_99_n225) );
  FA_X1 DP_mult_99_U97 ( .A(DP_mult_99_n296), .B(DP_mult_99_n274), .CI(
        DP_mult_99_n330), .CO(DP_mult_99_n222), .S(DP_mult_99_n223) );
  FA_X1 DP_mult_99_U96 ( .A(DP_mult_99_n285), .B(DP_mult_99_n318), .CI(
        DP_mult_99_n307), .CO(DP_mult_99_n220), .S(DP_mult_99_n221) );
  FA_X1 DP_mult_99_U95 ( .A(DP_mult_99_n228), .B(DP_mult_99_n230), .CI(
        DP_mult_99_n223), .CO(DP_mult_99_n218), .S(DP_mult_99_n219) );
  FA_X1 DP_mult_99_U94 ( .A(DP_mult_99_n226), .B(DP_mult_99_n221), .CI(
        DP_mult_99_n219), .CO(DP_mult_99_n216), .S(DP_mult_99_n217) );
  HA_X1 DP_mult_99_U93 ( .A(DP_mult_99_n256), .B(DP_mult_99_n273), .CO(
        DP_mult_99_n214), .S(DP_mult_99_n215) );
  FA_X1 DP_mult_99_U92 ( .A(DP_mult_99_n284), .B(DP_mult_99_n306), .CI(
        DP_mult_99_n329), .CO(DP_mult_99_n212), .S(DP_mult_99_n213) );
  FA_X1 DP_mult_99_U91 ( .A(DP_mult_99_n295), .B(DP_mult_99_n317), .CI(
        DP_mult_99_n215), .CO(DP_mult_99_n210), .S(DP_mult_99_n211) );
  FA_X1 DP_mult_99_U90 ( .A(DP_mult_99_n220), .B(DP_mult_99_n222), .CI(
        DP_mult_99_n213), .CO(DP_mult_99_n208), .S(DP_mult_99_n209) );
  FA_X1 DP_mult_99_U89 ( .A(DP_mult_99_n218), .B(DP_mult_99_n211), .CI(
        DP_mult_99_n209), .CO(DP_mult_99_n206), .S(DP_mult_99_n207) );
  HA_X1 DP_mult_99_U88 ( .A(DP_mult_99_n272), .B(DP_mult_99_n283), .CO(
        DP_mult_99_n204), .S(DP_mult_99_n205) );
  FA_X1 DP_mult_99_U87 ( .A(DP_mult_99_n328), .B(DP_mult_99_n305), .CI(
        DP_mult_99_n294), .CO(DP_mult_99_n202), .S(DP_mult_99_n203) );
  FA_X1 DP_mult_99_U86 ( .A(DP_mult_99_n214), .B(DP_mult_99_n316), .CI(
        DP_mult_99_n205), .CO(DP_mult_99_n200), .S(DP_mult_99_n201) );
  FA_X1 DP_mult_99_U85 ( .A(DP_mult_99_n203), .B(DP_mult_99_n212), .CI(
        DP_mult_99_n210), .CO(DP_mult_99_n198), .S(DP_mult_99_n199) );
  FA_X1 DP_mult_99_U84 ( .A(DP_mult_99_n208), .B(DP_mult_99_n201), .CI(
        DP_mult_99_n199), .CO(DP_mult_99_n196), .S(DP_mult_99_n197) );
  FA_X1 DP_mult_99_U81 ( .A(DP_mult_99_n271), .B(DP_mult_99_n293), .CI(
        DP_mult_99_n327), .CO(DP_mult_99_n192), .S(DP_mult_99_n193) );
  FA_X1 DP_mult_99_U80 ( .A(DP_mult_99_n204), .B(DP_mult_99_n315), .CI(
        DP_mult_99_n195), .CO(DP_mult_99_n190), .S(DP_mult_99_n191) );
  FA_X1 DP_mult_99_U79 ( .A(DP_mult_99_n193), .B(DP_mult_99_n202), .CI(
        DP_mult_99_n200), .CO(DP_mult_99_n188), .S(DP_mult_99_n189) );
  FA_X1 DP_mult_99_U78 ( .A(DP_mult_99_n198), .B(DP_mult_99_n191), .CI(
        DP_mult_99_n189), .CO(DP_mult_99_n186), .S(DP_mult_99_n187) );
  FA_X1 DP_mult_99_U76 ( .A(DP_mult_99_n303), .B(DP_mult_99_n281), .CI(
        DP_mult_99_n185), .CO(DP_mult_99_n182), .S(DP_mult_99_n183) );
  FA_X1 DP_mult_99_U75 ( .A(DP_mult_99_n270), .B(DP_mult_99_n292), .CI(
        DP_mult_99_n194), .CO(DP_mult_99_n180), .S(DP_mult_99_n181) );
  FA_X1 DP_mult_99_U74 ( .A(DP_mult_99_n190), .B(DP_mult_99_n192), .CI(
        DP_mult_99_n183), .CO(DP_mult_99_n178), .S(DP_mult_99_n179) );
  FA_X1 DP_mult_99_U73 ( .A(DP_mult_99_n188), .B(DP_mult_99_n181), .CI(
        DP_mult_99_n179), .CO(DP_mult_99_n176), .S(DP_mult_99_n177) );
  FA_X1 DP_mult_99_U72 ( .A(DP_mult_99_n184), .B(DP_mult_99_n269), .CI(
        DP_mult_99_n314), .CO(DP_mult_99_n174), .S(DP_mult_99_n175) );
  FA_X1 DP_mult_99_U71 ( .A(DP_mult_99_n280), .B(DP_mult_99_n302), .CI(
        DP_mult_99_n291), .CO(DP_mult_99_n172), .S(DP_mult_99_n173) );
  FA_X1 DP_mult_99_U70 ( .A(DP_mult_99_n180), .B(DP_mult_99_n182), .CI(
        DP_mult_99_n173), .CO(DP_mult_99_n170), .S(DP_mult_99_n171) );
  FA_X1 DP_mult_99_U69 ( .A(DP_mult_99_n178), .B(DP_mult_99_n175), .CI(
        DP_mult_99_n171), .CO(DP_mult_99_n168), .S(DP_mult_99_n169) );
  FA_X1 DP_mult_99_U67 ( .A(DP_mult_99_n268), .B(DP_mult_99_n279), .CI(
        DP_mult_99_n167), .CO(DP_mult_99_n164), .S(DP_mult_99_n165) );
  FA_X1 DP_mult_99_U66 ( .A(DP_mult_99_n174), .B(DP_mult_99_n290), .CI(
        DP_mult_99_n172), .CO(DP_mult_99_n162), .S(DP_mult_99_n163) );
  FA_X1 DP_mult_99_U65 ( .A(DP_mult_99_n170), .B(DP_mult_99_n165), .CI(
        DP_mult_99_n163), .CO(DP_mult_99_n160), .S(DP_mult_99_n161) );
  FA_X1 DP_mult_99_U64 ( .A(DP_mult_99_n166), .B(DP_mult_99_n267), .CI(
        DP_mult_99_n301), .CO(DP_mult_99_n158), .S(DP_mult_99_n159) );
  FA_X1 DP_mult_99_U63 ( .A(DP_mult_99_n278), .B(DP_mult_99_n289), .CI(
        DP_mult_99_n164), .CO(DP_mult_99_n156), .S(DP_mult_99_n157) );
  FA_X1 DP_mult_99_U62 ( .A(DP_mult_99_n162), .B(DP_mult_99_n159), .CI(
        DP_mult_99_n157), .CO(DP_mult_99_n154), .S(DP_mult_99_n155) );
  FA_X1 DP_mult_99_U60 ( .A(DP_mult_99_n266), .B(DP_mult_99_n277), .CI(
        DP_mult_99_n153), .CO(DP_mult_99_n150), .S(DP_mult_99_n151) );
  FA_X1 DP_mult_99_U59 ( .A(DP_mult_99_n151), .B(DP_mult_99_n158), .CI(
        DP_mult_99_n156), .CO(DP_mult_99_n148), .S(DP_mult_99_n149) );
  FA_X1 DP_mult_99_U58 ( .A(DP_mult_99_n265), .B(DP_mult_99_n152), .CI(
        DP_mult_99_n288), .CO(DP_mult_99_n146), .S(DP_mult_99_n147) );
  FA_X1 DP_mult_99_U57 ( .A(DP_mult_99_n150), .B(DP_mult_99_n276), .CI(
        DP_mult_99_n147), .CO(DP_mult_99_n144), .S(DP_mult_99_n145) );
  FA_X1 DP_mult_99_U55 ( .A(DP_mult_99_n143), .B(DP_mult_99_n264), .CI(
        DP_mult_99_n146), .CO(DP_mult_99_n140), .S(DP_mult_99_n141) );
  FA_X1 DP_mult_99_U54 ( .A(DP_mult_99_n263), .B(DP_mult_99_n142), .CI(
        DP_mult_99_n275), .CO(DP_mult_99_n138), .S(DP_mult_99_n139) );
  FA_X1 DP_mult_99_U42 ( .A(DP_mult_99_n207), .B(DP_mult_99_n216), .CI(
        DP_mult_99_n126), .CO(DP_mult_99_n125), .S(DP_sw1_b2_0_) );
  FA_X1 DP_mult_99_U41 ( .A(DP_mult_99_n197), .B(DP_mult_99_n206), .CI(
        DP_mult_99_n125), .CO(DP_mult_99_n124), .S(DP_sw1_b2_1_) );
  FA_X1 DP_mult_99_U40 ( .A(DP_mult_99_n187), .B(DP_mult_99_n196), .CI(
        DP_mult_99_n124), .CO(DP_mult_99_n123), .S(DP_sw1_b2_2_) );
  FA_X1 DP_mult_99_U39 ( .A(DP_mult_99_n177), .B(DP_mult_99_n186), .CI(
        DP_mult_99_n123), .CO(DP_mult_99_n122), .S(DP_sw1_b2_3_) );
  FA_X1 DP_mult_99_U38 ( .A(DP_mult_99_n169), .B(DP_mult_99_n176), .CI(
        DP_mult_99_n122), .CO(DP_mult_99_n121), .S(DP_sw1_b2_4_) );
  FA_X1 DP_mult_99_U37 ( .A(DP_mult_99_n161), .B(DP_mult_99_n168), .CI(
        DP_mult_99_n121), .CO(DP_mult_99_n120), .S(DP_sw1_b2_5_) );
  FA_X1 DP_mult_99_U36 ( .A(DP_mult_99_n155), .B(DP_mult_99_n160), .CI(
        DP_mult_99_n120), .CO(DP_mult_99_n119), .S(DP_sw1_b2_6_) );
  FA_X1 DP_mult_99_U30 ( .A(DP_mult_99_n149), .B(DP_mult_99_n154), .CI(
        DP_mult_99_n119), .CO(DP_mult_99_n118), .S(DP_sw1_b2_7_) );
  FA_X1 DP_mult_99_U20 ( .A(DP_mult_99_n145), .B(DP_mult_99_n148), .CI(
        DP_mult_99_n118), .CO(DP_mult_99_n117), .S(DP_sw1_b2_8_) );
  FA_X1 DP_mult_99_U10 ( .A(DP_mult_99_n141), .B(DP_mult_99_n144), .CI(
        DP_mult_99_n117), .CO(DP_mult_99_n116), .S(DP_sw1_b2_9_) );
  FA_X1 DP_mult_99_U9 ( .A(DP_mult_99_n140), .B(DP_mult_99_n139), .CI(
        DP_mult_99_n116), .CO(DP_mult_99_n115), .S(DP_sw1_b2_10_) );
  XOR2_X1 DP_mult_96_U563 ( .A(DP_a_int[9]), .B(DP_a_int[10]), .Z(
        DP_mult_96_n653) );
  INV_X1 DP_mult_96_U562 ( .A(DP_a_int[10]), .ZN(DP_mult_96_n543) );
  NOR2_X1 DP_mult_96_U561 ( .A1(DP_mult_96_n543), .A2(DP_sw0_1_), .ZN(
        DP_mult_96_n658) );
  INV_X1 DP_mult_96_U560 ( .A(DP_mult_96_n658), .ZN(DP_mult_96_n660) );
  NAND2_X1 DP_mult_96_U559 ( .A1(DP_a_int[10]), .A2(DP_mult_96_n532), .ZN(
        DP_mult_96_n530) );
  XNOR2_X1 DP_mult_96_U558 ( .A(DP_sw0_2_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n529) );
  OAI22_X1 DP_mult_96_U557 ( .A1(DP_mult_96_n660), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n529), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n659) );
  NAND2_X1 DP_mult_96_U556 ( .A1(DP_mult_96_n653), .A2(DP_mult_96_n659), .ZN(
        DP_mult_96_n656) );
  NAND2_X1 DP_mult_96_U555 ( .A1(DP_mult_96_n658), .A2(DP_mult_96_n659), .ZN(
        DP_mult_96_n657) );
  INV_X1 DP_mult_96_U554 ( .A(DP_sw0_0_), .ZN(DP_mult_96_n560) );
  MUX2_X1 DP_mult_96_U553 ( .A(DP_mult_96_n656), .B(DP_mult_96_n657), .S(
        DP_mult_96_n560), .Z(DP_mult_96_n655) );
  INV_X1 DP_mult_96_U552 ( .A(DP_mult_96_n655), .ZN(DP_mult_96_n650) );
  INV_X1 DP_mult_96_U551 ( .A(DP_a_int[8]), .ZN(DP_mult_96_n632) );
  XNOR2_X1 DP_mult_96_U550 ( .A(DP_mult_96_n632), .B(DP_a_int[9]), .ZN(
        DP_mult_96_n654) );
  NAND2_X1 DP_mult_96_U549 ( .A1(DP_mult_96_n546), .A2(DP_mult_96_n654), .ZN(
        DP_mult_96_n545) );
  NAND3_X1 DP_mult_96_U548 ( .A1(DP_mult_96_n653), .A2(DP_mult_96_n560), .A3(
        DP_a_int[8]), .ZN(DP_mult_96_n652) );
  OAI21_X1 DP_mult_96_U547 ( .B1(DP_mult_96_n632), .B2(DP_mult_96_n545), .A(
        DP_mult_96_n652), .ZN(DP_mult_96_n651) );
  AOI222_X1 DP_mult_96_U546 ( .A1(DP_mult_96_n650), .A2(DP_mult_96_n255), .B1(
        DP_mult_96_n651), .B2(DP_mult_96_n650), .C1(DP_mult_96_n651), .C2(
        DP_mult_96_n255), .ZN(DP_mult_96_n649) );
  INV_X1 DP_mult_96_U545 ( .A(DP_mult_96_n649), .ZN(DP_mult_96_n648) );
  AOI222_X1 DP_mult_96_U544 ( .A1(DP_mult_96_n648), .A2(DP_mult_96_n253), .B1(
        DP_mult_96_n648), .B2(DP_mult_96_n254), .C1(DP_mult_96_n254), .C2(
        DP_mult_96_n253), .ZN(DP_mult_96_n647) );
  INV_X1 DP_mult_96_U543 ( .A(DP_mult_96_n647), .ZN(DP_mult_96_n646) );
  AOI222_X1 DP_mult_96_U542 ( .A1(DP_mult_96_n646), .A2(DP_mult_96_n249), .B1(
        DP_mult_96_n646), .B2(DP_mult_96_n252), .C1(DP_mult_96_n252), .C2(
        DP_mult_96_n249), .ZN(DP_mult_96_n645) );
  INV_X1 DP_mult_96_U541 ( .A(DP_mult_96_n645), .ZN(DP_mult_96_n644) );
  AOI222_X1 DP_mult_96_U540 ( .A1(DP_mult_96_n644), .A2(DP_mult_96_n245), .B1(
        DP_mult_96_n644), .B2(DP_mult_96_n248), .C1(DP_mult_96_n248), .C2(
        DP_mult_96_n245), .ZN(DP_mult_96_n643) );
  INV_X1 DP_mult_96_U539 ( .A(DP_mult_96_n643), .ZN(DP_mult_96_n642) );
  AOI222_X1 DP_mult_96_U538 ( .A1(DP_mult_96_n642), .A2(DP_mult_96_n239), .B1(
        DP_mult_96_n642), .B2(DP_mult_96_n244), .C1(DP_mult_96_n244), .C2(
        DP_mult_96_n239), .ZN(DP_mult_96_n639) );
  INV_X1 DP_mult_96_U537 ( .A(DP_mult_96_n233), .ZN(DP_mult_96_n640) );
  INV_X1 DP_mult_96_U536 ( .A(DP_mult_96_n238), .ZN(DP_mult_96_n641) );
  OAI222_X1 DP_mult_96_U535 ( .A1(DP_mult_96_n639), .A2(DP_mult_96_n640), .B1(
        DP_mult_96_n639), .B2(DP_mult_96_n641), .C1(DP_mult_96_n641), .C2(
        DP_mult_96_n640), .ZN(DP_mult_96_n638) );
  AOI222_X1 DP_mult_96_U534 ( .A1(DP_mult_96_n638), .A2(DP_mult_96_n225), .B1(
        DP_mult_96_n638), .B2(DP_mult_96_n232), .C1(DP_mult_96_n232), .C2(
        DP_mult_96_n225), .ZN(DP_mult_96_n635) );
  INV_X1 DP_mult_96_U533 ( .A(DP_mult_96_n217), .ZN(DP_mult_96_n636) );
  INV_X1 DP_mult_96_U532 ( .A(DP_mult_96_n224), .ZN(DP_mult_96_n637) );
  OAI222_X1 DP_mult_96_U531 ( .A1(DP_mult_96_n635), .A2(DP_mult_96_n636), .B1(
        DP_mult_96_n635), .B2(DP_mult_96_n637), .C1(DP_mult_96_n637), .C2(
        DP_mult_96_n636), .ZN(DP_mult_96_n126) );
  XNOR2_X1 DP_mult_96_U530 ( .A(DP_sw0_11_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n606) );
  INV_X1 DP_mult_96_U529 ( .A(DP_a_int[4]), .ZN(DP_mult_96_n622) );
  INV_X1 DP_mult_96_U528 ( .A(DP_a_int[2]), .ZN(DP_mult_96_n624) );
  XNOR2_X1 DP_mult_96_U527 ( .A(DP_mult_96_n624), .B(DP_a_int[3]), .ZN(
        DP_mult_96_n634) );
  NAND2_X1 DP_mult_96_U526 ( .A1(DP_mult_96_n593), .A2(DP_mult_96_n634), .ZN(
        DP_mult_96_n595) );
  XNOR2_X1 DP_mult_96_U525 ( .A(DP_sw0_12_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n608) );
  OAI22_X1 DP_mult_96_U524 ( .A1(DP_mult_96_n606), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n608), .ZN(DP_mult_96_n142) );
  INV_X1 DP_mult_96_U523 ( .A(DP_mult_96_n142), .ZN(DP_mult_96_n143) );
  XNOR2_X1 DP_mult_96_U522 ( .A(DP_sw0_11_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n590) );
  INV_X1 DP_mult_96_U521 ( .A(DP_a_int[6]), .ZN(DP_mult_96_n620) );
  XNOR2_X1 DP_mult_96_U520 ( .A(DP_mult_96_n622), .B(DP_a_int[5]), .ZN(
        DP_mult_96_n633) );
  NAND2_X1 DP_mult_96_U519 ( .A1(DP_mult_96_n577), .A2(DP_mult_96_n633), .ZN(
        DP_mult_96_n579) );
  XNOR2_X1 DP_mult_96_U518 ( .A(DP_sw0_12_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n592) );
  OAI22_X1 DP_mult_96_U517 ( .A1(DP_mult_96_n590), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n592), .ZN(DP_mult_96_n152) );
  INV_X1 DP_mult_96_U516 ( .A(DP_mult_96_n152), .ZN(DP_mult_96_n153) );
  XNOR2_X1 DP_mult_96_U515 ( .A(DP_sw0_11_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n574) );
  XNOR2_X1 DP_mult_96_U514 ( .A(DP_mult_96_n620), .B(DP_a_int[7]), .ZN(
        DP_mult_96_n631) );
  NAND2_X1 DP_mult_96_U513 ( .A1(DP_mult_96_n561), .A2(DP_mult_96_n631), .ZN(
        DP_mult_96_n563) );
  XNOR2_X1 DP_mult_96_U512 ( .A(DP_sw0_12_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n576) );
  OAI22_X1 DP_mult_96_U511 ( .A1(DP_mult_96_n574), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n576), .ZN(DP_mult_96_n166) );
  INV_X1 DP_mult_96_U510 ( .A(DP_mult_96_n166), .ZN(DP_mult_96_n167) );
  XNOR2_X1 DP_mult_96_U509 ( .A(DP_sw0_11_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n557) );
  XNOR2_X1 DP_mult_96_U508 ( .A(DP_sw0_12_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n559) );
  OAI22_X1 DP_mult_96_U507 ( .A1(DP_mult_96_n557), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n559), .ZN(DP_mult_96_n184) );
  INV_X1 DP_mult_96_U506 ( .A(DP_mult_96_n184), .ZN(DP_mult_96_n185) );
  XNOR2_X1 DP_mult_96_U505 ( .A(DP_sw0_4_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n599) );
  XNOR2_X1 DP_mult_96_U504 ( .A(DP_sw0_5_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n600) );
  OAI22_X1 DP_mult_96_U503 ( .A1(DP_mult_96_n599), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n600), .ZN(DP_mult_96_n629) );
  XNOR2_X1 DP_mult_96_U502 ( .A(DP_sw0_8_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n571) );
  XNOR2_X1 DP_mult_96_U501 ( .A(DP_sw0_9_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n572) );
  OAI22_X1 DP_mult_96_U500 ( .A1(DP_mult_96_n571), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n572), .ZN(DP_mult_96_n630) );
  OR2_X1 DP_mult_96_U499 ( .A1(DP_mult_96_n629), .A2(DP_mult_96_n630), .ZN(
        DP_mult_96_n194) );
  XNOR2_X1 DP_mult_96_U498 ( .A(DP_mult_96_n629), .B(DP_mult_96_n630), .ZN(
        DP_mult_96_n195) );
  INV_X1 DP_mult_96_U497 ( .A(DP_a_int[0]), .ZN(DP_mult_96_n626) );
  XNOR2_X1 DP_mult_96_U496 ( .A(DP_mult_96_n626), .B(DP_a_int[1]), .ZN(
        DP_mult_96_n628) );
  NAND2_X1 DP_mult_96_U495 ( .A1(DP_mult_96_n526), .A2(DP_mult_96_n628), .ZN(
        DP_mult_96_n525) );
  OR3_X1 DP_mult_96_U494 ( .A1(DP_mult_96_n526), .A2(DP_sw0_0_), .A3(
        DP_mult_96_n626), .ZN(DP_mult_96_n627) );
  OAI21_X1 DP_mult_96_U493 ( .B1(DP_mult_96_n626), .B2(DP_mult_96_n525), .A(
        DP_mult_96_n627), .ZN(DP_mult_96_n256) );
  OR3_X1 DP_mult_96_U492 ( .A1(DP_mult_96_n593), .A2(DP_sw0_0_), .A3(
        DP_mult_96_n624), .ZN(DP_mult_96_n625) );
  OAI21_X1 DP_mult_96_U491 ( .B1(DP_mult_96_n624), .B2(DP_mult_96_n595), .A(
        DP_mult_96_n625), .ZN(DP_mult_96_n257) );
  OR3_X1 DP_mult_96_U490 ( .A1(DP_mult_96_n577), .A2(DP_sw0_0_), .A3(
        DP_mult_96_n622), .ZN(DP_mult_96_n623) );
  OAI21_X1 DP_mult_96_U489 ( .B1(DP_mult_96_n622), .B2(DP_mult_96_n579), .A(
        DP_mult_96_n623), .ZN(DP_mult_96_n258) );
  OR3_X1 DP_mult_96_U488 ( .A1(DP_mult_96_n561), .A2(DP_sw0_0_), .A3(
        DP_mult_96_n620), .ZN(DP_mult_96_n621) );
  OAI21_X1 DP_mult_96_U487 ( .B1(DP_mult_96_n620), .B2(DP_mult_96_n563), .A(
        DP_mult_96_n621), .ZN(DP_mult_96_n259) );
  XNOR2_X1 DP_mult_96_U486 ( .A(DP_sw0_10_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n619) );
  XNOR2_X1 DP_mult_96_U485 ( .A(DP_sw0_11_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n528) );
  OAI22_X1 DP_mult_96_U484 ( .A1(DP_mult_96_n619), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n528), .ZN(DP_mult_96_n263) );
  XNOR2_X1 DP_mult_96_U483 ( .A(DP_sw0_9_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n618) );
  OAI22_X1 DP_mult_96_U482 ( .A1(DP_mult_96_n618), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n619), .ZN(DP_mult_96_n264) );
  XNOR2_X1 DP_mult_96_U481 ( .A(DP_sw0_8_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n617) );
  OAI22_X1 DP_mult_96_U480 ( .A1(DP_mult_96_n617), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n618), .ZN(DP_mult_96_n265) );
  XNOR2_X1 DP_mult_96_U479 ( .A(DP_sw0_7_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n616) );
  OAI22_X1 DP_mult_96_U478 ( .A1(DP_mult_96_n616), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n617), .ZN(DP_mult_96_n266) );
  XNOR2_X1 DP_mult_96_U477 ( .A(DP_sw0_6_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n615) );
  OAI22_X1 DP_mult_96_U476 ( .A1(DP_mult_96_n615), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n616), .ZN(DP_mult_96_n267) );
  XNOR2_X1 DP_mult_96_U475 ( .A(DP_sw0_5_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n614) );
  OAI22_X1 DP_mult_96_U474 ( .A1(DP_mult_96_n614), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n615), .ZN(DP_mult_96_n268) );
  XNOR2_X1 DP_mult_96_U473 ( .A(DP_sw0_4_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n613) );
  OAI22_X1 DP_mult_96_U472 ( .A1(DP_mult_96_n613), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n614), .ZN(DP_mult_96_n269) );
  XNOR2_X1 DP_mult_96_U471 ( .A(DP_sw0_3_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n612) );
  OAI22_X1 DP_mult_96_U470 ( .A1(DP_mult_96_n612), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n613), .ZN(DP_mult_96_n270) );
  XNOR2_X1 DP_mult_96_U469 ( .A(DP_sw0_2_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n611) );
  OAI22_X1 DP_mult_96_U468 ( .A1(DP_mult_96_n611), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n612), .ZN(DP_mult_96_n271) );
  XNOR2_X1 DP_mult_96_U467 ( .A(DP_sw0_1_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n610) );
  OAI22_X1 DP_mult_96_U466 ( .A1(DP_mult_96_n610), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n611), .ZN(DP_mult_96_n272) );
  XNOR2_X1 DP_mult_96_U465 ( .A(DP_sw0_0_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n609) );
  OAI22_X1 DP_mult_96_U464 ( .A1(DP_mult_96_n609), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n610), .ZN(DP_mult_96_n273) );
  NOR2_X1 DP_mult_96_U463 ( .A1(DP_mult_96_n560), .A2(DP_mult_96_n526), .ZN(
        DP_mult_96_n274) );
  AOI21_X1 DP_mult_96_U462 ( .B1(DP_mult_96_n595), .B2(DP_mult_96_n593), .A(
        DP_mult_96_n608), .ZN(DP_mult_96_n607) );
  INV_X1 DP_mult_96_U461 ( .A(DP_mult_96_n607), .ZN(DP_mult_96_n275) );
  XNOR2_X1 DP_mult_96_U460 ( .A(DP_sw0_10_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n605) );
  OAI22_X1 DP_mult_96_U459 ( .A1(DP_mult_96_n605), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n606), .ZN(DP_mult_96_n276) );
  XNOR2_X1 DP_mult_96_U458 ( .A(DP_sw0_9_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n604) );
  OAI22_X1 DP_mult_96_U457 ( .A1(DP_mult_96_n604), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n605), .ZN(DP_mult_96_n277) );
  XNOR2_X1 DP_mult_96_U456 ( .A(DP_sw0_8_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n603) );
  OAI22_X1 DP_mult_96_U455 ( .A1(DP_mult_96_n603), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n604), .ZN(DP_mult_96_n278) );
  XNOR2_X1 DP_mult_96_U454 ( .A(DP_sw0_7_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n602) );
  OAI22_X1 DP_mult_96_U453 ( .A1(DP_mult_96_n602), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n603), .ZN(DP_mult_96_n279) );
  XNOR2_X1 DP_mult_96_U452 ( .A(DP_sw0_6_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n601) );
  OAI22_X1 DP_mult_96_U451 ( .A1(DP_mult_96_n601), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n602), .ZN(DP_mult_96_n280) );
  OAI22_X1 DP_mult_96_U450 ( .A1(DP_mult_96_n600), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n601), .ZN(DP_mult_96_n281) );
  XNOR2_X1 DP_mult_96_U449 ( .A(DP_sw0_3_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n598) );
  OAI22_X1 DP_mult_96_U448 ( .A1(DP_mult_96_n598), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n599), .ZN(DP_mult_96_n283) );
  XNOR2_X1 DP_mult_96_U447 ( .A(DP_sw0_2_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n597) );
  OAI22_X1 DP_mult_96_U446 ( .A1(DP_mult_96_n597), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n598), .ZN(DP_mult_96_n284) );
  XNOR2_X1 DP_mult_96_U445 ( .A(DP_sw0_1_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n596) );
  OAI22_X1 DP_mult_96_U444 ( .A1(DP_mult_96_n596), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n597), .ZN(DP_mult_96_n285) );
  XNOR2_X1 DP_mult_96_U443 ( .A(DP_sw0_0_), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n594) );
  OAI22_X1 DP_mult_96_U442 ( .A1(DP_mult_96_n594), .A2(DP_mult_96_n595), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n286) );
  NOR2_X1 DP_mult_96_U441 ( .A1(DP_mult_96_n560), .A2(DP_mult_96_n593), .ZN(
        DP_mult_96_n287) );
  AOI21_X1 DP_mult_96_U440 ( .B1(DP_mult_96_n579), .B2(DP_mult_96_n577), .A(
        DP_mult_96_n592), .ZN(DP_mult_96_n591) );
  INV_X1 DP_mult_96_U439 ( .A(DP_mult_96_n591), .ZN(DP_mult_96_n288) );
  XNOR2_X1 DP_mult_96_U438 ( .A(DP_sw0_10_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n589) );
  OAI22_X1 DP_mult_96_U437 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n590), .ZN(DP_mult_96_n289) );
  XNOR2_X1 DP_mult_96_U436 ( .A(DP_sw0_9_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n588) );
  OAI22_X1 DP_mult_96_U435 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n589), .ZN(DP_mult_96_n290) );
  XNOR2_X1 DP_mult_96_U434 ( .A(DP_sw0_8_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n587) );
  OAI22_X1 DP_mult_96_U433 ( .A1(DP_mult_96_n587), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n588), .ZN(DP_mult_96_n291) );
  XNOR2_X1 DP_mult_96_U432 ( .A(DP_sw0_7_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n586) );
  OAI22_X1 DP_mult_96_U431 ( .A1(DP_mult_96_n586), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n587), .ZN(DP_mult_96_n292) );
  XNOR2_X1 DP_mult_96_U430 ( .A(DP_sw0_6_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n585) );
  OAI22_X1 DP_mult_96_U429 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n586), .ZN(DP_mult_96_n293) );
  XNOR2_X1 DP_mult_96_U428 ( .A(DP_sw0_5_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n584) );
  OAI22_X1 DP_mult_96_U427 ( .A1(DP_mult_96_n584), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n585), .ZN(DP_mult_96_n294) );
  XNOR2_X1 DP_mult_96_U426 ( .A(DP_sw0_4_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n583) );
  OAI22_X1 DP_mult_96_U425 ( .A1(DP_mult_96_n583), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n584), .ZN(DP_mult_96_n295) );
  XNOR2_X1 DP_mult_96_U424 ( .A(DP_sw0_3_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n582) );
  OAI22_X1 DP_mult_96_U423 ( .A1(DP_mult_96_n582), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n583), .ZN(DP_mult_96_n296) );
  XNOR2_X1 DP_mult_96_U422 ( .A(DP_sw0_2_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n581) );
  OAI22_X1 DP_mult_96_U421 ( .A1(DP_mult_96_n581), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n582), .ZN(DP_mult_96_n297) );
  XNOR2_X1 DP_mult_96_U420 ( .A(DP_sw0_1_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n580) );
  OAI22_X1 DP_mult_96_U419 ( .A1(DP_mult_96_n580), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n581), .ZN(DP_mult_96_n298) );
  XNOR2_X1 DP_mult_96_U418 ( .A(DP_sw0_0_), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n578) );
  OAI22_X1 DP_mult_96_U417 ( .A1(DP_mult_96_n578), .A2(DP_mult_96_n579), .B1(
        DP_mult_96_n577), .B2(DP_mult_96_n580), .ZN(DP_mult_96_n299) );
  NOR2_X1 DP_mult_96_U416 ( .A1(DP_mult_96_n560), .A2(DP_mult_96_n577), .ZN(
        DP_mult_96_n300) );
  AOI21_X1 DP_mult_96_U415 ( .B1(DP_mult_96_n563), .B2(DP_mult_96_n561), .A(
        DP_mult_96_n576), .ZN(DP_mult_96_n575) );
  INV_X1 DP_mult_96_U414 ( .A(DP_mult_96_n575), .ZN(DP_mult_96_n301) );
  XNOR2_X1 DP_mult_96_U413 ( .A(DP_sw0_10_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n573) );
  OAI22_X1 DP_mult_96_U412 ( .A1(DP_mult_96_n573), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n574), .ZN(DP_mult_96_n302) );
  OAI22_X1 DP_mult_96_U411 ( .A1(DP_mult_96_n572), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n573), .ZN(DP_mult_96_n303) );
  XNOR2_X1 DP_mult_96_U410 ( .A(DP_sw0_7_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n570) );
  OAI22_X1 DP_mult_96_U409 ( .A1(DP_mult_96_n570), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n571), .ZN(DP_mult_96_n305) );
  XNOR2_X1 DP_mult_96_U408 ( .A(DP_sw0_6_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n569) );
  OAI22_X1 DP_mult_96_U407 ( .A1(DP_mult_96_n569), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n570), .ZN(DP_mult_96_n306) );
  XNOR2_X1 DP_mult_96_U406 ( .A(DP_sw0_5_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n568) );
  OAI22_X1 DP_mult_96_U405 ( .A1(DP_mult_96_n568), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n569), .ZN(DP_mult_96_n307) );
  XNOR2_X1 DP_mult_96_U404 ( .A(DP_sw0_4_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n567) );
  OAI22_X1 DP_mult_96_U403 ( .A1(DP_mult_96_n567), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n568), .ZN(DP_mult_96_n308) );
  XNOR2_X1 DP_mult_96_U402 ( .A(DP_sw0_3_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n566) );
  OAI22_X1 DP_mult_96_U401 ( .A1(DP_mult_96_n566), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n567), .ZN(DP_mult_96_n309) );
  XNOR2_X1 DP_mult_96_U400 ( .A(DP_sw0_2_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n565) );
  OAI22_X1 DP_mult_96_U399 ( .A1(DP_mult_96_n565), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n566), .ZN(DP_mult_96_n310) );
  XNOR2_X1 DP_mult_96_U398 ( .A(DP_sw0_1_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n564) );
  OAI22_X1 DP_mult_96_U397 ( .A1(DP_mult_96_n564), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n565), .ZN(DP_mult_96_n311) );
  XNOR2_X1 DP_mult_96_U396 ( .A(DP_sw0_0_), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n562) );
  OAI22_X1 DP_mult_96_U395 ( .A1(DP_mult_96_n562), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n564), .ZN(DP_mult_96_n312) );
  NOR2_X1 DP_mult_96_U394 ( .A1(DP_mult_96_n560), .A2(DP_mult_96_n561), .ZN(
        DP_mult_96_n313) );
  AOI21_X1 DP_mult_96_U393 ( .B1(DP_mult_96_n545), .B2(DP_mult_96_n546), .A(
        DP_mult_96_n559), .ZN(DP_mult_96_n558) );
  INV_X1 DP_mult_96_U392 ( .A(DP_mult_96_n558), .ZN(DP_mult_96_n314) );
  XNOR2_X1 DP_mult_96_U391 ( .A(DP_sw0_10_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n556) );
  OAI22_X1 DP_mult_96_U390 ( .A1(DP_mult_96_n556), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n557), .ZN(DP_mult_96_n315) );
  XNOR2_X1 DP_mult_96_U389 ( .A(DP_sw0_9_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n555) );
  OAI22_X1 DP_mult_96_U388 ( .A1(DP_mult_96_n555), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n556), .ZN(DP_mult_96_n316) );
  XNOR2_X1 DP_mult_96_U387 ( .A(DP_sw0_8_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n554) );
  OAI22_X1 DP_mult_96_U386 ( .A1(DP_mult_96_n554), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n555), .ZN(DP_mult_96_n317) );
  XNOR2_X1 DP_mult_96_U385 ( .A(DP_sw0_7_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n553) );
  OAI22_X1 DP_mult_96_U384 ( .A1(DP_mult_96_n553), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n554), .ZN(DP_mult_96_n318) );
  XNOR2_X1 DP_mult_96_U383 ( .A(DP_sw0_6_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n552) );
  OAI22_X1 DP_mult_96_U382 ( .A1(DP_mult_96_n552), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n553), .ZN(DP_mult_96_n319) );
  XNOR2_X1 DP_mult_96_U381 ( .A(DP_sw0_5_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n551) );
  OAI22_X1 DP_mult_96_U380 ( .A1(DP_mult_96_n551), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n552), .ZN(DP_mult_96_n320) );
  XNOR2_X1 DP_mult_96_U379 ( .A(DP_sw0_4_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n550) );
  OAI22_X1 DP_mult_96_U378 ( .A1(DP_mult_96_n550), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n551), .ZN(DP_mult_96_n321) );
  XNOR2_X1 DP_mult_96_U377 ( .A(DP_sw0_3_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n549) );
  OAI22_X1 DP_mult_96_U376 ( .A1(DP_mult_96_n549), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n550), .ZN(DP_mult_96_n322) );
  XNOR2_X1 DP_mult_96_U375 ( .A(DP_sw0_2_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n548) );
  OAI22_X1 DP_mult_96_U374 ( .A1(DP_mult_96_n548), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n549), .ZN(DP_mult_96_n323) );
  XNOR2_X1 DP_mult_96_U373 ( .A(DP_sw0_1_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n547) );
  OAI22_X1 DP_mult_96_U372 ( .A1(DP_mult_96_n547), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n548), .ZN(DP_mult_96_n324) );
  XNOR2_X1 DP_mult_96_U371 ( .A(DP_sw0_0_), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n544) );
  OAI22_X1 DP_mult_96_U370 ( .A1(DP_mult_96_n544), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n546), .B2(DP_mult_96_n547), .ZN(DP_mult_96_n325) );
  XOR2_X1 DP_mult_96_U369 ( .A(DP_sw0_12_), .B(DP_mult_96_n543), .Z(
        DP_mult_96_n541) );
  AOI21_X1 DP_mult_96_U368 ( .B1(DP_mult_96_n530), .B2(DP_mult_96_n532), .A(
        DP_mult_96_n541), .ZN(DP_mult_96_n542) );
  INV_X1 DP_mult_96_U367 ( .A(DP_mult_96_n542), .ZN(DP_mult_96_n327) );
  XNOR2_X1 DP_mult_96_U366 ( .A(DP_sw0_11_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n540) );
  OAI22_X1 DP_mult_96_U365 ( .A1(DP_mult_96_n540), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n541), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n328) );
  XNOR2_X1 DP_mult_96_U364 ( .A(DP_sw0_10_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n539) );
  OAI22_X1 DP_mult_96_U363 ( .A1(DP_mult_96_n539), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n540), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n329) );
  XNOR2_X1 DP_mult_96_U362 ( .A(DP_sw0_9_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n538) );
  OAI22_X1 DP_mult_96_U361 ( .A1(DP_mult_96_n538), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n539), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n330) );
  XNOR2_X1 DP_mult_96_U360 ( .A(DP_sw0_8_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n537) );
  OAI22_X1 DP_mult_96_U359 ( .A1(DP_mult_96_n537), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n538), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n331) );
  XNOR2_X1 DP_mult_96_U358 ( .A(DP_sw0_7_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n536) );
  OAI22_X1 DP_mult_96_U357 ( .A1(DP_mult_96_n536), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n537), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n332) );
  XNOR2_X1 DP_mult_96_U356 ( .A(DP_sw0_6_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n535) );
  OAI22_X1 DP_mult_96_U355 ( .A1(DP_mult_96_n535), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n536), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n333) );
  XNOR2_X1 DP_mult_96_U354 ( .A(DP_sw0_5_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n534) );
  OAI22_X1 DP_mult_96_U353 ( .A1(DP_mult_96_n534), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n535), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n334) );
  XNOR2_X1 DP_mult_96_U352 ( .A(DP_sw0_4_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n533) );
  OAI22_X1 DP_mult_96_U351 ( .A1(DP_mult_96_n533), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n534), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n335) );
  XNOR2_X1 DP_mult_96_U350 ( .A(DP_sw0_3_), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n531) );
  OAI22_X1 DP_mult_96_U349 ( .A1(DP_mult_96_n531), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n533), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n336) );
  OAI22_X1 DP_mult_96_U348 ( .A1(DP_mult_96_n529), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n531), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n337) );
  XNOR2_X1 DP_mult_96_U347 ( .A(DP_sw0_12_), .B(DP_a_int[0]), .ZN(
        DP_mult_96_n527) );
  OAI22_X1 DP_mult_96_U346 ( .A1(DP_mult_96_n528), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n526), .B2(DP_mult_96_n527), .ZN(DP_mult_96_n519) );
  AOI21_X1 DP_mult_96_U345 ( .B1(DP_mult_96_n525), .B2(DP_mult_96_n526), .A(
        DP_mult_96_n527), .ZN(DP_mult_96_n522) );
  INV_X1 DP_mult_96_U344 ( .A(DP_mult_96_n522), .ZN(DP_mult_96_n520) );
  INV_X1 DP_mult_96_U343 ( .A(DP_mult_96_n519), .ZN(DP_mult_96_n524) );
  AOI222_X1 DP_mult_96_U342 ( .A1(DP_mult_96_n115), .A2(DP_mult_96_n138), .B1(
        DP_mult_96_n524), .B2(DP_mult_96_n115), .C1(DP_mult_96_n524), .C2(
        DP_mult_96_n138), .ZN(DP_mult_96_n523) );
  OAI22_X1 DP_mult_96_U341 ( .A1(DP_mult_96_n522), .A2(DP_mult_96_n523), .B1(
        DP_mult_96_n524), .B2(DP_mult_96_n523), .ZN(DP_mult_96_n521) );
  AOI21_X1 DP_mult_96_U340 ( .B1(DP_mult_96_n519), .B2(DP_mult_96_n520), .A(
        DP_mult_96_n521), .ZN(DP_sw0_a1_11_) );
  XOR2_X2 DP_mult_96_U339 ( .A(DP_a_int[3]), .B(DP_mult_96_n622), .Z(
        DP_mult_96_n593) );
  XOR2_X2 DP_mult_96_U338 ( .A(DP_a_int[5]), .B(DP_mult_96_n620), .Z(
        DP_mult_96_n577) );
  XOR2_X2 DP_mult_96_U337 ( .A(DP_a_int[7]), .B(DP_mult_96_n632), .Z(
        DP_mult_96_n561) );
  XOR2_X2 DP_mult_96_U336 ( .A(DP_a_int[1]), .B(DP_mult_96_n624), .Z(
        DP_mult_96_n526) );
  INV_X1 DP_mult_96_U335 ( .A(DP_a_int[11]), .ZN(DP_mult_96_n532) );
  INV_X1 DP_mult_96_U334 ( .A(DP_mult_96_n653), .ZN(DP_mult_96_n546) );
  HA_X1 DP_mult_96_U120 ( .A(DP_mult_96_n325), .B(DP_mult_96_n337), .CO(
        DP_mult_96_n254), .S(DP_mult_96_n255) );
  FA_X1 DP_mult_96_U119 ( .A(DP_mult_96_n336), .B(DP_mult_96_n313), .CI(
        DP_mult_96_n324), .CO(DP_mult_96_n252), .S(DP_mult_96_n253) );
  HA_X1 DP_mult_96_U118 ( .A(DP_mult_96_n259), .B(DP_mult_96_n312), .CO(
        DP_mult_96_n250), .S(DP_mult_96_n251) );
  FA_X1 DP_mult_96_U117 ( .A(DP_mult_96_n323), .B(DP_mult_96_n335), .CI(
        DP_mult_96_n251), .CO(DP_mult_96_n248), .S(DP_mult_96_n249) );
  FA_X1 DP_mult_96_U109 ( .A(DP_mult_96_n334), .B(DP_mult_96_n300), .CI(
        DP_mult_96_n322), .CO(DP_mult_96_n246), .S(DP_mult_96_n247) );
  FA_X1 DP_mult_96_U108 ( .A(DP_mult_96_n250), .B(DP_mult_96_n311), .CI(
        DP_mult_96_n247), .CO(DP_mult_96_n244), .S(DP_mult_96_n245) );
  HA_X1 DP_mult_96_U107 ( .A(DP_mult_96_n258), .B(DP_mult_96_n299), .CO(
        DP_mult_96_n242), .S(DP_mult_96_n243) );
  FA_X1 DP_mult_96_U106 ( .A(DP_mult_96_n310), .B(DP_mult_96_n333), .CI(
        DP_mult_96_n321), .CO(DP_mult_96_n240), .S(DP_mult_96_n241) );
  FA_X1 DP_mult_96_U105 ( .A(DP_mult_96_n246), .B(DP_mult_96_n243), .CI(
        DP_mult_96_n241), .CO(DP_mult_96_n238), .S(DP_mult_96_n239) );
  FA_X1 DP_mult_96_U104 ( .A(DP_mult_96_n309), .B(DP_mult_96_n287), .CI(
        DP_mult_96_n332), .CO(DP_mult_96_n236), .S(DP_mult_96_n237) );
  FA_X1 DP_mult_96_U103 ( .A(DP_mult_96_n298), .B(DP_mult_96_n320), .CI(
        DP_mult_96_n242), .CO(DP_mult_96_n234), .S(DP_mult_96_n235) );
  FA_X1 DP_mult_96_U102 ( .A(DP_mult_96_n237), .B(DP_mult_96_n240), .CI(
        DP_mult_96_n235), .CO(DP_mult_96_n232), .S(DP_mult_96_n233) );
  HA_X1 DP_mult_96_U101 ( .A(DP_mult_96_n257), .B(DP_mult_96_n286), .CO(
        DP_mult_96_n230), .S(DP_mult_96_n231) );
  FA_X1 DP_mult_96_U100 ( .A(DP_mult_96_n297), .B(DP_mult_96_n308), .CI(
        DP_mult_96_n319), .CO(DP_mult_96_n228), .S(DP_mult_96_n229) );
  FA_X1 DP_mult_96_U99 ( .A(DP_mult_96_n231), .B(DP_mult_96_n331), .CI(
        DP_mult_96_n236), .CO(DP_mult_96_n226), .S(DP_mult_96_n227) );
  FA_X1 DP_mult_96_U98 ( .A(DP_mult_96_n229), .B(DP_mult_96_n234), .CI(
        DP_mult_96_n227), .CO(DP_mult_96_n224), .S(DP_mult_96_n225) );
  FA_X1 DP_mult_96_U97 ( .A(DP_mult_96_n296), .B(DP_mult_96_n274), .CI(
        DP_mult_96_n330), .CO(DP_mult_96_n222), .S(DP_mult_96_n223) );
  FA_X1 DP_mult_96_U96 ( .A(DP_mult_96_n285), .B(DP_mult_96_n318), .CI(
        DP_mult_96_n307), .CO(DP_mult_96_n220), .S(DP_mult_96_n221) );
  FA_X1 DP_mult_96_U95 ( .A(DP_mult_96_n228), .B(DP_mult_96_n230), .CI(
        DP_mult_96_n223), .CO(DP_mult_96_n218), .S(DP_mult_96_n219) );
  FA_X1 DP_mult_96_U94 ( .A(DP_mult_96_n226), .B(DP_mult_96_n221), .CI(
        DP_mult_96_n219), .CO(DP_mult_96_n216), .S(DP_mult_96_n217) );
  HA_X1 DP_mult_96_U93 ( .A(DP_mult_96_n256), .B(DP_mult_96_n273), .CO(
        DP_mult_96_n214), .S(DP_mult_96_n215) );
  FA_X1 DP_mult_96_U92 ( .A(DP_mult_96_n284), .B(DP_mult_96_n306), .CI(
        DP_mult_96_n329), .CO(DP_mult_96_n212), .S(DP_mult_96_n213) );
  FA_X1 DP_mult_96_U91 ( .A(DP_mult_96_n295), .B(DP_mult_96_n317), .CI(
        DP_mult_96_n215), .CO(DP_mult_96_n210), .S(DP_mult_96_n211) );
  FA_X1 DP_mult_96_U90 ( .A(DP_mult_96_n220), .B(DP_mult_96_n222), .CI(
        DP_mult_96_n213), .CO(DP_mult_96_n208), .S(DP_mult_96_n209) );
  FA_X1 DP_mult_96_U89 ( .A(DP_mult_96_n218), .B(DP_mult_96_n211), .CI(
        DP_mult_96_n209), .CO(DP_mult_96_n206), .S(DP_mult_96_n207) );
  HA_X1 DP_mult_96_U88 ( .A(DP_mult_96_n272), .B(DP_mult_96_n283), .CO(
        DP_mult_96_n204), .S(DP_mult_96_n205) );
  FA_X1 DP_mult_96_U87 ( .A(DP_mult_96_n328), .B(DP_mult_96_n305), .CI(
        DP_mult_96_n294), .CO(DP_mult_96_n202), .S(DP_mult_96_n203) );
  FA_X1 DP_mult_96_U86 ( .A(DP_mult_96_n214), .B(DP_mult_96_n316), .CI(
        DP_mult_96_n205), .CO(DP_mult_96_n200), .S(DP_mult_96_n201) );
  FA_X1 DP_mult_96_U85 ( .A(DP_mult_96_n203), .B(DP_mult_96_n212), .CI(
        DP_mult_96_n210), .CO(DP_mult_96_n198), .S(DP_mult_96_n199) );
  FA_X1 DP_mult_96_U84 ( .A(DP_mult_96_n208), .B(DP_mult_96_n201), .CI(
        DP_mult_96_n199), .CO(DP_mult_96_n196), .S(DP_mult_96_n197) );
  FA_X1 DP_mult_96_U81 ( .A(DP_mult_96_n271), .B(DP_mult_96_n293), .CI(
        DP_mult_96_n327), .CO(DP_mult_96_n192), .S(DP_mult_96_n193) );
  FA_X1 DP_mult_96_U80 ( .A(DP_mult_96_n204), .B(DP_mult_96_n315), .CI(
        DP_mult_96_n195), .CO(DP_mult_96_n190), .S(DP_mult_96_n191) );
  FA_X1 DP_mult_96_U79 ( .A(DP_mult_96_n193), .B(DP_mult_96_n202), .CI(
        DP_mult_96_n200), .CO(DP_mult_96_n188), .S(DP_mult_96_n189) );
  FA_X1 DP_mult_96_U78 ( .A(DP_mult_96_n198), .B(DP_mult_96_n191), .CI(
        DP_mult_96_n189), .CO(DP_mult_96_n186), .S(DP_mult_96_n187) );
  FA_X1 DP_mult_96_U76 ( .A(DP_mult_96_n303), .B(DP_mult_96_n281), .CI(
        DP_mult_96_n185), .CO(DP_mult_96_n182), .S(DP_mult_96_n183) );
  FA_X1 DP_mult_96_U75 ( .A(DP_mult_96_n270), .B(DP_mult_96_n292), .CI(
        DP_mult_96_n194), .CO(DP_mult_96_n180), .S(DP_mult_96_n181) );
  FA_X1 DP_mult_96_U74 ( .A(DP_mult_96_n190), .B(DP_mult_96_n192), .CI(
        DP_mult_96_n183), .CO(DP_mult_96_n178), .S(DP_mult_96_n179) );
  FA_X1 DP_mult_96_U73 ( .A(DP_mult_96_n188), .B(DP_mult_96_n181), .CI(
        DP_mult_96_n179), .CO(DP_mult_96_n176), .S(DP_mult_96_n177) );
  FA_X1 DP_mult_96_U72 ( .A(DP_mult_96_n184), .B(DP_mult_96_n269), .CI(
        DP_mult_96_n314), .CO(DP_mult_96_n174), .S(DP_mult_96_n175) );
  FA_X1 DP_mult_96_U71 ( .A(DP_mult_96_n280), .B(DP_mult_96_n302), .CI(
        DP_mult_96_n291), .CO(DP_mult_96_n172), .S(DP_mult_96_n173) );
  FA_X1 DP_mult_96_U70 ( .A(DP_mult_96_n180), .B(DP_mult_96_n182), .CI(
        DP_mult_96_n173), .CO(DP_mult_96_n170), .S(DP_mult_96_n171) );
  FA_X1 DP_mult_96_U69 ( .A(DP_mult_96_n178), .B(DP_mult_96_n175), .CI(
        DP_mult_96_n171), .CO(DP_mult_96_n168), .S(DP_mult_96_n169) );
  FA_X1 DP_mult_96_U67 ( .A(DP_mult_96_n268), .B(DP_mult_96_n279), .CI(
        DP_mult_96_n167), .CO(DP_mult_96_n164), .S(DP_mult_96_n165) );
  FA_X1 DP_mult_96_U66 ( .A(DP_mult_96_n174), .B(DP_mult_96_n290), .CI(
        DP_mult_96_n172), .CO(DP_mult_96_n162), .S(DP_mult_96_n163) );
  FA_X1 DP_mult_96_U65 ( .A(DP_mult_96_n170), .B(DP_mult_96_n165), .CI(
        DP_mult_96_n163), .CO(DP_mult_96_n160), .S(DP_mult_96_n161) );
  FA_X1 DP_mult_96_U64 ( .A(DP_mult_96_n166), .B(DP_mult_96_n267), .CI(
        DP_mult_96_n301), .CO(DP_mult_96_n158), .S(DP_mult_96_n159) );
  FA_X1 DP_mult_96_U63 ( .A(DP_mult_96_n278), .B(DP_mult_96_n289), .CI(
        DP_mult_96_n164), .CO(DP_mult_96_n156), .S(DP_mult_96_n157) );
  FA_X1 DP_mult_96_U62 ( .A(DP_mult_96_n162), .B(DP_mult_96_n159), .CI(
        DP_mult_96_n157), .CO(DP_mult_96_n154), .S(DP_mult_96_n155) );
  FA_X1 DP_mult_96_U60 ( .A(DP_mult_96_n266), .B(DP_mult_96_n277), .CI(
        DP_mult_96_n153), .CO(DP_mult_96_n150), .S(DP_mult_96_n151) );
  FA_X1 DP_mult_96_U59 ( .A(DP_mult_96_n151), .B(DP_mult_96_n158), .CI(
        DP_mult_96_n156), .CO(DP_mult_96_n148), .S(DP_mult_96_n149) );
  FA_X1 DP_mult_96_U58 ( .A(DP_mult_96_n265), .B(DP_mult_96_n152), .CI(
        DP_mult_96_n288), .CO(DP_mult_96_n146), .S(DP_mult_96_n147) );
  FA_X1 DP_mult_96_U57 ( .A(DP_mult_96_n150), .B(DP_mult_96_n276), .CI(
        DP_mult_96_n147), .CO(DP_mult_96_n144), .S(DP_mult_96_n145) );
  FA_X1 DP_mult_96_U55 ( .A(DP_mult_96_n143), .B(DP_mult_96_n264), .CI(
        DP_mult_96_n146), .CO(DP_mult_96_n140), .S(DP_mult_96_n141) );
  FA_X1 DP_mult_96_U54 ( .A(DP_mult_96_n263), .B(DP_mult_96_n142), .CI(
        DP_mult_96_n275), .CO(DP_mult_96_n138), .S(DP_mult_96_n139) );
  FA_X1 DP_mult_96_U42 ( .A(DP_mult_96_n207), .B(DP_mult_96_n216), .CI(
        DP_mult_96_n126), .CO(DP_mult_96_n125), .S(DP_sw0_a1_0_) );
  FA_X1 DP_mult_96_U41 ( .A(DP_mult_96_n197), .B(DP_mult_96_n206), .CI(
        DP_mult_96_n125), .CO(DP_mult_96_n124), .S(DP_sw0_a1_1_) );
  FA_X1 DP_mult_96_U40 ( .A(DP_mult_96_n187), .B(DP_mult_96_n196), .CI(
        DP_mult_96_n124), .CO(DP_mult_96_n123), .S(DP_sw0_a1_2_) );
  FA_X1 DP_mult_96_U39 ( .A(DP_mult_96_n177), .B(DP_mult_96_n186), .CI(
        DP_mult_96_n123), .CO(DP_mult_96_n122), .S(DP_sw0_a1_3_) );
  FA_X1 DP_mult_96_U38 ( .A(DP_mult_96_n169), .B(DP_mult_96_n176), .CI(
        DP_mult_96_n122), .CO(DP_mult_96_n121), .S(DP_sw0_a1_4_) );
  FA_X1 DP_mult_96_U37 ( .A(DP_mult_96_n161), .B(DP_mult_96_n168), .CI(
        DP_mult_96_n121), .CO(DP_mult_96_n120), .S(DP_sw0_a1_5_) );
  FA_X1 DP_mult_96_U36 ( .A(DP_mult_96_n155), .B(DP_mult_96_n160), .CI(
        DP_mult_96_n120), .CO(DP_mult_96_n119), .S(DP_sw0_a1_6_) );
  FA_X1 DP_mult_96_U30 ( .A(DP_mult_96_n149), .B(DP_mult_96_n154), .CI(
        DP_mult_96_n119), .CO(DP_mult_96_n118), .S(DP_sw0_a1_7_) );
  FA_X1 DP_mult_96_U20 ( .A(DP_mult_96_n145), .B(DP_mult_96_n148), .CI(
        DP_mult_96_n118), .CO(DP_mult_96_n117), .S(DP_sw0_a1_8_) );
  FA_X1 DP_mult_96_U10 ( .A(DP_mult_96_n141), .B(DP_mult_96_n144), .CI(
        DP_mult_96_n117), .CO(DP_mult_96_n116), .S(DP_sw0_a1_9_) );
  FA_X1 DP_mult_96_U9 ( .A(DP_mult_96_n140), .B(DP_mult_96_n139), .CI(
        DP_mult_96_n116), .CO(DP_mult_96_n115), .S(DP_sw0_a1_10_) );
  XOR2_X1 DP_mult_98_U563 ( .A(DP_b_int[21]), .B(DP_b_int[22]), .Z(
        DP_mult_98_n653) );
  INV_X1 DP_mult_98_U562 ( .A(DP_b_int[22]), .ZN(DP_mult_98_n543) );
  NOR2_X1 DP_mult_98_U561 ( .A1(DP_mult_98_n543), .A2(DP_sw0_1_), .ZN(
        DP_mult_98_n658) );
  INV_X1 DP_mult_98_U560 ( .A(DP_mult_98_n658), .ZN(DP_mult_98_n660) );
  NAND2_X1 DP_mult_98_U559 ( .A1(DP_b_int[22]), .A2(DP_mult_98_n532), .ZN(
        DP_mult_98_n530) );
  XNOR2_X1 DP_mult_98_U558 ( .A(DP_sw0_2_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n529) );
  OAI22_X1 DP_mult_98_U557 ( .A1(DP_mult_98_n660), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n529), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n659) );
  NAND2_X1 DP_mult_98_U556 ( .A1(DP_mult_98_n653), .A2(DP_mult_98_n659), .ZN(
        DP_mult_98_n656) );
  NAND2_X1 DP_mult_98_U555 ( .A1(DP_mult_98_n658), .A2(DP_mult_98_n659), .ZN(
        DP_mult_98_n657) );
  INV_X1 DP_mult_98_U554 ( .A(DP_sw0_0_), .ZN(DP_mult_98_n560) );
  MUX2_X1 DP_mult_98_U553 ( .A(DP_mult_98_n656), .B(DP_mult_98_n657), .S(
        DP_mult_98_n560), .Z(DP_mult_98_n655) );
  INV_X1 DP_mult_98_U552 ( .A(DP_mult_98_n655), .ZN(DP_mult_98_n650) );
  INV_X1 DP_mult_98_U551 ( .A(DP_b_int[20]), .ZN(DP_mult_98_n632) );
  XNOR2_X1 DP_mult_98_U550 ( .A(DP_mult_98_n632), .B(DP_b_int[21]), .ZN(
        DP_mult_98_n654) );
  NAND2_X1 DP_mult_98_U549 ( .A1(DP_mult_98_n546), .A2(DP_mult_98_n654), .ZN(
        DP_mult_98_n545) );
  NAND3_X1 DP_mult_98_U548 ( .A1(DP_mult_98_n653), .A2(DP_mult_98_n560), .A3(
        DP_b_int[20]), .ZN(DP_mult_98_n652) );
  OAI21_X1 DP_mult_98_U547 ( .B1(DP_mult_98_n632), .B2(DP_mult_98_n545), .A(
        DP_mult_98_n652), .ZN(DP_mult_98_n651) );
  AOI222_X1 DP_mult_98_U546 ( .A1(DP_mult_98_n650), .A2(DP_mult_98_n255), .B1(
        DP_mult_98_n651), .B2(DP_mult_98_n650), .C1(DP_mult_98_n651), .C2(
        DP_mult_98_n255), .ZN(DP_mult_98_n649) );
  INV_X1 DP_mult_98_U545 ( .A(DP_mult_98_n649), .ZN(DP_mult_98_n648) );
  AOI222_X1 DP_mult_98_U544 ( .A1(DP_mult_98_n648), .A2(DP_mult_98_n253), .B1(
        DP_mult_98_n648), .B2(DP_mult_98_n254), .C1(DP_mult_98_n254), .C2(
        DP_mult_98_n253), .ZN(DP_mult_98_n647) );
  INV_X1 DP_mult_98_U543 ( .A(DP_mult_98_n647), .ZN(DP_mult_98_n646) );
  AOI222_X1 DP_mult_98_U542 ( .A1(DP_mult_98_n646), .A2(DP_mult_98_n249), .B1(
        DP_mult_98_n646), .B2(DP_mult_98_n252), .C1(DP_mult_98_n252), .C2(
        DP_mult_98_n249), .ZN(DP_mult_98_n645) );
  INV_X1 DP_mult_98_U541 ( .A(DP_mult_98_n645), .ZN(DP_mult_98_n644) );
  AOI222_X1 DP_mult_98_U540 ( .A1(DP_mult_98_n644), .A2(DP_mult_98_n245), .B1(
        DP_mult_98_n644), .B2(DP_mult_98_n248), .C1(DP_mult_98_n248), .C2(
        DP_mult_98_n245), .ZN(DP_mult_98_n643) );
  INV_X1 DP_mult_98_U539 ( .A(DP_mult_98_n643), .ZN(DP_mult_98_n642) );
  AOI222_X1 DP_mult_98_U538 ( .A1(DP_mult_98_n642), .A2(DP_mult_98_n239), .B1(
        DP_mult_98_n642), .B2(DP_mult_98_n244), .C1(DP_mult_98_n244), .C2(
        DP_mult_98_n239), .ZN(DP_mult_98_n639) );
  INV_X1 DP_mult_98_U537 ( .A(DP_mult_98_n233), .ZN(DP_mult_98_n640) );
  INV_X1 DP_mult_98_U536 ( .A(DP_mult_98_n238), .ZN(DP_mult_98_n641) );
  OAI222_X1 DP_mult_98_U535 ( .A1(DP_mult_98_n639), .A2(DP_mult_98_n640), .B1(
        DP_mult_98_n639), .B2(DP_mult_98_n641), .C1(DP_mult_98_n641), .C2(
        DP_mult_98_n640), .ZN(DP_mult_98_n638) );
  AOI222_X1 DP_mult_98_U534 ( .A1(DP_mult_98_n638), .A2(DP_mult_98_n225), .B1(
        DP_mult_98_n638), .B2(DP_mult_98_n232), .C1(DP_mult_98_n232), .C2(
        DP_mult_98_n225), .ZN(DP_mult_98_n635) );
  INV_X1 DP_mult_98_U533 ( .A(DP_mult_98_n217), .ZN(DP_mult_98_n636) );
  INV_X1 DP_mult_98_U532 ( .A(DP_mult_98_n224), .ZN(DP_mult_98_n637) );
  OAI222_X1 DP_mult_98_U531 ( .A1(DP_mult_98_n635), .A2(DP_mult_98_n636), .B1(
        DP_mult_98_n635), .B2(DP_mult_98_n637), .C1(DP_mult_98_n637), .C2(
        DP_mult_98_n636), .ZN(DP_mult_98_n126) );
  XNOR2_X1 DP_mult_98_U530 ( .A(DP_sw0_11_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n606) );
  INV_X1 DP_mult_98_U529 ( .A(DP_b_int[16]), .ZN(DP_mult_98_n622) );
  INV_X1 DP_mult_98_U528 ( .A(DP_b_int[14]), .ZN(DP_mult_98_n624) );
  XNOR2_X1 DP_mult_98_U527 ( .A(DP_mult_98_n624), .B(DP_b_int[15]), .ZN(
        DP_mult_98_n634) );
  NAND2_X1 DP_mult_98_U526 ( .A1(DP_mult_98_n593), .A2(DP_mult_98_n634), .ZN(
        DP_mult_98_n595) );
  XNOR2_X1 DP_mult_98_U525 ( .A(DP_sw0_12_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n608) );
  OAI22_X1 DP_mult_98_U524 ( .A1(DP_mult_98_n606), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n608), .ZN(DP_mult_98_n142) );
  INV_X1 DP_mult_98_U523 ( .A(DP_mult_98_n142), .ZN(DP_mult_98_n143) );
  XNOR2_X1 DP_mult_98_U522 ( .A(DP_sw0_11_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n590) );
  INV_X1 DP_mult_98_U521 ( .A(DP_b_int[18]), .ZN(DP_mult_98_n620) );
  XNOR2_X1 DP_mult_98_U520 ( .A(DP_mult_98_n622), .B(DP_b_int[17]), .ZN(
        DP_mult_98_n633) );
  NAND2_X1 DP_mult_98_U519 ( .A1(DP_mult_98_n577), .A2(DP_mult_98_n633), .ZN(
        DP_mult_98_n579) );
  XNOR2_X1 DP_mult_98_U518 ( .A(DP_sw0_12_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n592) );
  OAI22_X1 DP_mult_98_U517 ( .A1(DP_mult_98_n590), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n592), .ZN(DP_mult_98_n152) );
  INV_X1 DP_mult_98_U516 ( .A(DP_mult_98_n152), .ZN(DP_mult_98_n153) );
  XNOR2_X1 DP_mult_98_U515 ( .A(DP_sw0_11_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n574) );
  XNOR2_X1 DP_mult_98_U514 ( .A(DP_mult_98_n620), .B(DP_b_int[19]), .ZN(
        DP_mult_98_n631) );
  NAND2_X1 DP_mult_98_U513 ( .A1(DP_mult_98_n561), .A2(DP_mult_98_n631), .ZN(
        DP_mult_98_n563) );
  XNOR2_X1 DP_mult_98_U512 ( .A(DP_sw0_12_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n576) );
  OAI22_X1 DP_mult_98_U511 ( .A1(DP_mult_98_n574), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n576), .ZN(DP_mult_98_n166) );
  INV_X1 DP_mult_98_U510 ( .A(DP_mult_98_n166), .ZN(DP_mult_98_n167) );
  XNOR2_X1 DP_mult_98_U509 ( .A(DP_sw0_11_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n557) );
  XNOR2_X1 DP_mult_98_U508 ( .A(DP_sw0_12_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n559) );
  OAI22_X1 DP_mult_98_U507 ( .A1(DP_mult_98_n557), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n559), .ZN(DP_mult_98_n184) );
  INV_X1 DP_mult_98_U506 ( .A(DP_mult_98_n184), .ZN(DP_mult_98_n185) );
  XNOR2_X1 DP_mult_98_U505 ( .A(DP_sw0_4_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n599) );
  XNOR2_X1 DP_mult_98_U504 ( .A(DP_sw0_5_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n600) );
  OAI22_X1 DP_mult_98_U503 ( .A1(DP_mult_98_n599), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n600), .ZN(DP_mult_98_n629) );
  XNOR2_X1 DP_mult_98_U502 ( .A(DP_sw0_8_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n571) );
  XNOR2_X1 DP_mult_98_U501 ( .A(DP_sw0_9_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n572) );
  OAI22_X1 DP_mult_98_U500 ( .A1(DP_mult_98_n571), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n572), .ZN(DP_mult_98_n630) );
  OR2_X1 DP_mult_98_U499 ( .A1(DP_mult_98_n629), .A2(DP_mult_98_n630), .ZN(
        DP_mult_98_n194) );
  XNOR2_X1 DP_mult_98_U498 ( .A(DP_mult_98_n629), .B(DP_mult_98_n630), .ZN(
        DP_mult_98_n195) );
  INV_X1 DP_mult_98_U497 ( .A(DP_b_int[12]), .ZN(DP_mult_98_n626) );
  XNOR2_X1 DP_mult_98_U496 ( .A(DP_mult_98_n626), .B(DP_b_int[13]), .ZN(
        DP_mult_98_n628) );
  NAND2_X1 DP_mult_98_U495 ( .A1(DP_mult_98_n526), .A2(DP_mult_98_n628), .ZN(
        DP_mult_98_n525) );
  OR3_X1 DP_mult_98_U494 ( .A1(DP_mult_98_n526), .A2(DP_sw0_0_), .A3(
        DP_mult_98_n626), .ZN(DP_mult_98_n627) );
  OAI21_X1 DP_mult_98_U493 ( .B1(DP_mult_98_n626), .B2(DP_mult_98_n525), .A(
        DP_mult_98_n627), .ZN(DP_mult_98_n256) );
  OR3_X1 DP_mult_98_U492 ( .A1(DP_mult_98_n593), .A2(DP_sw0_0_), .A3(
        DP_mult_98_n624), .ZN(DP_mult_98_n625) );
  OAI21_X1 DP_mult_98_U491 ( .B1(DP_mult_98_n624), .B2(DP_mult_98_n595), .A(
        DP_mult_98_n625), .ZN(DP_mult_98_n257) );
  OR3_X1 DP_mult_98_U490 ( .A1(DP_mult_98_n577), .A2(DP_sw0_0_), .A3(
        DP_mult_98_n622), .ZN(DP_mult_98_n623) );
  OAI21_X1 DP_mult_98_U489 ( .B1(DP_mult_98_n622), .B2(DP_mult_98_n579), .A(
        DP_mult_98_n623), .ZN(DP_mult_98_n258) );
  OR3_X1 DP_mult_98_U488 ( .A1(DP_mult_98_n561), .A2(DP_sw0_0_), .A3(
        DP_mult_98_n620), .ZN(DP_mult_98_n621) );
  OAI21_X1 DP_mult_98_U487 ( .B1(DP_mult_98_n620), .B2(DP_mult_98_n563), .A(
        DP_mult_98_n621), .ZN(DP_mult_98_n259) );
  XNOR2_X1 DP_mult_98_U486 ( .A(DP_sw0_10_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n619) );
  XNOR2_X1 DP_mult_98_U485 ( .A(DP_sw0_11_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n528) );
  OAI22_X1 DP_mult_98_U484 ( .A1(DP_mult_98_n619), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n528), .ZN(DP_mult_98_n263) );
  XNOR2_X1 DP_mult_98_U483 ( .A(DP_sw0_9_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n618) );
  OAI22_X1 DP_mult_98_U482 ( .A1(DP_mult_98_n618), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n619), .ZN(DP_mult_98_n264) );
  XNOR2_X1 DP_mult_98_U481 ( .A(DP_sw0_8_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n617) );
  OAI22_X1 DP_mult_98_U480 ( .A1(DP_mult_98_n617), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n618), .ZN(DP_mult_98_n265) );
  XNOR2_X1 DP_mult_98_U479 ( .A(DP_sw0_7_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n616) );
  OAI22_X1 DP_mult_98_U478 ( .A1(DP_mult_98_n616), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n617), .ZN(DP_mult_98_n266) );
  XNOR2_X1 DP_mult_98_U477 ( .A(DP_sw0_6_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n615) );
  OAI22_X1 DP_mult_98_U476 ( .A1(DP_mult_98_n615), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n616), .ZN(DP_mult_98_n267) );
  XNOR2_X1 DP_mult_98_U475 ( .A(DP_sw0_5_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n614) );
  OAI22_X1 DP_mult_98_U474 ( .A1(DP_mult_98_n614), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n615), .ZN(DP_mult_98_n268) );
  XNOR2_X1 DP_mult_98_U473 ( .A(DP_sw0_4_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n613) );
  OAI22_X1 DP_mult_98_U472 ( .A1(DP_mult_98_n613), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n614), .ZN(DP_mult_98_n269) );
  XNOR2_X1 DP_mult_98_U471 ( .A(DP_sw0_3_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n612) );
  OAI22_X1 DP_mult_98_U470 ( .A1(DP_mult_98_n612), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n613), .ZN(DP_mult_98_n270) );
  XNOR2_X1 DP_mult_98_U469 ( .A(DP_sw0_2_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n611) );
  OAI22_X1 DP_mult_98_U468 ( .A1(DP_mult_98_n611), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n612), .ZN(DP_mult_98_n271) );
  XNOR2_X1 DP_mult_98_U467 ( .A(DP_sw0_1_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n610) );
  OAI22_X1 DP_mult_98_U466 ( .A1(DP_mult_98_n610), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n611), .ZN(DP_mult_98_n272) );
  XNOR2_X1 DP_mult_98_U465 ( .A(DP_sw0_0_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n609) );
  OAI22_X1 DP_mult_98_U464 ( .A1(DP_mult_98_n609), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n610), .ZN(DP_mult_98_n273) );
  NOR2_X1 DP_mult_98_U463 ( .A1(DP_mult_98_n560), .A2(DP_mult_98_n526), .ZN(
        DP_mult_98_n274) );
  AOI21_X1 DP_mult_98_U462 ( .B1(DP_mult_98_n595), .B2(DP_mult_98_n593), .A(
        DP_mult_98_n608), .ZN(DP_mult_98_n607) );
  INV_X1 DP_mult_98_U461 ( .A(DP_mult_98_n607), .ZN(DP_mult_98_n275) );
  XNOR2_X1 DP_mult_98_U460 ( .A(DP_sw0_10_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n605) );
  OAI22_X1 DP_mult_98_U459 ( .A1(DP_mult_98_n605), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n606), .ZN(DP_mult_98_n276) );
  XNOR2_X1 DP_mult_98_U458 ( .A(DP_sw0_9_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n604) );
  OAI22_X1 DP_mult_98_U457 ( .A1(DP_mult_98_n604), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n605), .ZN(DP_mult_98_n277) );
  XNOR2_X1 DP_mult_98_U456 ( .A(DP_sw0_8_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n603) );
  OAI22_X1 DP_mult_98_U455 ( .A1(DP_mult_98_n603), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n604), .ZN(DP_mult_98_n278) );
  XNOR2_X1 DP_mult_98_U454 ( .A(DP_sw0_7_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n602) );
  OAI22_X1 DP_mult_98_U453 ( .A1(DP_mult_98_n602), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n603), .ZN(DP_mult_98_n279) );
  XNOR2_X1 DP_mult_98_U452 ( .A(DP_sw0_6_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n601) );
  OAI22_X1 DP_mult_98_U451 ( .A1(DP_mult_98_n601), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n602), .ZN(DP_mult_98_n280) );
  OAI22_X1 DP_mult_98_U450 ( .A1(DP_mult_98_n600), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n601), .ZN(DP_mult_98_n281) );
  XNOR2_X1 DP_mult_98_U449 ( .A(DP_sw0_3_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n598) );
  OAI22_X1 DP_mult_98_U448 ( .A1(DP_mult_98_n598), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n599), .ZN(DP_mult_98_n283) );
  XNOR2_X1 DP_mult_98_U447 ( .A(DP_sw0_2_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n597) );
  OAI22_X1 DP_mult_98_U446 ( .A1(DP_mult_98_n597), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n598), .ZN(DP_mult_98_n284) );
  XNOR2_X1 DP_mult_98_U445 ( .A(DP_sw0_1_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n596) );
  OAI22_X1 DP_mult_98_U444 ( .A1(DP_mult_98_n596), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n597), .ZN(DP_mult_98_n285) );
  XNOR2_X1 DP_mult_98_U443 ( .A(DP_sw0_0_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n594) );
  OAI22_X1 DP_mult_98_U442 ( .A1(DP_mult_98_n594), .A2(DP_mult_98_n595), .B1(
        DP_mult_98_n593), .B2(DP_mult_98_n596), .ZN(DP_mult_98_n286) );
  NOR2_X1 DP_mult_98_U441 ( .A1(DP_mult_98_n560), .A2(DP_mult_98_n593), .ZN(
        DP_mult_98_n287) );
  AOI21_X1 DP_mult_98_U440 ( .B1(DP_mult_98_n579), .B2(DP_mult_98_n577), .A(
        DP_mult_98_n592), .ZN(DP_mult_98_n591) );
  INV_X1 DP_mult_98_U439 ( .A(DP_mult_98_n591), .ZN(DP_mult_98_n288) );
  XNOR2_X1 DP_mult_98_U438 ( .A(DP_sw0_10_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n589) );
  OAI22_X1 DP_mult_98_U437 ( .A1(DP_mult_98_n589), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n590), .ZN(DP_mult_98_n289) );
  XNOR2_X1 DP_mult_98_U436 ( .A(DP_sw0_9_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n588) );
  OAI22_X1 DP_mult_98_U435 ( .A1(DP_mult_98_n588), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n589), .ZN(DP_mult_98_n290) );
  XNOR2_X1 DP_mult_98_U434 ( .A(DP_sw0_8_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n587) );
  OAI22_X1 DP_mult_98_U433 ( .A1(DP_mult_98_n587), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n588), .ZN(DP_mult_98_n291) );
  XNOR2_X1 DP_mult_98_U432 ( .A(DP_sw0_7_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n586) );
  OAI22_X1 DP_mult_98_U431 ( .A1(DP_mult_98_n586), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n587), .ZN(DP_mult_98_n292) );
  XNOR2_X1 DP_mult_98_U430 ( .A(DP_sw0_6_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n585) );
  OAI22_X1 DP_mult_98_U429 ( .A1(DP_mult_98_n585), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n586), .ZN(DP_mult_98_n293) );
  XNOR2_X1 DP_mult_98_U428 ( .A(DP_sw0_5_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n584) );
  OAI22_X1 DP_mult_98_U427 ( .A1(DP_mult_98_n584), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n585), .ZN(DP_mult_98_n294) );
  XNOR2_X1 DP_mult_98_U426 ( .A(DP_sw0_4_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n583) );
  OAI22_X1 DP_mult_98_U425 ( .A1(DP_mult_98_n583), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n584), .ZN(DP_mult_98_n295) );
  XNOR2_X1 DP_mult_98_U424 ( .A(DP_sw0_3_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n582) );
  OAI22_X1 DP_mult_98_U423 ( .A1(DP_mult_98_n582), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n583), .ZN(DP_mult_98_n296) );
  XNOR2_X1 DP_mult_98_U422 ( .A(DP_sw0_2_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n581) );
  OAI22_X1 DP_mult_98_U421 ( .A1(DP_mult_98_n581), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n582), .ZN(DP_mult_98_n297) );
  XNOR2_X1 DP_mult_98_U420 ( .A(DP_sw0_1_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n580) );
  OAI22_X1 DP_mult_98_U419 ( .A1(DP_mult_98_n580), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n581), .ZN(DP_mult_98_n298) );
  XNOR2_X1 DP_mult_98_U418 ( .A(DP_sw0_0_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n578) );
  OAI22_X1 DP_mult_98_U417 ( .A1(DP_mult_98_n578), .A2(DP_mult_98_n579), .B1(
        DP_mult_98_n577), .B2(DP_mult_98_n580), .ZN(DP_mult_98_n299) );
  NOR2_X1 DP_mult_98_U416 ( .A1(DP_mult_98_n560), .A2(DP_mult_98_n577), .ZN(
        DP_mult_98_n300) );
  AOI21_X1 DP_mult_98_U415 ( .B1(DP_mult_98_n563), .B2(DP_mult_98_n561), .A(
        DP_mult_98_n576), .ZN(DP_mult_98_n575) );
  INV_X1 DP_mult_98_U414 ( .A(DP_mult_98_n575), .ZN(DP_mult_98_n301) );
  XNOR2_X1 DP_mult_98_U413 ( .A(DP_sw0_10_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n573) );
  OAI22_X1 DP_mult_98_U412 ( .A1(DP_mult_98_n573), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n574), .ZN(DP_mult_98_n302) );
  OAI22_X1 DP_mult_98_U411 ( .A1(DP_mult_98_n572), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n573), .ZN(DP_mult_98_n303) );
  XNOR2_X1 DP_mult_98_U410 ( .A(DP_sw0_7_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n570) );
  OAI22_X1 DP_mult_98_U409 ( .A1(DP_mult_98_n570), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n571), .ZN(DP_mult_98_n305) );
  XNOR2_X1 DP_mult_98_U408 ( .A(DP_sw0_6_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n569) );
  OAI22_X1 DP_mult_98_U407 ( .A1(DP_mult_98_n569), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n570), .ZN(DP_mult_98_n306) );
  XNOR2_X1 DP_mult_98_U406 ( .A(DP_sw0_5_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n568) );
  OAI22_X1 DP_mult_98_U405 ( .A1(DP_mult_98_n568), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n569), .ZN(DP_mult_98_n307) );
  XNOR2_X1 DP_mult_98_U404 ( .A(DP_sw0_4_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n567) );
  OAI22_X1 DP_mult_98_U403 ( .A1(DP_mult_98_n567), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n568), .ZN(DP_mult_98_n308) );
  XNOR2_X1 DP_mult_98_U402 ( .A(DP_sw0_3_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n566) );
  OAI22_X1 DP_mult_98_U401 ( .A1(DP_mult_98_n566), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n567), .ZN(DP_mult_98_n309) );
  XNOR2_X1 DP_mult_98_U400 ( .A(DP_sw0_2_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n565) );
  OAI22_X1 DP_mult_98_U399 ( .A1(DP_mult_98_n565), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n566), .ZN(DP_mult_98_n310) );
  XNOR2_X1 DP_mult_98_U398 ( .A(DP_sw0_1_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n564) );
  OAI22_X1 DP_mult_98_U397 ( .A1(DP_mult_98_n564), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n565), .ZN(DP_mult_98_n311) );
  XNOR2_X1 DP_mult_98_U396 ( .A(DP_sw0_0_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n562) );
  OAI22_X1 DP_mult_98_U395 ( .A1(DP_mult_98_n562), .A2(DP_mult_98_n563), .B1(
        DP_mult_98_n561), .B2(DP_mult_98_n564), .ZN(DP_mult_98_n312) );
  NOR2_X1 DP_mult_98_U394 ( .A1(DP_mult_98_n560), .A2(DP_mult_98_n561), .ZN(
        DP_mult_98_n313) );
  AOI21_X1 DP_mult_98_U393 ( .B1(DP_mult_98_n545), .B2(DP_mult_98_n546), .A(
        DP_mult_98_n559), .ZN(DP_mult_98_n558) );
  INV_X1 DP_mult_98_U392 ( .A(DP_mult_98_n558), .ZN(DP_mult_98_n314) );
  XNOR2_X1 DP_mult_98_U391 ( .A(DP_sw0_10_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n556) );
  OAI22_X1 DP_mult_98_U390 ( .A1(DP_mult_98_n556), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n557), .ZN(DP_mult_98_n315) );
  XNOR2_X1 DP_mult_98_U389 ( .A(DP_sw0_9_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n555) );
  OAI22_X1 DP_mult_98_U388 ( .A1(DP_mult_98_n555), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n556), .ZN(DP_mult_98_n316) );
  XNOR2_X1 DP_mult_98_U387 ( .A(DP_sw0_8_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n554) );
  OAI22_X1 DP_mult_98_U386 ( .A1(DP_mult_98_n554), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n555), .ZN(DP_mult_98_n317) );
  XNOR2_X1 DP_mult_98_U385 ( .A(DP_sw0_7_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n553) );
  OAI22_X1 DP_mult_98_U384 ( .A1(DP_mult_98_n553), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n554), .ZN(DP_mult_98_n318) );
  XNOR2_X1 DP_mult_98_U383 ( .A(DP_sw0_6_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n552) );
  OAI22_X1 DP_mult_98_U382 ( .A1(DP_mult_98_n552), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n553), .ZN(DP_mult_98_n319) );
  XNOR2_X1 DP_mult_98_U381 ( .A(DP_sw0_5_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n551) );
  OAI22_X1 DP_mult_98_U380 ( .A1(DP_mult_98_n551), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n552), .ZN(DP_mult_98_n320) );
  XNOR2_X1 DP_mult_98_U379 ( .A(DP_sw0_4_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n550) );
  OAI22_X1 DP_mult_98_U378 ( .A1(DP_mult_98_n550), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n551), .ZN(DP_mult_98_n321) );
  XNOR2_X1 DP_mult_98_U377 ( .A(DP_sw0_3_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n549) );
  OAI22_X1 DP_mult_98_U376 ( .A1(DP_mult_98_n549), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n550), .ZN(DP_mult_98_n322) );
  XNOR2_X1 DP_mult_98_U375 ( .A(DP_sw0_2_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n548) );
  OAI22_X1 DP_mult_98_U374 ( .A1(DP_mult_98_n548), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n549), .ZN(DP_mult_98_n323) );
  XNOR2_X1 DP_mult_98_U373 ( .A(DP_sw0_1_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n547) );
  OAI22_X1 DP_mult_98_U372 ( .A1(DP_mult_98_n547), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n548), .ZN(DP_mult_98_n324) );
  XNOR2_X1 DP_mult_98_U371 ( .A(DP_sw0_0_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n544) );
  OAI22_X1 DP_mult_98_U370 ( .A1(DP_mult_98_n544), .A2(DP_mult_98_n545), .B1(
        DP_mult_98_n546), .B2(DP_mult_98_n547), .ZN(DP_mult_98_n325) );
  XOR2_X1 DP_mult_98_U369 ( .A(DP_sw0_12_), .B(DP_mult_98_n543), .Z(
        DP_mult_98_n541) );
  AOI21_X1 DP_mult_98_U368 ( .B1(DP_mult_98_n530), .B2(DP_mult_98_n532), .A(
        DP_mult_98_n541), .ZN(DP_mult_98_n542) );
  INV_X1 DP_mult_98_U367 ( .A(DP_mult_98_n542), .ZN(DP_mult_98_n327) );
  XNOR2_X1 DP_mult_98_U366 ( .A(DP_sw0_11_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n540) );
  OAI22_X1 DP_mult_98_U365 ( .A1(DP_mult_98_n540), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n541), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n328) );
  XNOR2_X1 DP_mult_98_U364 ( .A(DP_sw0_10_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n539) );
  OAI22_X1 DP_mult_98_U363 ( .A1(DP_mult_98_n539), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n540), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n329) );
  XNOR2_X1 DP_mult_98_U362 ( .A(DP_sw0_9_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n538) );
  OAI22_X1 DP_mult_98_U361 ( .A1(DP_mult_98_n538), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n539), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n330) );
  XNOR2_X1 DP_mult_98_U360 ( .A(DP_sw0_8_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n537) );
  OAI22_X1 DP_mult_98_U359 ( .A1(DP_mult_98_n537), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n538), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n331) );
  XNOR2_X1 DP_mult_98_U358 ( .A(DP_sw0_7_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n536) );
  OAI22_X1 DP_mult_98_U357 ( .A1(DP_mult_98_n536), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n537), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n332) );
  XNOR2_X1 DP_mult_98_U356 ( .A(DP_sw0_6_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n535) );
  OAI22_X1 DP_mult_98_U355 ( .A1(DP_mult_98_n535), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n536), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n333) );
  XNOR2_X1 DP_mult_98_U354 ( .A(DP_sw0_5_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n534) );
  OAI22_X1 DP_mult_98_U353 ( .A1(DP_mult_98_n534), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n535), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n334) );
  XNOR2_X1 DP_mult_98_U352 ( .A(DP_sw0_4_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n533) );
  OAI22_X1 DP_mult_98_U351 ( .A1(DP_mult_98_n533), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n534), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n335) );
  XNOR2_X1 DP_mult_98_U350 ( .A(DP_sw0_3_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n531) );
  OAI22_X1 DP_mult_98_U349 ( .A1(DP_mult_98_n531), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n533), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n336) );
  OAI22_X1 DP_mult_98_U348 ( .A1(DP_mult_98_n529), .A2(DP_mult_98_n530), .B1(
        DP_mult_98_n531), .B2(DP_mult_98_n532), .ZN(DP_mult_98_n337) );
  XNOR2_X1 DP_mult_98_U347 ( .A(DP_sw0_12_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n527) );
  OAI22_X1 DP_mult_98_U346 ( .A1(DP_mult_98_n528), .A2(DP_mult_98_n525), .B1(
        DP_mult_98_n526), .B2(DP_mult_98_n527), .ZN(DP_mult_98_n519) );
  AOI21_X1 DP_mult_98_U345 ( .B1(DP_mult_98_n525), .B2(DP_mult_98_n526), .A(
        DP_mult_98_n527), .ZN(DP_mult_98_n522) );
  INV_X1 DP_mult_98_U344 ( .A(DP_mult_98_n522), .ZN(DP_mult_98_n520) );
  INV_X1 DP_mult_98_U343 ( .A(DP_mult_98_n519), .ZN(DP_mult_98_n524) );
  AOI222_X1 DP_mult_98_U342 ( .A1(DP_mult_98_n115), .A2(DP_mult_98_n138), .B1(
        DP_mult_98_n524), .B2(DP_mult_98_n115), .C1(DP_mult_98_n524), .C2(
        DP_mult_98_n138), .ZN(DP_mult_98_n523) );
  OAI22_X1 DP_mult_98_U341 ( .A1(DP_mult_98_n522), .A2(DP_mult_98_n523), .B1(
        DP_mult_98_n524), .B2(DP_mult_98_n523), .ZN(DP_mult_98_n521) );
  AOI21_X1 DP_mult_98_U340 ( .B1(DP_mult_98_n519), .B2(DP_mult_98_n520), .A(
        DP_mult_98_n521), .ZN(DP_sw0_b1_11_) );
  XOR2_X2 DP_mult_98_U339 ( .A(DP_b_int[15]), .B(DP_mult_98_n622), .Z(
        DP_mult_98_n593) );
  XOR2_X2 DP_mult_98_U338 ( .A(DP_b_int[17]), .B(DP_mult_98_n620), .Z(
        DP_mult_98_n577) );
  XOR2_X2 DP_mult_98_U337 ( .A(DP_b_int[19]), .B(DP_mult_98_n632), .Z(
        DP_mult_98_n561) );
  XOR2_X2 DP_mult_98_U336 ( .A(DP_b_int[13]), .B(DP_mult_98_n624), .Z(
        DP_mult_98_n526) );
  INV_X1 DP_mult_98_U335 ( .A(DP_b_int[23]), .ZN(DP_mult_98_n532) );
  INV_X1 DP_mult_98_U334 ( .A(DP_mult_98_n653), .ZN(DP_mult_98_n546) );
  HA_X1 DP_mult_98_U120 ( .A(DP_mult_98_n325), .B(DP_mult_98_n337), .CO(
        DP_mult_98_n254), .S(DP_mult_98_n255) );
  FA_X1 DP_mult_98_U119 ( .A(DP_mult_98_n336), .B(DP_mult_98_n313), .CI(
        DP_mult_98_n324), .CO(DP_mult_98_n252), .S(DP_mult_98_n253) );
  HA_X1 DP_mult_98_U118 ( .A(DP_mult_98_n259), .B(DP_mult_98_n312), .CO(
        DP_mult_98_n250), .S(DP_mult_98_n251) );
  FA_X1 DP_mult_98_U117 ( .A(DP_mult_98_n323), .B(DP_mult_98_n335), .CI(
        DP_mult_98_n251), .CO(DP_mult_98_n248), .S(DP_mult_98_n249) );
  FA_X1 DP_mult_98_U109 ( .A(DP_mult_98_n334), .B(DP_mult_98_n300), .CI(
        DP_mult_98_n322), .CO(DP_mult_98_n246), .S(DP_mult_98_n247) );
  FA_X1 DP_mult_98_U108 ( .A(DP_mult_98_n250), .B(DP_mult_98_n311), .CI(
        DP_mult_98_n247), .CO(DP_mult_98_n244), .S(DP_mult_98_n245) );
  HA_X1 DP_mult_98_U107 ( .A(DP_mult_98_n258), .B(DP_mult_98_n299), .CO(
        DP_mult_98_n242), .S(DP_mult_98_n243) );
  FA_X1 DP_mult_98_U106 ( .A(DP_mult_98_n310), .B(DP_mult_98_n333), .CI(
        DP_mult_98_n321), .CO(DP_mult_98_n240), .S(DP_mult_98_n241) );
  FA_X1 DP_mult_98_U105 ( .A(DP_mult_98_n246), .B(DP_mult_98_n243), .CI(
        DP_mult_98_n241), .CO(DP_mult_98_n238), .S(DP_mult_98_n239) );
  FA_X1 DP_mult_98_U104 ( .A(DP_mult_98_n309), .B(DP_mult_98_n287), .CI(
        DP_mult_98_n332), .CO(DP_mult_98_n236), .S(DP_mult_98_n237) );
  FA_X1 DP_mult_98_U103 ( .A(DP_mult_98_n298), .B(DP_mult_98_n320), .CI(
        DP_mult_98_n242), .CO(DP_mult_98_n234), .S(DP_mult_98_n235) );
  FA_X1 DP_mult_98_U102 ( .A(DP_mult_98_n237), .B(DP_mult_98_n240), .CI(
        DP_mult_98_n235), .CO(DP_mult_98_n232), .S(DP_mult_98_n233) );
  HA_X1 DP_mult_98_U101 ( .A(DP_mult_98_n257), .B(DP_mult_98_n286), .CO(
        DP_mult_98_n230), .S(DP_mult_98_n231) );
  FA_X1 DP_mult_98_U100 ( .A(DP_mult_98_n297), .B(DP_mult_98_n308), .CI(
        DP_mult_98_n319), .CO(DP_mult_98_n228), .S(DP_mult_98_n229) );
  FA_X1 DP_mult_98_U99 ( .A(DP_mult_98_n231), .B(DP_mult_98_n331), .CI(
        DP_mult_98_n236), .CO(DP_mult_98_n226), .S(DP_mult_98_n227) );
  FA_X1 DP_mult_98_U98 ( .A(DP_mult_98_n229), .B(DP_mult_98_n234), .CI(
        DP_mult_98_n227), .CO(DP_mult_98_n224), .S(DP_mult_98_n225) );
  FA_X1 DP_mult_98_U97 ( .A(DP_mult_98_n296), .B(DP_mult_98_n274), .CI(
        DP_mult_98_n330), .CO(DP_mult_98_n222), .S(DP_mult_98_n223) );
  FA_X1 DP_mult_98_U96 ( .A(DP_mult_98_n285), .B(DP_mult_98_n318), .CI(
        DP_mult_98_n307), .CO(DP_mult_98_n220), .S(DP_mult_98_n221) );
  FA_X1 DP_mult_98_U95 ( .A(DP_mult_98_n228), .B(DP_mult_98_n230), .CI(
        DP_mult_98_n223), .CO(DP_mult_98_n218), .S(DP_mult_98_n219) );
  FA_X1 DP_mult_98_U94 ( .A(DP_mult_98_n226), .B(DP_mult_98_n221), .CI(
        DP_mult_98_n219), .CO(DP_mult_98_n216), .S(DP_mult_98_n217) );
  HA_X1 DP_mult_98_U93 ( .A(DP_mult_98_n256), .B(DP_mult_98_n273), .CO(
        DP_mult_98_n214), .S(DP_mult_98_n215) );
  FA_X1 DP_mult_98_U92 ( .A(DP_mult_98_n284), .B(DP_mult_98_n306), .CI(
        DP_mult_98_n329), .CO(DP_mult_98_n212), .S(DP_mult_98_n213) );
  FA_X1 DP_mult_98_U91 ( .A(DP_mult_98_n295), .B(DP_mult_98_n317), .CI(
        DP_mult_98_n215), .CO(DP_mult_98_n210), .S(DP_mult_98_n211) );
  FA_X1 DP_mult_98_U90 ( .A(DP_mult_98_n220), .B(DP_mult_98_n222), .CI(
        DP_mult_98_n213), .CO(DP_mult_98_n208), .S(DP_mult_98_n209) );
  FA_X1 DP_mult_98_U89 ( .A(DP_mult_98_n218), .B(DP_mult_98_n211), .CI(
        DP_mult_98_n209), .CO(DP_mult_98_n206), .S(DP_mult_98_n207) );
  HA_X1 DP_mult_98_U88 ( .A(DP_mult_98_n272), .B(DP_mult_98_n283), .CO(
        DP_mult_98_n204), .S(DP_mult_98_n205) );
  FA_X1 DP_mult_98_U87 ( .A(DP_mult_98_n328), .B(DP_mult_98_n305), .CI(
        DP_mult_98_n294), .CO(DP_mult_98_n202), .S(DP_mult_98_n203) );
  FA_X1 DP_mult_98_U86 ( .A(DP_mult_98_n214), .B(DP_mult_98_n316), .CI(
        DP_mult_98_n205), .CO(DP_mult_98_n200), .S(DP_mult_98_n201) );
  FA_X1 DP_mult_98_U85 ( .A(DP_mult_98_n203), .B(DP_mult_98_n212), .CI(
        DP_mult_98_n210), .CO(DP_mult_98_n198), .S(DP_mult_98_n199) );
  FA_X1 DP_mult_98_U84 ( .A(DP_mult_98_n208), .B(DP_mult_98_n201), .CI(
        DP_mult_98_n199), .CO(DP_mult_98_n196), .S(DP_mult_98_n197) );
  FA_X1 DP_mult_98_U81 ( .A(DP_mult_98_n271), .B(DP_mult_98_n293), .CI(
        DP_mult_98_n327), .CO(DP_mult_98_n192), .S(DP_mult_98_n193) );
  FA_X1 DP_mult_98_U80 ( .A(DP_mult_98_n204), .B(DP_mult_98_n315), .CI(
        DP_mult_98_n195), .CO(DP_mult_98_n190), .S(DP_mult_98_n191) );
  FA_X1 DP_mult_98_U79 ( .A(DP_mult_98_n193), .B(DP_mult_98_n202), .CI(
        DP_mult_98_n200), .CO(DP_mult_98_n188), .S(DP_mult_98_n189) );
  FA_X1 DP_mult_98_U78 ( .A(DP_mult_98_n198), .B(DP_mult_98_n191), .CI(
        DP_mult_98_n189), .CO(DP_mult_98_n186), .S(DP_mult_98_n187) );
  FA_X1 DP_mult_98_U76 ( .A(DP_mult_98_n303), .B(DP_mult_98_n281), .CI(
        DP_mult_98_n185), .CO(DP_mult_98_n182), .S(DP_mult_98_n183) );
  FA_X1 DP_mult_98_U75 ( .A(DP_mult_98_n270), .B(DP_mult_98_n292), .CI(
        DP_mult_98_n194), .CO(DP_mult_98_n180), .S(DP_mult_98_n181) );
  FA_X1 DP_mult_98_U74 ( .A(DP_mult_98_n190), .B(DP_mult_98_n192), .CI(
        DP_mult_98_n183), .CO(DP_mult_98_n178), .S(DP_mult_98_n179) );
  FA_X1 DP_mult_98_U73 ( .A(DP_mult_98_n188), .B(DP_mult_98_n181), .CI(
        DP_mult_98_n179), .CO(DP_mult_98_n176), .S(DP_mult_98_n177) );
  FA_X1 DP_mult_98_U72 ( .A(DP_mult_98_n184), .B(DP_mult_98_n269), .CI(
        DP_mult_98_n314), .CO(DP_mult_98_n174), .S(DP_mult_98_n175) );
  FA_X1 DP_mult_98_U71 ( .A(DP_mult_98_n280), .B(DP_mult_98_n302), .CI(
        DP_mult_98_n291), .CO(DP_mult_98_n172), .S(DP_mult_98_n173) );
  FA_X1 DP_mult_98_U70 ( .A(DP_mult_98_n180), .B(DP_mult_98_n182), .CI(
        DP_mult_98_n173), .CO(DP_mult_98_n170), .S(DP_mult_98_n171) );
  FA_X1 DP_mult_98_U69 ( .A(DP_mult_98_n178), .B(DP_mult_98_n175), .CI(
        DP_mult_98_n171), .CO(DP_mult_98_n168), .S(DP_mult_98_n169) );
  FA_X1 DP_mult_98_U67 ( .A(DP_mult_98_n268), .B(DP_mult_98_n279), .CI(
        DP_mult_98_n167), .CO(DP_mult_98_n164), .S(DP_mult_98_n165) );
  FA_X1 DP_mult_98_U66 ( .A(DP_mult_98_n174), .B(DP_mult_98_n290), .CI(
        DP_mult_98_n172), .CO(DP_mult_98_n162), .S(DP_mult_98_n163) );
  FA_X1 DP_mult_98_U65 ( .A(DP_mult_98_n170), .B(DP_mult_98_n165), .CI(
        DP_mult_98_n163), .CO(DP_mult_98_n160), .S(DP_mult_98_n161) );
  FA_X1 DP_mult_98_U64 ( .A(DP_mult_98_n166), .B(DP_mult_98_n267), .CI(
        DP_mult_98_n301), .CO(DP_mult_98_n158), .S(DP_mult_98_n159) );
  FA_X1 DP_mult_98_U63 ( .A(DP_mult_98_n278), .B(DP_mult_98_n289), .CI(
        DP_mult_98_n164), .CO(DP_mult_98_n156), .S(DP_mult_98_n157) );
  FA_X1 DP_mult_98_U62 ( .A(DP_mult_98_n162), .B(DP_mult_98_n159), .CI(
        DP_mult_98_n157), .CO(DP_mult_98_n154), .S(DP_mult_98_n155) );
  FA_X1 DP_mult_98_U60 ( .A(DP_mult_98_n266), .B(DP_mult_98_n277), .CI(
        DP_mult_98_n153), .CO(DP_mult_98_n150), .S(DP_mult_98_n151) );
  FA_X1 DP_mult_98_U59 ( .A(DP_mult_98_n151), .B(DP_mult_98_n158), .CI(
        DP_mult_98_n156), .CO(DP_mult_98_n148), .S(DP_mult_98_n149) );
  FA_X1 DP_mult_98_U58 ( .A(DP_mult_98_n265), .B(DP_mult_98_n152), .CI(
        DP_mult_98_n288), .CO(DP_mult_98_n146), .S(DP_mult_98_n147) );
  FA_X1 DP_mult_98_U57 ( .A(DP_mult_98_n150), .B(DP_mult_98_n276), .CI(
        DP_mult_98_n147), .CO(DP_mult_98_n144), .S(DP_mult_98_n145) );
  FA_X1 DP_mult_98_U55 ( .A(DP_mult_98_n143), .B(DP_mult_98_n264), .CI(
        DP_mult_98_n146), .CO(DP_mult_98_n140), .S(DP_mult_98_n141) );
  FA_X1 DP_mult_98_U54 ( .A(DP_mult_98_n263), .B(DP_mult_98_n142), .CI(
        DP_mult_98_n275), .CO(DP_mult_98_n138), .S(DP_mult_98_n139) );
  FA_X1 DP_mult_98_U42 ( .A(DP_mult_98_n207), .B(DP_mult_98_n216), .CI(
        DP_mult_98_n126), .CO(DP_mult_98_n125), .S(DP_sw0_b1_0_) );
  FA_X1 DP_mult_98_U41 ( .A(DP_mult_98_n197), .B(DP_mult_98_n206), .CI(
        DP_mult_98_n125), .CO(DP_mult_98_n124), .S(DP_sw0_b1_1_) );
  FA_X1 DP_mult_98_U40 ( .A(DP_mult_98_n187), .B(DP_mult_98_n196), .CI(
        DP_mult_98_n124), .CO(DP_mult_98_n123), .S(DP_sw0_b1_2_) );
  FA_X1 DP_mult_98_U39 ( .A(DP_mult_98_n177), .B(DP_mult_98_n186), .CI(
        DP_mult_98_n123), .CO(DP_mult_98_n122), .S(DP_sw0_b1_3_) );
  FA_X1 DP_mult_98_U38 ( .A(DP_mult_98_n169), .B(DP_mult_98_n176), .CI(
        DP_mult_98_n122), .CO(DP_mult_98_n121), .S(DP_sw0_b1_4_) );
  FA_X1 DP_mult_98_U37 ( .A(DP_mult_98_n161), .B(DP_mult_98_n168), .CI(
        DP_mult_98_n121), .CO(DP_mult_98_n120), .S(DP_sw0_b1_5_) );
  FA_X1 DP_mult_98_U36 ( .A(DP_mult_98_n155), .B(DP_mult_98_n160), .CI(
        DP_mult_98_n120), .CO(DP_mult_98_n119), .S(DP_sw0_b1_6_) );
  FA_X1 DP_mult_98_U30 ( .A(DP_mult_98_n149), .B(DP_mult_98_n154), .CI(
        DP_mult_98_n119), .CO(DP_mult_98_n118), .S(DP_sw0_b1_7_) );
  FA_X1 DP_mult_98_U20 ( .A(DP_mult_98_n145), .B(DP_mult_98_n148), .CI(
        DP_mult_98_n118), .CO(DP_mult_98_n117), .S(DP_sw0_b1_8_) );
  FA_X1 DP_mult_98_U10 ( .A(DP_mult_98_n141), .B(DP_mult_98_n144), .CI(
        DP_mult_98_n117), .CO(DP_mult_98_n116), .S(DP_sw0_b1_9_) );
  FA_X1 DP_mult_98_U9 ( .A(DP_mult_98_n140), .B(DP_mult_98_n139), .CI(
        DP_mult_98_n116), .CO(DP_mult_98_n115), .S(DP_sw0_b1_10_) );
  XOR2_X1 CU_U4 ( .A(vOut), .B(CU_presentState_0_), .Z(sw_out_regs_en_int) );
  XOR2_X1 CU_U3 ( .A(vIn), .B(sw_out_regs_en_int), .Z(CU_nextState_0_) );
  DFFR_X1 CU_presentState_reg_1_ ( .D(sw_out_regs_en_int), .CK(clk), .RN(rst_n), .Q(vOut) );
  DFFR_X1 CU_presentState_reg_0_ ( .D(CU_nextState_0_), .CK(clk), .RN(rst_n), 
        .Q(CU_presentState_0_) );
endmodule

