
module iir_filter_DW01_add_3 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   B_0_, carry_23_, carry_22_, carry_21_, carry_20_, carry_19_,
         carry_18_, carry_17_, carry_16_, carry_15_, carry_14_, carry_13_,
         carry_12_, carry_11_, carry_10_, carry_9_, carry_8_, carry_7_,
         carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, carry_1_, B_not_23_,
         B_not_22_, B_not_21_, B_not_20_, B_not_19_, B_not_18_, B_not_17_,
         B_not_16_, B_not_15_, B_not_14_, B_not_13_, B_not_12_, B_not_11_,
         B_not_10_, B_not_9_, B_not_8_, B_not_7_, B_not_6_, B_not_5_, B_not_4_,
         B_not_3_, B_not_2_, B_not_1_;
  assign DIFF[0] = B_0_;
  assign B_0_ = B[0];

  FA_X1 U2_23 ( .A(A[23]), .B(B_not_23_), .CI(carry_23_), .S(DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(B_not_22_), .CI(carry_22_), .CO(carry_23_), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(B_not_21_), .CI(carry_21_), .CO(carry_22_), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(B_not_20_), .CI(carry_20_), .CO(carry_21_), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(B_not_19_), .CI(carry_19_), .CO(carry_20_), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(B_not_18_), .CI(carry_18_), .CO(carry_19_), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(B_not_17_), .CI(carry_17_), .CO(carry_18_), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(B_not_16_), .CI(carry_16_), .CO(carry_17_), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(B_not_15_), .CI(carry_15_), .CO(carry_16_), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(B_not_14_), .CI(carry_14_), .CO(carry_15_), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(B_not_13_), .CI(carry_13_), .CO(carry_14_), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(B_not_12_), .CI(carry_12_), .CO(carry_13_), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(B_not_11_), .CI(carry_11_), .CO(carry_12_), .S(
        DIFF[11]) );
  AND2_X1 U1 ( .A1(carry_10_), .A2(B_not_10_), .ZN(carry_11_) );
  XOR2_X1 U2 ( .A(B_not_10_), .B(carry_10_), .Z(DIFF[10]) );
  AND2_X1 U3 ( .A1(carry_9_), .A2(B_not_9_), .ZN(carry_10_) );
  XOR2_X1 U4 ( .A(B_not_9_), .B(carry_9_), .Z(DIFF[9]) );
  AND2_X1 U5 ( .A1(carry_8_), .A2(B_not_8_), .ZN(carry_9_) );
  XOR2_X1 U6 ( .A(B_not_8_), .B(carry_8_), .Z(DIFF[8]) );
  AND2_X1 U7 ( .A1(carry_7_), .A2(B_not_7_), .ZN(carry_8_) );
  XOR2_X1 U8 ( .A(B_not_7_), .B(carry_7_), .Z(DIFF[7]) );
  AND2_X1 U9 ( .A1(carry_6_), .A2(B_not_6_), .ZN(carry_7_) );
  XOR2_X1 U10 ( .A(B_not_6_), .B(carry_6_), .Z(DIFF[6]) );
  AND2_X1 U11 ( .A1(carry_5_), .A2(B_not_5_), .ZN(carry_6_) );
  XOR2_X1 U12 ( .A(B_not_5_), .B(carry_5_), .Z(DIFF[5]) );
  AND2_X1 U13 ( .A1(carry_4_), .A2(B_not_4_), .ZN(carry_5_) );
  XOR2_X1 U14 ( .A(B_not_4_), .B(carry_4_), .Z(DIFF[4]) );
  AND2_X1 U15 ( .A1(carry_3_), .A2(B_not_3_), .ZN(carry_4_) );
  XOR2_X1 U16 ( .A(B_not_3_), .B(carry_3_), .Z(DIFF[3]) );
  AND2_X1 U17 ( .A1(carry_2_), .A2(B_not_2_), .ZN(carry_3_) );
  XOR2_X1 U18 ( .A(B_not_2_), .B(carry_2_), .Z(DIFF[2]) );
  AND2_X1 U19 ( .A1(carry_1_), .A2(B_not_1_), .ZN(carry_2_) );
  XOR2_X1 U20 ( .A(B_not_1_), .B(carry_1_), .Z(DIFF[1]) );
  INV_X1 U21 ( .A(B_0_), .ZN(carry_1_) );
  INV_X1 U22 ( .A(B[9]), .ZN(B_not_9_) );
  INV_X1 U23 ( .A(B[8]), .ZN(B_not_8_) );
  INV_X1 U24 ( .A(B[7]), .ZN(B_not_7_) );
  INV_X1 U25 ( .A(B[6]), .ZN(B_not_6_) );
  INV_X1 U26 ( .A(B[5]), .ZN(B_not_5_) );
  INV_X1 U27 ( .A(B[4]), .ZN(B_not_4_) );
  INV_X1 U28 ( .A(B[3]), .ZN(B_not_3_) );
  INV_X1 U29 ( .A(B[2]), .ZN(B_not_2_) );
  INV_X1 U30 ( .A(B[23]), .ZN(B_not_23_) );
  INV_X1 U31 ( .A(B[22]), .ZN(B_not_22_) );
  INV_X1 U32 ( .A(B[21]), .ZN(B_not_21_) );
  INV_X1 U33 ( .A(B[20]), .ZN(B_not_20_) );
  INV_X1 U34 ( .A(B[1]), .ZN(B_not_1_) );
  INV_X1 U35 ( .A(B[19]), .ZN(B_not_19_) );
  INV_X1 U36 ( .A(B[18]), .ZN(B_not_18_) );
  INV_X1 U37 ( .A(B[17]), .ZN(B_not_17_) );
  INV_X1 U38 ( .A(B[16]), .ZN(B_not_16_) );
  INV_X1 U39 ( .A(B[15]), .ZN(B_not_15_) );
  INV_X1 U40 ( .A(B[14]), .ZN(B_not_14_) );
  INV_X1 U41 ( .A(B[13]), .ZN(B_not_13_) );
  INV_X1 U42 ( .A(B[12]), .ZN(B_not_12_) );
  INV_X1 U43 ( .A(B[11]), .ZN(B_not_11_) );
  INV_X1 U44 ( .A(B[10]), .ZN(B_not_10_) );
endmodule


module iir_filter_DW_mult_tc_5 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(product[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(product[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(product[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(product[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(product[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(product[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(product[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(product[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(product[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(product[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(product[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(product[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(product[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(product[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(product[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(product[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(product[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(product[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(product[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(product[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(product[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(product[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(product[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1598), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1600), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1602), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1604), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1606), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1608), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1610), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(b[22]), .B(n1614), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(b[21]), .B(b[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(b[20]), .B(b[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(b[19]), .B(b[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(b[18]), .B(b[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(b[17]), .B(b[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(b[16]), .B(b[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(b[15]), .B(b[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(b[14]), .B(b[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(b[13]), .B(b[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(b[12]), .B(b[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(b[11]), .B(b[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(b[10]), .B(b[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(b[9]), .B(b[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(b[8]), .B(b[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(b[7]), .B(b[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(b[6]), .B(b[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(b[5]), .B(b[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(b[4]), .B(b[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(b[3]), .B(b[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(b[2]), .B(b[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(b[1]), .B(b[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(b[0]), .B(b[1]), .CO(n727), .S(n1397) );
  INV_X1 U1137 ( .A(n1533), .ZN(n1570) );
  INV_X1 U1138 ( .A(n1536), .ZN(n1568) );
  INV_X1 U1139 ( .A(n1535), .ZN(n1561) );
  INV_X1 U1140 ( .A(n1534), .ZN(n1569) );
  BUF_X1 U1141 ( .A(n1654), .Z(n1572) );
  INV_X1 U1142 ( .A(n1546), .ZN(n1560) );
  INV_X1 U1143 ( .A(n1544), .ZN(n1558) );
  INV_X1 U1144 ( .A(n1537), .ZN(n1580) );
  INV_X1 U1145 ( .A(n1550), .ZN(n1575) );
  INV_X1 U1146 ( .A(n1549), .ZN(n1585) );
  INV_X1 U1147 ( .A(n1547), .ZN(n1595) );
  INV_X1 U1148 ( .A(n1548), .ZN(n1590) );
  INV_X1 U1149 ( .A(n1538), .ZN(n1559) );
  INV_X1 U1150 ( .A(n1545), .ZN(n1593) );
  INV_X1 U1151 ( .A(n1552), .ZN(n1583) );
  INV_X1 U1152 ( .A(n1551), .ZN(n1588) );
  INV_X1 U1153 ( .A(n1553), .ZN(n1578) );
  INV_X1 U1154 ( .A(n1554), .ZN(n1573) );
  BUF_X1 U1155 ( .A(n1654), .Z(n1571) );
  BUF_X1 U1156 ( .A(n1629), .Z(n1557) );
  BUF_X1 U1157 ( .A(n1967), .Z(n1596) );
  BUF_X1 U1158 ( .A(n1912), .Z(n1591) );
  BUF_X1 U1159 ( .A(n1857), .Z(n1586) );
  BUF_X1 U1160 ( .A(n1802), .Z(n1581) );
  BUF_X1 U1161 ( .A(n1747), .Z(n1576) );
  BUF_X1 U1162 ( .A(n1912), .Z(n1592) );
  BUF_X1 U1163 ( .A(n1857), .Z(n1587) );
  BUF_X1 U1164 ( .A(n1802), .Z(n1582) );
  BUF_X1 U1165 ( .A(n1747), .Z(n1577) );
  BUF_X1 U1166 ( .A(n1967), .Z(n1597) );
  INV_X1 U1167 ( .A(n1615), .ZN(n1614) );
  INV_X1 U1168 ( .A(n1540), .ZN(n1589) );
  INV_X1 U1169 ( .A(n1541), .ZN(n1584) );
  INV_X1 U1170 ( .A(n1542), .ZN(n1579) );
  INV_X1 U1171 ( .A(n1543), .ZN(n1574) );
  BUF_X1 U1172 ( .A(n1629), .Z(n1556) );
  INV_X1 U1173 ( .A(n1539), .ZN(n1594) );
  NAND3_X1 U1174 ( .A1(n2157), .A2(n2158), .A3(n2159), .ZN(n1639) );
  INV_X1 U1175 ( .A(n1555), .ZN(n1564) );
  OR2_X1 U1176 ( .A1(n1738), .A2(n1739), .ZN(n1533) );
  OR2_X1 U1177 ( .A1(n1740), .A2(n1741), .ZN(n1534) );
  OR2_X1 U1178 ( .A1(n2158), .A2(n2157), .ZN(n1535) );
  AND2_X1 U1179 ( .A1(n1738), .A2(n1740), .ZN(n1536) );
  INV_X1 U1180 ( .A(n1611), .ZN(n1610) );
  INV_X1 U1181 ( .A(n1607), .ZN(n1606) );
  INV_X1 U1182 ( .A(n1609), .ZN(n1608) );
  INV_X1 U1183 ( .A(n1605), .ZN(n1604) );
  INV_X1 U1184 ( .A(n1603), .ZN(n1602) );
  OR2_X1 U1185 ( .A1(n1849), .A2(n1850), .ZN(n1537) );
  BUF_X1 U1186 ( .A(n1636), .Z(n1562) );
  BUF_X1 U1187 ( .A(n1636), .Z(n1563) );
  BUF_X1 U1188 ( .A(n1647), .Z(n1565) );
  BUF_X1 U1189 ( .A(n1647), .Z(n1566) );
  OR2_X1 U1190 ( .A1(n2068), .A2(n2067), .ZN(n1538) );
  OR2_X1 U1191 ( .A1(n2016), .A2(n2017), .ZN(n1539) );
  OR2_X1 U1192 ( .A1(n1961), .A2(n1962), .ZN(n1540) );
  OR2_X1 U1193 ( .A1(n1906), .A2(n1907), .ZN(n1541) );
  OR2_X1 U1194 ( .A1(n1851), .A2(n1852), .ZN(n1542) );
  OR2_X1 U1195 ( .A1(n1796), .A2(n1797), .ZN(n1543) );
  AND2_X1 U1196 ( .A1(n2070), .A2(n2068), .ZN(n1544) );
  AND2_X1 U1197 ( .A1(n2014), .A2(n2016), .ZN(n1545) );
  OR2_X1 U1198 ( .A1(n2070), .A2(n2069), .ZN(n1546) );
  OR2_X1 U1199 ( .A1(n2014), .A2(n2015), .ZN(n1547) );
  OR2_X1 U1200 ( .A1(n1959), .A2(n1960), .ZN(n1548) );
  OR2_X1 U1201 ( .A1(n1904), .A2(n1905), .ZN(n1549) );
  OR2_X1 U1202 ( .A1(n1794), .A2(n1795), .ZN(n1550) );
  AND2_X1 U1203 ( .A1(n1959), .A2(n1961), .ZN(n1551) );
  AND2_X1 U1204 ( .A1(n1904), .A2(n1906), .ZN(n1552) );
  AND2_X1 U1205 ( .A1(n1849), .A2(n1851), .ZN(n1553) );
  AND2_X1 U1206 ( .A1(n1794), .A2(n1796), .ZN(n1554) );
  BUF_X1 U1207 ( .A(n1647), .Z(n1567) );
  INV_X1 U1208 ( .A(n1599), .ZN(n1598) );
  AND2_X1 U1209 ( .A1(a[0]), .A2(n2157), .ZN(n1555) );
  BUF_X1 U1210 ( .A(a[20]), .Z(n1600) );
  INV_X1 U1211 ( .A(a[23]), .ZN(n1599) );
  INV_X1 U1212 ( .A(a[5]), .ZN(n1611) );
  INV_X1 U1213 ( .A(a[11]), .ZN(n1607) );
  INV_X1 U1214 ( .A(a[8]), .ZN(n1609) );
  INV_X1 U1215 ( .A(a[14]), .ZN(n1605) );
  INV_X1 U1216 ( .A(a[17]), .ZN(n1603) );
  BUF_X1 U1217 ( .A(a[20]), .Z(n1601) );
  CLKBUF_X1 U1218 ( .A(b[23]), .Z(n1612) );
  CLKBUF_X1 U1219 ( .A(b[23]), .Z(n1613) );
  INV_X1 U1220 ( .A(b[23]), .ZN(n1615) );
  INV_X1 U1221 ( .A(n1612), .ZN(n1616) );
  INV_X1 U1222 ( .A(n1612), .ZN(n1617) );
  INV_X1 U1223 ( .A(n1612), .ZN(n1618) );
  INV_X1 U1224 ( .A(n1613), .ZN(n1619) );
  INV_X1 U1225 ( .A(n1613), .ZN(n1620) );
  AOI21_X1 U1226 ( .B1(n1621), .B2(n1622), .A(n1623), .ZN(product[47]) );
  OAI22_X1 U1227 ( .A1(n1624), .A2(n1625), .B1(n1624), .B2(n1626), .ZN(n1623)
         );
  INV_X1 U1228 ( .A(n1622), .ZN(n1626) );
  AOI222_X1 U1229 ( .A1(n1627), .A2(n303), .B1(n1625), .B2(n303), .C1(n1627), 
        .C2(n1625), .ZN(n1624) );
  XOR2_X1 U1230 ( .A(n1628), .B(n1599), .Z(n1622) );
  OAI221_X1 U1231 ( .B1(n1617), .B2(n1557), .C1(n1620), .C2(n1558), .A(n1630), 
        .ZN(n1628) );
  OAI21_X1 U1232 ( .B1(n1559), .B2(n1560), .A(n1614), .ZN(n1630) );
  INV_X1 U1233 ( .A(n1625), .ZN(n1621) );
  XOR2_X1 U1234 ( .A(a[23]), .B(n1631), .Z(n1625) );
  AOI221_X1 U1235 ( .B1(n1613), .B2(n1559), .C1(n1560), .C2(n1614), .A(n1632), 
        .ZN(n1631) );
  OAI22_X1 U1236 ( .A1(n1558), .A2(n1633), .B1(n1557), .B2(n1634), .ZN(n1632)
         );
  XNOR2_X1 U1237 ( .A(a[2]), .B(n1635), .ZN(n908) );
  AOI221_X1 U1238 ( .B1(n1561), .B2(b[22]), .C1(n1563), .C2(b[21]), .A(n1637), 
        .ZN(n1635) );
  OAI22_X1 U1239 ( .A1(n1564), .A2(n1638), .B1(n1639), .B2(n1640), .ZN(n1637)
         );
  INV_X1 U1240 ( .A(n1376), .ZN(n1638) );
  XNOR2_X1 U1241 ( .A(a[2]), .B(n1641), .ZN(n907) );
  AOI221_X1 U1242 ( .B1(n1563), .B2(b[22]), .C1(n1555), .C2(n1375), .A(n1642), 
        .ZN(n1641) );
  OAI22_X1 U1243 ( .A1(n1643), .A2(n1639), .B1(n1617), .B2(n1535), .ZN(n1642)
         );
  XNOR2_X1 U1244 ( .A(a[2]), .B(n1644), .ZN(n906) );
  AOI221_X1 U1245 ( .B1(n1561), .B2(n1613), .C1(n1563), .C2(n1614), .A(n1645), 
        .ZN(n1644) );
  OAI22_X1 U1246 ( .A1(n1633), .A2(n1564), .B1(n1634), .B2(n1639), .ZN(n1645)
         );
  XNOR2_X1 U1247 ( .A(n1646), .B(n1611), .ZN(n904) );
  OAI22_X1 U1248 ( .A1(n1565), .A2(n1534), .B1(n1568), .B2(n1567), .ZN(n1646)
         );
  XNOR2_X1 U1249 ( .A(n1648), .B(n1611), .ZN(n903) );
  OAI222_X1 U1250 ( .A1(n1534), .A2(n1649), .B1(n1566), .B2(n1533), .C1(n1568), 
        .C2(n1650), .ZN(n1648) );
  XNOR2_X1 U1251 ( .A(n1610), .B(n1651), .ZN(n902) );
  AOI221_X1 U1252 ( .B1(b[2]), .B2(n1569), .C1(b[1]), .C2(n1570), .A(n1652), 
        .ZN(n1651) );
  OAI22_X1 U1253 ( .A1(n1568), .A2(n1653), .B1(n1565), .B2(n1572), .ZN(n1652)
         );
  XNOR2_X1 U1254 ( .A(n1610), .B(n1655), .ZN(n901) );
  AOI221_X1 U1255 ( .B1(b[3]), .B2(n1569), .C1(b[2]), .C2(n1570), .A(n1656), 
        .ZN(n1655) );
  OAI22_X1 U1256 ( .A1(n1568), .A2(n1657), .B1(n1649), .B2(n1572), .ZN(n1656)
         );
  XNOR2_X1 U1257 ( .A(n1610), .B(n1658), .ZN(n900) );
  AOI221_X1 U1258 ( .B1(b[4]), .B2(n1569), .C1(b[3]), .C2(n1570), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1259 ( .A1(n1568), .A2(n1660), .B1(n1661), .B2(n1572), .ZN(n1659)
         );
  XNOR2_X1 U1260 ( .A(n1610), .B(n1662), .ZN(n899) );
  AOI221_X1 U1261 ( .B1(b[5]), .B2(n1569), .C1(b[4]), .C2(n1570), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1262 ( .A1(n1568), .A2(n1664), .B1(n1572), .B2(n1665), .ZN(n1663)
         );
  XNOR2_X1 U1263 ( .A(n1610), .B(n1666), .ZN(n898) );
  AOI221_X1 U1264 ( .B1(b[6]), .B2(n1569), .C1(b[5]), .C2(n1570), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1265 ( .A1(n1568), .A2(n1668), .B1(n1572), .B2(n1669), .ZN(n1667)
         );
  XNOR2_X1 U1266 ( .A(n1610), .B(n1670), .ZN(n897) );
  AOI221_X1 U1267 ( .B1(b[7]), .B2(n1569), .C1(b[6]), .C2(n1570), .A(n1671), 
        .ZN(n1670) );
  OAI22_X1 U1268 ( .A1(n1568), .A2(n1672), .B1(n1572), .B2(n1673), .ZN(n1671)
         );
  XNOR2_X1 U1269 ( .A(n1610), .B(n1674), .ZN(n896) );
  AOI221_X1 U1270 ( .B1(b[8]), .B2(n1569), .C1(b[7]), .C2(n1570), .A(n1675), 
        .ZN(n1674) );
  OAI22_X1 U1271 ( .A1(n1568), .A2(n1676), .B1(n1571), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1272 ( .A(n1610), .B(n1678), .ZN(n895) );
  AOI221_X1 U1273 ( .B1(b[9]), .B2(n1569), .C1(b[8]), .C2(n1570), .A(n1679), 
        .ZN(n1678) );
  OAI22_X1 U1274 ( .A1(n1568), .A2(n1680), .B1(n1572), .B2(n1681), .ZN(n1679)
         );
  XNOR2_X1 U1275 ( .A(n1610), .B(n1682), .ZN(n894) );
  AOI221_X1 U1276 ( .B1(b[10]), .B2(n1569), .C1(b[9]), .C2(n1570), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1277 ( .A1(n1568), .A2(n1684), .B1(n1572), .B2(n1685), .ZN(n1683)
         );
  XNOR2_X1 U1278 ( .A(n1610), .B(n1686), .ZN(n893) );
  AOI221_X1 U1279 ( .B1(b[11]), .B2(n1569), .C1(b[10]), .C2(n1570), .A(n1687), 
        .ZN(n1686) );
  OAI22_X1 U1280 ( .A1(n1568), .A2(n1688), .B1(n1571), .B2(n1689), .ZN(n1687)
         );
  XNOR2_X1 U1281 ( .A(n1610), .B(n1690), .ZN(n892) );
  AOI221_X1 U1282 ( .B1(b[12]), .B2(n1569), .C1(b[11]), .C2(n1570), .A(n1691), 
        .ZN(n1690) );
  OAI22_X1 U1283 ( .A1(n1568), .A2(n1692), .B1(n1571), .B2(n1693), .ZN(n1691)
         );
  XNOR2_X1 U1284 ( .A(n1610), .B(n1694), .ZN(n891) );
  AOI221_X1 U1285 ( .B1(b[13]), .B2(n1569), .C1(b[12]), .C2(n1570), .A(n1695), 
        .ZN(n1694) );
  OAI22_X1 U1286 ( .A1(n1568), .A2(n1696), .B1(n1571), .B2(n1697), .ZN(n1695)
         );
  XNOR2_X1 U1287 ( .A(n1610), .B(n1698), .ZN(n890) );
  AOI221_X1 U1288 ( .B1(b[14]), .B2(n1569), .C1(b[13]), .C2(n1570), .A(n1699), 
        .ZN(n1698) );
  OAI22_X1 U1289 ( .A1(n1568), .A2(n1700), .B1(n1571), .B2(n1701), .ZN(n1699)
         );
  XNOR2_X1 U1290 ( .A(n1610), .B(n1702), .ZN(n889) );
  AOI221_X1 U1291 ( .B1(b[15]), .B2(n1569), .C1(b[14]), .C2(n1570), .A(n1703), 
        .ZN(n1702) );
  OAI22_X1 U1292 ( .A1(n1568), .A2(n1704), .B1(n1571), .B2(n1705), .ZN(n1703)
         );
  XNOR2_X1 U1293 ( .A(n1610), .B(n1706), .ZN(n888) );
  AOI221_X1 U1294 ( .B1(b[16]), .B2(n1569), .C1(b[15]), .C2(n1570), .A(n1707), 
        .ZN(n1706) );
  OAI22_X1 U1295 ( .A1(n1568), .A2(n1708), .B1(n1571), .B2(n1709), .ZN(n1707)
         );
  XNOR2_X1 U1296 ( .A(n1610), .B(n1710), .ZN(n887) );
  AOI221_X1 U1297 ( .B1(b[17]), .B2(n1569), .C1(b[16]), .C2(n1570), .A(n1711), 
        .ZN(n1710) );
  OAI22_X1 U1298 ( .A1(n1568), .A2(n1712), .B1(n1571), .B2(n1713), .ZN(n1711)
         );
  XNOR2_X1 U1299 ( .A(n1610), .B(n1714), .ZN(n886) );
  AOI221_X1 U1300 ( .B1(b[18]), .B2(n1569), .C1(b[17]), .C2(n1570), .A(n1715), 
        .ZN(n1714) );
  OAI22_X1 U1301 ( .A1(n1568), .A2(n1716), .B1(n1571), .B2(n1717), .ZN(n1715)
         );
  XNOR2_X1 U1302 ( .A(n1610), .B(n1718), .ZN(n885) );
  AOI221_X1 U1303 ( .B1(b[19]), .B2(n1569), .C1(b[18]), .C2(n1570), .A(n1719), 
        .ZN(n1718) );
  OAI22_X1 U1304 ( .A1(n1568), .A2(n1720), .B1(n1571), .B2(n1721), .ZN(n1719)
         );
  XNOR2_X1 U1305 ( .A(a[5]), .B(n1722), .ZN(n884) );
  AOI221_X1 U1306 ( .B1(n1569), .B2(b[20]), .C1(b[19]), .C2(n1570), .A(n1723), 
        .ZN(n1722) );
  OAI22_X1 U1307 ( .A1(n1568), .A2(n1724), .B1(n1571), .B2(n1725), .ZN(n1723)
         );
  XNOR2_X1 U1308 ( .A(a[5]), .B(n1726), .ZN(n883) );
  AOI221_X1 U1309 ( .B1(n1569), .B2(b[21]), .C1(n1570), .C2(b[20]), .A(n1727), 
        .ZN(n1726) );
  OAI22_X1 U1310 ( .A1(n1568), .A2(n1728), .B1(n1571), .B2(n1729), .ZN(n1727)
         );
  XNOR2_X1 U1311 ( .A(a[5]), .B(n1730), .ZN(n882) );
  AOI221_X1 U1312 ( .B1(n1569), .B2(b[22]), .C1(n1536), .C2(n1376), .A(n1731), 
        .ZN(n1730) );
  OAI22_X1 U1313 ( .A1(n1640), .A2(n1572), .B1(n1643), .B2(n1533), .ZN(n1731)
         );
  XNOR2_X1 U1314 ( .A(a[5]), .B(n1732), .ZN(n881) );
  AOI221_X1 U1315 ( .B1(n1570), .B2(b[22]), .C1(n1536), .C2(n1375), .A(n1733), 
        .ZN(n1732) );
  OAI22_X1 U1316 ( .A1(n1615), .A2(n1534), .B1(n1643), .B2(n1572), .ZN(n1733)
         );
  XNOR2_X1 U1317 ( .A(a[5]), .B(n1734), .ZN(n880) );
  AOI221_X1 U1318 ( .B1(n1569), .B2(n1613), .C1(n1570), .C2(n1614), .A(n1735), 
        .ZN(n1734) );
  OAI22_X1 U1319 ( .A1(n1633), .A2(n1568), .B1(n1634), .B2(n1572), .ZN(n1735)
         );
  XNOR2_X1 U1320 ( .A(n1610), .B(n1736), .ZN(n879) );
  OAI221_X1 U1321 ( .B1(n1616), .B2(n1572), .C1(n1620), .C2(n1568), .A(n1737), 
        .ZN(n1736) );
  OAI21_X1 U1322 ( .B1(n1569), .B2(n1570), .A(n1614), .ZN(n1737) );
  INV_X1 U1323 ( .A(n1741), .ZN(n1738) );
  NAND3_X1 U1324 ( .A1(n1741), .A2(n1740), .A3(n1739), .ZN(n1654) );
  XNOR2_X1 U1325 ( .A(a[3]), .B(a[4]), .ZN(n1739) );
  XNOR2_X1 U1326 ( .A(a[4]), .B(n1611), .ZN(n1740) );
  XOR2_X1 U1327 ( .A(a[3]), .B(n1742), .Z(n1741) );
  XNOR2_X1 U1328 ( .A(n1743), .B(n1609), .ZN(n878) );
  OAI22_X1 U1329 ( .A1(n1565), .A2(n1543), .B1(n1565), .B2(n1573), .ZN(n1743)
         );
  XNOR2_X1 U1330 ( .A(n1744), .B(n1609), .ZN(n877) );
  OAI222_X1 U1331 ( .A1(n1649), .A2(n1543), .B1(n1566), .B2(n1550), .C1(n1650), 
        .C2(n1573), .ZN(n1744) );
  XNOR2_X1 U1332 ( .A(n1608), .B(n1745), .ZN(n876) );
  AOI221_X1 U1333 ( .B1(n1574), .B2(b[2]), .C1(n1575), .C2(b[1]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1334 ( .A1(n1653), .A2(n1573), .B1(n1565), .B2(n1576), .ZN(n1746)
         );
  XNOR2_X1 U1335 ( .A(n1608), .B(n1748), .ZN(n875) );
  AOI221_X1 U1336 ( .B1(n1574), .B2(b[3]), .C1(n1575), .C2(b[2]), .A(n1749), 
        .ZN(n1748) );
  OAI22_X1 U1337 ( .A1(n1657), .A2(n1573), .B1(n1649), .B2(n1577), .ZN(n1749)
         );
  XNOR2_X1 U1338 ( .A(n1608), .B(n1750), .ZN(n874) );
  AOI221_X1 U1339 ( .B1(n1574), .B2(b[4]), .C1(n1575), .C2(b[3]), .A(n1751), 
        .ZN(n1750) );
  OAI22_X1 U1340 ( .A1(n1660), .A2(n1573), .B1(n1661), .B2(n1577), .ZN(n1751)
         );
  XNOR2_X1 U1341 ( .A(n1608), .B(n1752), .ZN(n873) );
  AOI221_X1 U1342 ( .B1(n1574), .B2(b[5]), .C1(n1575), .C2(b[4]), .A(n1753), 
        .ZN(n1752) );
  OAI22_X1 U1343 ( .A1(n1664), .A2(n1573), .B1(n1665), .B2(n1577), .ZN(n1753)
         );
  XNOR2_X1 U1344 ( .A(n1608), .B(n1754), .ZN(n872) );
  AOI221_X1 U1345 ( .B1(n1574), .B2(b[6]), .C1(n1575), .C2(b[5]), .A(n1755), 
        .ZN(n1754) );
  OAI22_X1 U1346 ( .A1(n1668), .A2(n1573), .B1(n1669), .B2(n1577), .ZN(n1755)
         );
  XNOR2_X1 U1347 ( .A(n1608), .B(n1756), .ZN(n871) );
  AOI221_X1 U1348 ( .B1(n1574), .B2(b[7]), .C1(n1575), .C2(b[6]), .A(n1757), 
        .ZN(n1756) );
  OAI22_X1 U1349 ( .A1(n1672), .A2(n1573), .B1(n1673), .B2(n1577), .ZN(n1757)
         );
  XNOR2_X1 U1350 ( .A(n1608), .B(n1758), .ZN(n870) );
  AOI221_X1 U1351 ( .B1(n1574), .B2(b[8]), .C1(n1575), .C2(b[7]), .A(n1759), 
        .ZN(n1758) );
  OAI22_X1 U1352 ( .A1(n1676), .A2(n1573), .B1(n1677), .B2(n1577), .ZN(n1759)
         );
  XNOR2_X1 U1353 ( .A(n1608), .B(n1760), .ZN(n869) );
  AOI221_X1 U1354 ( .B1(n1574), .B2(b[9]), .C1(n1575), .C2(b[8]), .A(n1761), 
        .ZN(n1760) );
  OAI22_X1 U1355 ( .A1(n1680), .A2(n1573), .B1(n1681), .B2(n1577), .ZN(n1761)
         );
  XNOR2_X1 U1356 ( .A(n1608), .B(n1762), .ZN(n868) );
  AOI221_X1 U1357 ( .B1(n1574), .B2(b[10]), .C1(n1575), .C2(b[9]), .A(n1763), 
        .ZN(n1762) );
  OAI22_X1 U1358 ( .A1(n1684), .A2(n1573), .B1(n1685), .B2(n1577), .ZN(n1763)
         );
  XNOR2_X1 U1359 ( .A(n1608), .B(n1764), .ZN(n867) );
  AOI221_X1 U1360 ( .B1(n1574), .B2(b[11]), .C1(n1575), .C2(b[10]), .A(n1765), 
        .ZN(n1764) );
  OAI22_X1 U1361 ( .A1(n1688), .A2(n1573), .B1(n1689), .B2(n1577), .ZN(n1765)
         );
  XNOR2_X1 U1362 ( .A(n1608), .B(n1766), .ZN(n866) );
  AOI221_X1 U1363 ( .B1(n1574), .B2(b[12]), .C1(n1575), .C2(b[11]), .A(n1767), 
        .ZN(n1766) );
  OAI22_X1 U1364 ( .A1(n1692), .A2(n1573), .B1(n1693), .B2(n1577), .ZN(n1767)
         );
  XNOR2_X1 U1365 ( .A(n1608), .B(n1768), .ZN(n865) );
  AOI221_X1 U1366 ( .B1(n1574), .B2(b[13]), .C1(n1575), .C2(b[12]), .A(n1769), 
        .ZN(n1768) );
  OAI22_X1 U1367 ( .A1(n1696), .A2(n1573), .B1(n1697), .B2(n1576), .ZN(n1769)
         );
  XNOR2_X1 U1368 ( .A(n1608), .B(n1770), .ZN(n864) );
  AOI221_X1 U1369 ( .B1(n1574), .B2(b[14]), .C1(n1575), .C2(b[13]), .A(n1771), 
        .ZN(n1770) );
  OAI22_X1 U1370 ( .A1(n1700), .A2(n1573), .B1(n1701), .B2(n1576), .ZN(n1771)
         );
  XNOR2_X1 U1371 ( .A(n1608), .B(n1772), .ZN(n863) );
  AOI221_X1 U1372 ( .B1(n1574), .B2(b[15]), .C1(n1575), .C2(b[14]), .A(n1773), 
        .ZN(n1772) );
  OAI22_X1 U1373 ( .A1(n1704), .A2(n1573), .B1(n1705), .B2(n1576), .ZN(n1773)
         );
  XNOR2_X1 U1374 ( .A(n1608), .B(n1774), .ZN(n862) );
  AOI221_X1 U1375 ( .B1(n1574), .B2(b[16]), .C1(n1575), .C2(b[15]), .A(n1775), 
        .ZN(n1774) );
  OAI22_X1 U1376 ( .A1(n1708), .A2(n1573), .B1(n1709), .B2(n1576), .ZN(n1775)
         );
  XNOR2_X1 U1377 ( .A(n1608), .B(n1776), .ZN(n861) );
  AOI221_X1 U1378 ( .B1(n1574), .B2(b[17]), .C1(n1575), .C2(b[16]), .A(n1777), 
        .ZN(n1776) );
  OAI22_X1 U1379 ( .A1(n1712), .A2(n1573), .B1(n1713), .B2(n1576), .ZN(n1777)
         );
  XNOR2_X1 U1380 ( .A(n1608), .B(n1778), .ZN(n860) );
  AOI221_X1 U1381 ( .B1(n1574), .B2(b[18]), .C1(n1575), .C2(b[17]), .A(n1779), 
        .ZN(n1778) );
  OAI22_X1 U1382 ( .A1(n1716), .A2(n1573), .B1(n1717), .B2(n1576), .ZN(n1779)
         );
  XNOR2_X1 U1383 ( .A(n1608), .B(n1780), .ZN(n859) );
  AOI221_X1 U1384 ( .B1(n1574), .B2(b[19]), .C1(n1575), .C2(b[18]), .A(n1781), 
        .ZN(n1780) );
  OAI22_X1 U1385 ( .A1(n1720), .A2(n1573), .B1(n1721), .B2(n1576), .ZN(n1781)
         );
  XNOR2_X1 U1386 ( .A(a[8]), .B(n1782), .ZN(n858) );
  AOI221_X1 U1387 ( .B1(n1574), .B2(b[20]), .C1(n1575), .C2(b[19]), .A(n1783), 
        .ZN(n1782) );
  OAI22_X1 U1388 ( .A1(n1724), .A2(n1573), .B1(n1725), .B2(n1576), .ZN(n1783)
         );
  XNOR2_X1 U1389 ( .A(a[8]), .B(n1784), .ZN(n857) );
  AOI221_X1 U1390 ( .B1(n1574), .B2(b[21]), .C1(n1575), .C2(b[20]), .A(n1785), 
        .ZN(n1784) );
  OAI22_X1 U1391 ( .A1(n1728), .A2(n1573), .B1(n1729), .B2(n1576), .ZN(n1785)
         );
  XNOR2_X1 U1392 ( .A(a[8]), .B(n1786), .ZN(n856) );
  AOI221_X1 U1393 ( .B1(n1574), .B2(b[22]), .C1(n1554), .C2(n1376), .A(n1787), 
        .ZN(n1786) );
  OAI22_X1 U1394 ( .A1(n1640), .A2(n1577), .B1(n1643), .B2(n1550), .ZN(n1787)
         );
  XNOR2_X1 U1395 ( .A(a[8]), .B(n1788), .ZN(n855) );
  AOI221_X1 U1396 ( .B1(n1575), .B2(b[22]), .C1(n1554), .C2(n1375), .A(n1789), 
        .ZN(n1788) );
  OAI22_X1 U1397 ( .A1(n1617), .A2(n1543), .B1(n1643), .B2(n1576), .ZN(n1789)
         );
  XNOR2_X1 U1398 ( .A(a[8]), .B(n1790), .ZN(n854) );
  AOI221_X1 U1399 ( .B1(n1574), .B2(n1613), .C1(n1575), .C2(n1614), .A(n1791), 
        .ZN(n1790) );
  OAI22_X1 U1400 ( .A1(n1633), .A2(n1573), .B1(n1634), .B2(n1576), .ZN(n1791)
         );
  XNOR2_X1 U1401 ( .A(n1608), .B(n1792), .ZN(n853) );
  OAI221_X1 U1402 ( .B1(n1616), .B2(n1577), .C1(n1617), .C2(n1573), .A(n1793), 
        .ZN(n1792) );
  OAI21_X1 U1403 ( .B1(n1574), .B2(n1575), .A(n1614), .ZN(n1793) );
  INV_X1 U1404 ( .A(n1797), .ZN(n1794) );
  NAND3_X1 U1405 ( .A1(n1797), .A2(n1796), .A3(n1795), .ZN(n1747) );
  XNOR2_X1 U1406 ( .A(a[6]), .B(a[7]), .ZN(n1795) );
  XNOR2_X1 U1407 ( .A(a[7]), .B(n1609), .ZN(n1796) );
  XOR2_X1 U1408 ( .A(a[6]), .B(n1611), .Z(n1797) );
  XNOR2_X1 U1409 ( .A(n1798), .B(n1607), .ZN(n852) );
  OAI22_X1 U1410 ( .A1(n1565), .A2(n1542), .B1(n1565), .B2(n1578), .ZN(n1798)
         );
  XNOR2_X1 U1411 ( .A(n1799), .B(n1607), .ZN(n851) );
  OAI222_X1 U1412 ( .A1(n1649), .A2(n1542), .B1(n1566), .B2(n1537), .C1(n1650), 
        .C2(n1578), .ZN(n1799) );
  XNOR2_X1 U1413 ( .A(n1606), .B(n1800), .ZN(n850) );
  AOI221_X1 U1414 ( .B1(n1579), .B2(b[2]), .C1(n1580), .C2(b[1]), .A(n1801), 
        .ZN(n1800) );
  OAI22_X1 U1415 ( .A1(n1653), .A2(n1578), .B1(n1566), .B2(n1581), .ZN(n1801)
         );
  XNOR2_X1 U1416 ( .A(n1606), .B(n1803), .ZN(n849) );
  AOI221_X1 U1417 ( .B1(n1579), .B2(b[3]), .C1(n1580), .C2(b[2]), .A(n1804), 
        .ZN(n1803) );
  OAI22_X1 U1418 ( .A1(n1657), .A2(n1578), .B1(n1649), .B2(n1582), .ZN(n1804)
         );
  XNOR2_X1 U1419 ( .A(n1606), .B(n1805), .ZN(n848) );
  AOI221_X1 U1420 ( .B1(n1579), .B2(b[4]), .C1(n1580), .C2(b[3]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1421 ( .A1(n1660), .A2(n1578), .B1(n1661), .B2(n1582), .ZN(n1806)
         );
  XNOR2_X1 U1422 ( .A(n1606), .B(n1807), .ZN(n847) );
  AOI221_X1 U1423 ( .B1(n1579), .B2(b[5]), .C1(n1580), .C2(b[4]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1424 ( .A1(n1664), .A2(n1578), .B1(n1665), .B2(n1582), .ZN(n1808)
         );
  XNOR2_X1 U1425 ( .A(n1606), .B(n1809), .ZN(n846) );
  AOI221_X1 U1426 ( .B1(n1579), .B2(b[6]), .C1(n1580), .C2(b[5]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1427 ( .A1(n1668), .A2(n1578), .B1(n1669), .B2(n1582), .ZN(n1810)
         );
  XNOR2_X1 U1428 ( .A(n1606), .B(n1811), .ZN(n845) );
  AOI221_X1 U1429 ( .B1(n1579), .B2(b[7]), .C1(n1580), .C2(b[6]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1430 ( .A1(n1672), .A2(n1578), .B1(n1673), .B2(n1582), .ZN(n1812)
         );
  XNOR2_X1 U1431 ( .A(n1606), .B(n1813), .ZN(n844) );
  AOI221_X1 U1432 ( .B1(n1579), .B2(b[8]), .C1(n1580), .C2(b[7]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1433 ( .A1(n1676), .A2(n1578), .B1(n1677), .B2(n1582), .ZN(n1814)
         );
  XNOR2_X1 U1434 ( .A(n1606), .B(n1815), .ZN(n843) );
  AOI221_X1 U1435 ( .B1(n1579), .B2(b[9]), .C1(n1580), .C2(b[8]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1436 ( .A1(n1680), .A2(n1578), .B1(n1681), .B2(n1582), .ZN(n1816)
         );
  XNOR2_X1 U1437 ( .A(n1606), .B(n1817), .ZN(n842) );
  AOI221_X1 U1438 ( .B1(n1579), .B2(b[10]), .C1(n1580), .C2(b[9]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1439 ( .A1(n1684), .A2(n1578), .B1(n1685), .B2(n1582), .ZN(n1818)
         );
  XNOR2_X1 U1440 ( .A(n1606), .B(n1819), .ZN(n841) );
  AOI221_X1 U1441 ( .B1(n1579), .B2(b[11]), .C1(n1580), .C2(b[10]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1442 ( .A1(n1688), .A2(n1578), .B1(n1689), .B2(n1582), .ZN(n1820)
         );
  XNOR2_X1 U1443 ( .A(n1606), .B(n1821), .ZN(n840) );
  AOI221_X1 U1444 ( .B1(n1579), .B2(b[12]), .C1(n1580), .C2(b[11]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1445 ( .A1(n1692), .A2(n1578), .B1(n1693), .B2(n1582), .ZN(n1822)
         );
  XNOR2_X1 U1446 ( .A(n1606), .B(n1823), .ZN(n839) );
  AOI221_X1 U1447 ( .B1(n1579), .B2(b[13]), .C1(n1580), .C2(b[12]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1448 ( .A1(n1696), .A2(n1578), .B1(n1697), .B2(n1581), .ZN(n1824)
         );
  XNOR2_X1 U1449 ( .A(n1606), .B(n1825), .ZN(n838) );
  AOI221_X1 U1450 ( .B1(n1579), .B2(b[14]), .C1(n1580), .C2(b[13]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1451 ( .A1(n1700), .A2(n1578), .B1(n1701), .B2(n1581), .ZN(n1826)
         );
  XNOR2_X1 U1452 ( .A(n1606), .B(n1827), .ZN(n837) );
  AOI221_X1 U1453 ( .B1(n1579), .B2(b[15]), .C1(n1580), .C2(b[14]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1454 ( .A1(n1704), .A2(n1578), .B1(n1705), .B2(n1581), .ZN(n1828)
         );
  XNOR2_X1 U1455 ( .A(n1606), .B(n1829), .ZN(n836) );
  AOI221_X1 U1456 ( .B1(n1579), .B2(b[16]), .C1(n1580), .C2(b[15]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1457 ( .A1(n1708), .A2(n1578), .B1(n1709), .B2(n1581), .ZN(n1830)
         );
  XNOR2_X1 U1458 ( .A(n1606), .B(n1831), .ZN(n835) );
  AOI221_X1 U1459 ( .B1(n1579), .B2(b[17]), .C1(n1580), .C2(b[16]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1460 ( .A1(n1712), .A2(n1578), .B1(n1713), .B2(n1581), .ZN(n1832)
         );
  XNOR2_X1 U1461 ( .A(n1606), .B(n1833), .ZN(n834) );
  AOI221_X1 U1462 ( .B1(n1579), .B2(b[18]), .C1(n1580), .C2(b[17]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1463 ( .A1(n1716), .A2(n1578), .B1(n1717), .B2(n1581), .ZN(n1834)
         );
  XNOR2_X1 U1464 ( .A(n1606), .B(n1835), .ZN(n833) );
  AOI221_X1 U1465 ( .B1(n1579), .B2(b[19]), .C1(n1580), .C2(b[18]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1466 ( .A1(n1720), .A2(n1578), .B1(n1721), .B2(n1581), .ZN(n1836)
         );
  XNOR2_X1 U1467 ( .A(n1606), .B(n1837), .ZN(n832) );
  AOI221_X1 U1468 ( .B1(n1579), .B2(b[20]), .C1(n1580), .C2(b[19]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1469 ( .A1(n1724), .A2(n1578), .B1(n1725), .B2(n1581), .ZN(n1838)
         );
  XNOR2_X1 U1470 ( .A(a[11]), .B(n1839), .ZN(n831) );
  AOI221_X1 U1471 ( .B1(n1579), .B2(b[21]), .C1(n1580), .C2(b[20]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1472 ( .A1(n1728), .A2(n1578), .B1(n1729), .B2(n1581), .ZN(n1840)
         );
  XNOR2_X1 U1473 ( .A(a[11]), .B(n1841), .ZN(n830) );
  AOI221_X1 U1474 ( .B1(n1579), .B2(b[22]), .C1(n1553), .C2(n1376), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1475 ( .A1(n1640), .A2(n1582), .B1(n1643), .B2(n1537), .ZN(n1842)
         );
  XNOR2_X1 U1476 ( .A(a[11]), .B(n1843), .ZN(n829) );
  AOI221_X1 U1477 ( .B1(n1580), .B2(b[22]), .C1(n1553), .C2(n1375), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1478 ( .A1(n1617), .A2(n1542), .B1(n1643), .B2(n1581), .ZN(n1844)
         );
  XNOR2_X1 U1479 ( .A(a[11]), .B(n1845), .ZN(n828) );
  AOI221_X1 U1480 ( .B1(n1579), .B2(n1614), .C1(n1580), .C2(n1614), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1481 ( .A1(n1633), .A2(n1578), .B1(n1634), .B2(n1581), .ZN(n1846)
         );
  XNOR2_X1 U1482 ( .A(a[11]), .B(n1847), .ZN(n827) );
  OAI221_X1 U1483 ( .B1(n1616), .B2(n1582), .C1(n1617), .C2(n1578), .A(n1848), 
        .ZN(n1847) );
  OAI21_X1 U1484 ( .B1(n1579), .B2(n1580), .A(n1614), .ZN(n1848) );
  INV_X1 U1485 ( .A(n1852), .ZN(n1849) );
  NAND3_X1 U1486 ( .A1(n1852), .A2(n1851), .A3(n1850), .ZN(n1802) );
  XNOR2_X1 U1487 ( .A(a[10]), .B(a[9]), .ZN(n1850) );
  XNOR2_X1 U1488 ( .A(a[10]), .B(n1607), .ZN(n1851) );
  XOR2_X1 U1489 ( .A(a[9]), .B(n1609), .Z(n1852) );
  XNOR2_X1 U1490 ( .A(n1853), .B(n1605), .ZN(n826) );
  OAI22_X1 U1491 ( .A1(n1565), .A2(n1541), .B1(n1565), .B2(n1583), .ZN(n1853)
         );
  XNOR2_X1 U1492 ( .A(n1854), .B(n1605), .ZN(n825) );
  OAI222_X1 U1493 ( .A1(n1649), .A2(n1541), .B1(n1566), .B2(n1549), .C1(n1650), 
        .C2(n1583), .ZN(n1854) );
  XNOR2_X1 U1494 ( .A(n1604), .B(n1855), .ZN(n824) );
  AOI221_X1 U1495 ( .B1(n1584), .B2(b[2]), .C1(n1585), .C2(b[1]), .A(n1856), 
        .ZN(n1855) );
  OAI22_X1 U1496 ( .A1(n1653), .A2(n1583), .B1(n1565), .B2(n1586), .ZN(n1856)
         );
  XNOR2_X1 U1497 ( .A(n1604), .B(n1858), .ZN(n823) );
  AOI221_X1 U1498 ( .B1(n1584), .B2(b[3]), .C1(n1585), .C2(b[2]), .A(n1859), 
        .ZN(n1858) );
  OAI22_X1 U1499 ( .A1(n1657), .A2(n1583), .B1(n1649), .B2(n1587), .ZN(n1859)
         );
  XNOR2_X1 U1500 ( .A(n1604), .B(n1860), .ZN(n822) );
  AOI221_X1 U1501 ( .B1(n1584), .B2(b[4]), .C1(n1585), .C2(b[3]), .A(n1861), 
        .ZN(n1860) );
  OAI22_X1 U1502 ( .A1(n1660), .A2(n1583), .B1(n1661), .B2(n1587), .ZN(n1861)
         );
  XNOR2_X1 U1503 ( .A(n1604), .B(n1862), .ZN(n821) );
  AOI221_X1 U1504 ( .B1(n1584), .B2(b[5]), .C1(n1585), .C2(b[4]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1505 ( .A1(n1664), .A2(n1583), .B1(n1665), .B2(n1587), .ZN(n1863)
         );
  XNOR2_X1 U1506 ( .A(n1604), .B(n1864), .ZN(n820) );
  AOI221_X1 U1507 ( .B1(n1584), .B2(b[6]), .C1(n1585), .C2(b[5]), .A(n1865), 
        .ZN(n1864) );
  OAI22_X1 U1508 ( .A1(n1668), .A2(n1583), .B1(n1669), .B2(n1587), .ZN(n1865)
         );
  XNOR2_X1 U1509 ( .A(n1604), .B(n1866), .ZN(n819) );
  AOI221_X1 U1510 ( .B1(n1584), .B2(b[7]), .C1(n1585), .C2(b[6]), .A(n1867), 
        .ZN(n1866) );
  OAI22_X1 U1511 ( .A1(n1672), .A2(n1583), .B1(n1673), .B2(n1587), .ZN(n1867)
         );
  XNOR2_X1 U1512 ( .A(n1604), .B(n1868), .ZN(n818) );
  AOI221_X1 U1513 ( .B1(n1584), .B2(b[8]), .C1(n1585), .C2(b[7]), .A(n1869), 
        .ZN(n1868) );
  OAI22_X1 U1514 ( .A1(n1676), .A2(n1583), .B1(n1677), .B2(n1587), .ZN(n1869)
         );
  XNOR2_X1 U1515 ( .A(n1604), .B(n1870), .ZN(n817) );
  AOI221_X1 U1516 ( .B1(n1584), .B2(b[9]), .C1(n1585), .C2(b[8]), .A(n1871), 
        .ZN(n1870) );
  OAI22_X1 U1517 ( .A1(n1680), .A2(n1583), .B1(n1681), .B2(n1587), .ZN(n1871)
         );
  XNOR2_X1 U1518 ( .A(n1604), .B(n1872), .ZN(n816) );
  AOI221_X1 U1519 ( .B1(n1584), .B2(b[10]), .C1(n1585), .C2(b[9]), .A(n1873), 
        .ZN(n1872) );
  OAI22_X1 U1520 ( .A1(n1684), .A2(n1583), .B1(n1685), .B2(n1587), .ZN(n1873)
         );
  XNOR2_X1 U1521 ( .A(n1604), .B(n1874), .ZN(n815) );
  AOI221_X1 U1522 ( .B1(n1584), .B2(b[11]), .C1(n1585), .C2(b[10]), .A(n1875), 
        .ZN(n1874) );
  OAI22_X1 U1523 ( .A1(n1688), .A2(n1583), .B1(n1689), .B2(n1587), .ZN(n1875)
         );
  XNOR2_X1 U1524 ( .A(n1604), .B(n1876), .ZN(n814) );
  AOI221_X1 U1525 ( .B1(n1584), .B2(b[12]), .C1(n1585), .C2(b[11]), .A(n1877), 
        .ZN(n1876) );
  OAI22_X1 U1526 ( .A1(n1692), .A2(n1583), .B1(n1693), .B2(n1587), .ZN(n1877)
         );
  XNOR2_X1 U1527 ( .A(n1604), .B(n1878), .ZN(n813) );
  AOI221_X1 U1528 ( .B1(n1584), .B2(b[13]), .C1(n1585), .C2(b[12]), .A(n1879), 
        .ZN(n1878) );
  OAI22_X1 U1529 ( .A1(n1696), .A2(n1583), .B1(n1697), .B2(n1586), .ZN(n1879)
         );
  XNOR2_X1 U1530 ( .A(n1604), .B(n1880), .ZN(n812) );
  AOI221_X1 U1531 ( .B1(n1584), .B2(b[14]), .C1(n1585), .C2(b[13]), .A(n1881), 
        .ZN(n1880) );
  OAI22_X1 U1532 ( .A1(n1700), .A2(n1583), .B1(n1701), .B2(n1586), .ZN(n1881)
         );
  XNOR2_X1 U1533 ( .A(n1604), .B(n1882), .ZN(n811) );
  AOI221_X1 U1534 ( .B1(n1584), .B2(b[15]), .C1(n1585), .C2(b[14]), .A(n1883), 
        .ZN(n1882) );
  OAI22_X1 U1535 ( .A1(n1704), .A2(n1583), .B1(n1705), .B2(n1586), .ZN(n1883)
         );
  XNOR2_X1 U1536 ( .A(n1604), .B(n1884), .ZN(n810) );
  AOI221_X1 U1537 ( .B1(n1584), .B2(b[16]), .C1(n1585), .C2(b[15]), .A(n1885), 
        .ZN(n1884) );
  OAI22_X1 U1538 ( .A1(n1708), .A2(n1583), .B1(n1709), .B2(n1586), .ZN(n1885)
         );
  XNOR2_X1 U1539 ( .A(n1604), .B(n1886), .ZN(n809) );
  AOI221_X1 U1540 ( .B1(n1584), .B2(b[17]), .C1(n1585), .C2(b[16]), .A(n1887), 
        .ZN(n1886) );
  OAI22_X1 U1541 ( .A1(n1712), .A2(n1583), .B1(n1713), .B2(n1586), .ZN(n1887)
         );
  XNOR2_X1 U1542 ( .A(n1604), .B(n1888), .ZN(n808) );
  AOI221_X1 U1543 ( .B1(n1584), .B2(b[18]), .C1(n1585), .C2(b[17]), .A(n1889), 
        .ZN(n1888) );
  OAI22_X1 U1544 ( .A1(n1716), .A2(n1583), .B1(n1717), .B2(n1586), .ZN(n1889)
         );
  XNOR2_X1 U1545 ( .A(n1604), .B(n1890), .ZN(n807) );
  AOI221_X1 U1546 ( .B1(n1584), .B2(b[19]), .C1(n1585), .C2(b[18]), .A(n1891), 
        .ZN(n1890) );
  OAI22_X1 U1547 ( .A1(n1720), .A2(n1583), .B1(n1721), .B2(n1586), .ZN(n1891)
         );
  XNOR2_X1 U1548 ( .A(n1604), .B(n1892), .ZN(n806) );
  AOI221_X1 U1549 ( .B1(n1584), .B2(b[20]), .C1(n1585), .C2(b[19]), .A(n1893), 
        .ZN(n1892) );
  OAI22_X1 U1550 ( .A1(n1724), .A2(n1583), .B1(n1725), .B2(n1586), .ZN(n1893)
         );
  XNOR2_X1 U1551 ( .A(a[14]), .B(n1894), .ZN(n805) );
  AOI221_X1 U1552 ( .B1(n1584), .B2(b[21]), .C1(n1585), .C2(b[20]), .A(n1895), 
        .ZN(n1894) );
  OAI22_X1 U1553 ( .A1(n1728), .A2(n1583), .B1(n1729), .B2(n1586), .ZN(n1895)
         );
  XNOR2_X1 U1554 ( .A(a[14]), .B(n1896), .ZN(n804) );
  AOI221_X1 U1555 ( .B1(n1584), .B2(b[22]), .C1(n1552), .C2(n1376), .A(n1897), 
        .ZN(n1896) );
  OAI22_X1 U1556 ( .A1(n1640), .A2(n1587), .B1(n1643), .B2(n1549), .ZN(n1897)
         );
  XNOR2_X1 U1557 ( .A(a[14]), .B(n1898), .ZN(n803) );
  AOI221_X1 U1558 ( .B1(n1585), .B2(b[22]), .C1(n1552), .C2(n1375), .A(n1899), 
        .ZN(n1898) );
  OAI22_X1 U1559 ( .A1(n1617), .A2(n1541), .B1(n1643), .B2(n1586), .ZN(n1899)
         );
  XNOR2_X1 U1560 ( .A(a[14]), .B(n1900), .ZN(n802) );
  AOI221_X1 U1561 ( .B1(n1584), .B2(n1614), .C1(n1585), .C2(n1614), .A(n1901), 
        .ZN(n1900) );
  OAI22_X1 U1562 ( .A1(n1633), .A2(n1583), .B1(n1634), .B2(n1586), .ZN(n1901)
         );
  XNOR2_X1 U1563 ( .A(a[14]), .B(n1902), .ZN(n801) );
  OAI221_X1 U1564 ( .B1(n1617), .B2(n1587), .C1(n1619), .C2(n1583), .A(n1903), 
        .ZN(n1902) );
  OAI21_X1 U1565 ( .B1(n1584), .B2(n1585), .A(n1614), .ZN(n1903) );
  INV_X1 U1566 ( .A(n1907), .ZN(n1904) );
  NAND3_X1 U1567 ( .A1(n1907), .A2(n1906), .A3(n1905), .ZN(n1857) );
  XNOR2_X1 U1568 ( .A(a[12]), .B(a[13]), .ZN(n1905) );
  XNOR2_X1 U1569 ( .A(a[13]), .B(n1605), .ZN(n1906) );
  XOR2_X1 U1570 ( .A(a[12]), .B(n1607), .Z(n1907) );
  XNOR2_X1 U1571 ( .A(n1908), .B(n1603), .ZN(n800) );
  OAI22_X1 U1572 ( .A1(n1565), .A2(n1540), .B1(n1566), .B2(n1588), .ZN(n1908)
         );
  XNOR2_X1 U1573 ( .A(n1909), .B(n1603), .ZN(n799) );
  OAI222_X1 U1574 ( .A1(n1649), .A2(n1540), .B1(n1566), .B2(n1548), .C1(n1650), 
        .C2(n1588), .ZN(n1909) );
  XNOR2_X1 U1575 ( .A(n1602), .B(n1910), .ZN(n798) );
  AOI221_X1 U1576 ( .B1(n1589), .B2(b[2]), .C1(n1590), .C2(b[1]), .A(n1911), 
        .ZN(n1910) );
  OAI22_X1 U1577 ( .A1(n1653), .A2(n1588), .B1(n1566), .B2(n1591), .ZN(n1911)
         );
  XNOR2_X1 U1578 ( .A(n1602), .B(n1913), .ZN(n797) );
  AOI221_X1 U1579 ( .B1(n1589), .B2(b[3]), .C1(n1590), .C2(b[2]), .A(n1914), 
        .ZN(n1913) );
  OAI22_X1 U1580 ( .A1(n1657), .A2(n1588), .B1(n1649), .B2(n1592), .ZN(n1914)
         );
  XNOR2_X1 U1581 ( .A(n1602), .B(n1915), .ZN(n796) );
  AOI221_X1 U1582 ( .B1(n1589), .B2(b[4]), .C1(n1590), .C2(b[3]), .A(n1916), 
        .ZN(n1915) );
  OAI22_X1 U1583 ( .A1(n1660), .A2(n1588), .B1(n1661), .B2(n1592), .ZN(n1916)
         );
  XNOR2_X1 U1584 ( .A(n1602), .B(n1917), .ZN(n795) );
  AOI221_X1 U1585 ( .B1(n1589), .B2(b[5]), .C1(n1590), .C2(b[4]), .A(n1918), 
        .ZN(n1917) );
  OAI22_X1 U1586 ( .A1(n1664), .A2(n1588), .B1(n1665), .B2(n1592), .ZN(n1918)
         );
  XNOR2_X1 U1587 ( .A(n1602), .B(n1919), .ZN(n794) );
  AOI221_X1 U1588 ( .B1(n1589), .B2(b[6]), .C1(n1590), .C2(b[5]), .A(n1920), 
        .ZN(n1919) );
  OAI22_X1 U1589 ( .A1(n1668), .A2(n1588), .B1(n1669), .B2(n1592), .ZN(n1920)
         );
  XNOR2_X1 U1590 ( .A(n1602), .B(n1921), .ZN(n793) );
  AOI221_X1 U1591 ( .B1(n1589), .B2(b[7]), .C1(n1590), .C2(b[6]), .A(n1922), 
        .ZN(n1921) );
  OAI22_X1 U1592 ( .A1(n1672), .A2(n1588), .B1(n1673), .B2(n1592), .ZN(n1922)
         );
  XNOR2_X1 U1593 ( .A(n1602), .B(n1923), .ZN(n792) );
  AOI221_X1 U1594 ( .B1(n1589), .B2(b[8]), .C1(n1590), .C2(b[7]), .A(n1924), 
        .ZN(n1923) );
  OAI22_X1 U1595 ( .A1(n1676), .A2(n1588), .B1(n1677), .B2(n1592), .ZN(n1924)
         );
  XNOR2_X1 U1596 ( .A(n1602), .B(n1925), .ZN(n791) );
  AOI221_X1 U1597 ( .B1(n1589), .B2(b[9]), .C1(n1590), .C2(b[8]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1598 ( .A1(n1680), .A2(n1588), .B1(n1681), .B2(n1592), .ZN(n1926)
         );
  XNOR2_X1 U1599 ( .A(n1602), .B(n1927), .ZN(n790) );
  AOI221_X1 U1600 ( .B1(n1589), .B2(b[10]), .C1(n1590), .C2(b[9]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1601 ( .A1(n1684), .A2(n1588), .B1(n1685), .B2(n1592), .ZN(n1928)
         );
  XNOR2_X1 U1602 ( .A(n1602), .B(n1929), .ZN(n789) );
  AOI221_X1 U1603 ( .B1(n1589), .B2(b[11]), .C1(n1590), .C2(b[10]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1604 ( .A1(n1688), .A2(n1588), .B1(n1689), .B2(n1592), .ZN(n1930)
         );
  XNOR2_X1 U1605 ( .A(n1602), .B(n1931), .ZN(n788) );
  AOI221_X1 U1606 ( .B1(n1589), .B2(b[12]), .C1(n1590), .C2(b[11]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1607 ( .A1(n1692), .A2(n1588), .B1(n1693), .B2(n1592), .ZN(n1932)
         );
  XNOR2_X1 U1608 ( .A(n1602), .B(n1933), .ZN(n787) );
  AOI221_X1 U1609 ( .B1(n1589), .B2(b[13]), .C1(n1590), .C2(b[12]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1610 ( .A1(n1696), .A2(n1588), .B1(n1697), .B2(n1591), .ZN(n1934)
         );
  XNOR2_X1 U1611 ( .A(n1602), .B(n1935), .ZN(n786) );
  AOI221_X1 U1612 ( .B1(n1589), .B2(b[14]), .C1(n1590), .C2(b[13]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1613 ( .A1(n1700), .A2(n1588), .B1(n1701), .B2(n1591), .ZN(n1936)
         );
  XNOR2_X1 U1614 ( .A(n1602), .B(n1937), .ZN(n785) );
  AOI221_X1 U1615 ( .B1(n1589), .B2(b[15]), .C1(n1590), .C2(b[14]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1616 ( .A1(n1704), .A2(n1588), .B1(n1705), .B2(n1591), .ZN(n1938)
         );
  XNOR2_X1 U1617 ( .A(n1602), .B(n1939), .ZN(n784) );
  AOI221_X1 U1618 ( .B1(n1589), .B2(b[16]), .C1(n1590), .C2(b[15]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1619 ( .A1(n1708), .A2(n1588), .B1(n1709), .B2(n1591), .ZN(n1940)
         );
  XNOR2_X1 U1620 ( .A(n1602), .B(n1941), .ZN(n783) );
  AOI221_X1 U1621 ( .B1(n1589), .B2(b[17]), .C1(n1590), .C2(b[16]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1622 ( .A1(n1712), .A2(n1588), .B1(n1713), .B2(n1591), .ZN(n1942)
         );
  XNOR2_X1 U1623 ( .A(n1602), .B(n1943), .ZN(n782) );
  AOI221_X1 U1624 ( .B1(n1589), .B2(b[18]), .C1(n1590), .C2(b[17]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1625 ( .A1(n1716), .A2(n1588), .B1(n1717), .B2(n1591), .ZN(n1944)
         );
  XNOR2_X1 U1626 ( .A(n1602), .B(n1945), .ZN(n781) );
  AOI221_X1 U1627 ( .B1(n1589), .B2(b[19]), .C1(n1590), .C2(b[18]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1628 ( .A1(n1720), .A2(n1588), .B1(n1721), .B2(n1591), .ZN(n1946)
         );
  XNOR2_X1 U1629 ( .A(n1602), .B(n1947), .ZN(n780) );
  AOI221_X1 U1630 ( .B1(n1589), .B2(b[20]), .C1(n1590), .C2(b[19]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1631 ( .A1(n1724), .A2(n1588), .B1(n1725), .B2(n1591), .ZN(n1948)
         );
  XNOR2_X1 U1632 ( .A(a[17]), .B(n1949), .ZN(n779) );
  AOI221_X1 U1633 ( .B1(n1589), .B2(b[21]), .C1(n1590), .C2(b[20]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1634 ( .A1(n1728), .A2(n1588), .B1(n1729), .B2(n1591), .ZN(n1950)
         );
  XNOR2_X1 U1635 ( .A(a[17]), .B(n1951), .ZN(n778) );
  AOI221_X1 U1636 ( .B1(n1589), .B2(b[22]), .C1(n1551), .C2(n1376), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1637 ( .A1(n1640), .A2(n1592), .B1(n1643), .B2(n1548), .ZN(n1952)
         );
  XNOR2_X1 U1638 ( .A(a[17]), .B(n1953), .ZN(n777) );
  AOI221_X1 U1639 ( .B1(n1590), .B2(b[22]), .C1(n1551), .C2(n1375), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1640 ( .A1(n1617), .A2(n1540), .B1(n1643), .B2(n1591), .ZN(n1954)
         );
  XNOR2_X1 U1641 ( .A(a[17]), .B(n1955), .ZN(n776) );
  AOI221_X1 U1642 ( .B1(n1589), .B2(n1613), .C1(n1590), .C2(n1614), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1643 ( .A1(n1633), .A2(n1588), .B1(n1634), .B2(n1591), .ZN(n1956)
         );
  XNOR2_X1 U1644 ( .A(a[17]), .B(n1957), .ZN(n775) );
  OAI221_X1 U1645 ( .B1(n1618), .B2(n1592), .C1(n1617), .C2(n1588), .A(n1958), 
        .ZN(n1957) );
  OAI21_X1 U1646 ( .B1(n1589), .B2(n1590), .A(n1614), .ZN(n1958) );
  INV_X1 U1647 ( .A(n1962), .ZN(n1959) );
  NAND3_X1 U1648 ( .A1(n1962), .A2(n1961), .A3(n1960), .ZN(n1912) );
  XNOR2_X1 U1649 ( .A(a[15]), .B(a[16]), .ZN(n1960) );
  XNOR2_X1 U1650 ( .A(a[16]), .B(n1603), .ZN(n1961) );
  XOR2_X1 U1651 ( .A(a[15]), .B(n1605), .Z(n1962) );
  XOR2_X1 U1652 ( .A(n1963), .B(n1600), .Z(n774) );
  OAI22_X1 U1653 ( .A1(n1565), .A2(n1539), .B1(n1566), .B2(n1593), .ZN(n1963)
         );
  XOR2_X1 U1654 ( .A(n1964), .B(n1600), .Z(n773) );
  OAI222_X1 U1655 ( .A1(n1649), .A2(n1539), .B1(n1566), .B2(n1547), .C1(n1650), 
        .C2(n1593), .ZN(n1964) );
  XNOR2_X1 U1656 ( .A(n1600), .B(n1965), .ZN(n772) );
  AOI221_X1 U1657 ( .B1(n1594), .B2(b[2]), .C1(n1595), .C2(b[1]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1658 ( .A1(n1653), .A2(n1593), .B1(n1566), .B2(n1596), .ZN(n1966)
         );
  XNOR2_X1 U1659 ( .A(n1600), .B(n1968), .ZN(n771) );
  AOI221_X1 U1660 ( .B1(n1594), .B2(b[3]), .C1(n1595), .C2(b[2]), .A(n1969), 
        .ZN(n1968) );
  OAI22_X1 U1661 ( .A1(n1657), .A2(n1593), .B1(n1649), .B2(n1597), .ZN(n1969)
         );
  XNOR2_X1 U1662 ( .A(n1600), .B(n1970), .ZN(n770) );
  AOI221_X1 U1663 ( .B1(n1594), .B2(b[4]), .C1(n1595), .C2(b[3]), .A(n1971), 
        .ZN(n1970) );
  OAI22_X1 U1664 ( .A1(n1660), .A2(n1593), .B1(n1661), .B2(n1597), .ZN(n1971)
         );
  XNOR2_X1 U1665 ( .A(n1600), .B(n1972), .ZN(n769) );
  AOI221_X1 U1666 ( .B1(n1594), .B2(b[5]), .C1(n1595), .C2(b[4]), .A(n1973), 
        .ZN(n1972) );
  OAI22_X1 U1667 ( .A1(n1664), .A2(n1593), .B1(n1665), .B2(n1597), .ZN(n1973)
         );
  XNOR2_X1 U1668 ( .A(n1600), .B(n1974), .ZN(n768) );
  AOI221_X1 U1669 ( .B1(n1594), .B2(b[6]), .C1(n1595), .C2(b[5]), .A(n1975), 
        .ZN(n1974) );
  OAI22_X1 U1670 ( .A1(n1668), .A2(n1593), .B1(n1669), .B2(n1597), .ZN(n1975)
         );
  XNOR2_X1 U1671 ( .A(n1600), .B(n1976), .ZN(n767) );
  AOI221_X1 U1672 ( .B1(n1594), .B2(b[7]), .C1(n1595), .C2(b[6]), .A(n1977), 
        .ZN(n1976) );
  OAI22_X1 U1673 ( .A1(n1672), .A2(n1593), .B1(n1673), .B2(n1597), .ZN(n1977)
         );
  XNOR2_X1 U1674 ( .A(n1600), .B(n1978), .ZN(n766) );
  AOI221_X1 U1675 ( .B1(n1594), .B2(b[8]), .C1(n1595), .C2(b[7]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1676 ( .A1(n1676), .A2(n1593), .B1(n1677), .B2(n1597), .ZN(n1979)
         );
  XNOR2_X1 U1677 ( .A(n1600), .B(n1980), .ZN(n765) );
  AOI221_X1 U1678 ( .B1(n1594), .B2(b[9]), .C1(n1595), .C2(b[8]), .A(n1981), 
        .ZN(n1980) );
  OAI22_X1 U1679 ( .A1(n1680), .A2(n1593), .B1(n1681), .B2(n1597), .ZN(n1981)
         );
  XNOR2_X1 U1680 ( .A(n1600), .B(n1982), .ZN(n764) );
  AOI221_X1 U1681 ( .B1(n1594), .B2(b[10]), .C1(n1595), .C2(b[9]), .A(n1983), 
        .ZN(n1982) );
  OAI22_X1 U1682 ( .A1(n1684), .A2(n1593), .B1(n1685), .B2(n1597), .ZN(n1983)
         );
  XNOR2_X1 U1683 ( .A(n1600), .B(n1984), .ZN(n763) );
  AOI221_X1 U1684 ( .B1(n1594), .B2(b[11]), .C1(n1595), .C2(b[10]), .A(n1985), 
        .ZN(n1984) );
  OAI22_X1 U1685 ( .A1(n1688), .A2(n1593), .B1(n1689), .B2(n1597), .ZN(n1985)
         );
  XNOR2_X1 U1686 ( .A(n1601), .B(n1986), .ZN(n762) );
  AOI221_X1 U1687 ( .B1(n1594), .B2(b[12]), .C1(n1595), .C2(b[11]), .A(n1987), 
        .ZN(n1986) );
  OAI22_X1 U1688 ( .A1(n1692), .A2(n1593), .B1(n1693), .B2(n1597), .ZN(n1987)
         );
  XNOR2_X1 U1689 ( .A(n1601), .B(n1988), .ZN(n761) );
  AOI221_X1 U1690 ( .B1(n1594), .B2(b[13]), .C1(n1595), .C2(b[12]), .A(n1989), 
        .ZN(n1988) );
  OAI22_X1 U1691 ( .A1(n1696), .A2(n1593), .B1(n1697), .B2(n1596), .ZN(n1989)
         );
  XNOR2_X1 U1692 ( .A(n1601), .B(n1990), .ZN(n760) );
  AOI221_X1 U1693 ( .B1(n1594), .B2(b[14]), .C1(n1595), .C2(b[13]), .A(n1991), 
        .ZN(n1990) );
  OAI22_X1 U1694 ( .A1(n1700), .A2(n1593), .B1(n1701), .B2(n1596), .ZN(n1991)
         );
  XNOR2_X1 U1695 ( .A(n1601), .B(n1992), .ZN(n759) );
  AOI221_X1 U1696 ( .B1(n1594), .B2(b[15]), .C1(n1595), .C2(b[14]), .A(n1993), 
        .ZN(n1992) );
  OAI22_X1 U1697 ( .A1(n1704), .A2(n1593), .B1(n1705), .B2(n1596), .ZN(n1993)
         );
  XNOR2_X1 U1698 ( .A(n1601), .B(n1994), .ZN(n758) );
  AOI221_X1 U1699 ( .B1(n1594), .B2(b[16]), .C1(n1595), .C2(b[15]), .A(n1995), 
        .ZN(n1994) );
  OAI22_X1 U1700 ( .A1(n1708), .A2(n1593), .B1(n1709), .B2(n1596), .ZN(n1995)
         );
  XNOR2_X1 U1701 ( .A(n1601), .B(n1996), .ZN(n757) );
  AOI221_X1 U1702 ( .B1(n1594), .B2(b[17]), .C1(n1595), .C2(b[16]), .A(n1997), 
        .ZN(n1996) );
  OAI22_X1 U1703 ( .A1(n1712), .A2(n1593), .B1(n1713), .B2(n1596), .ZN(n1997)
         );
  XNOR2_X1 U1704 ( .A(n1601), .B(n1998), .ZN(n756) );
  AOI221_X1 U1705 ( .B1(n1594), .B2(b[18]), .C1(n1595), .C2(b[17]), .A(n1999), 
        .ZN(n1998) );
  OAI22_X1 U1706 ( .A1(n1716), .A2(n1593), .B1(n1717), .B2(n1596), .ZN(n1999)
         );
  XNOR2_X1 U1707 ( .A(n1601), .B(n2000), .ZN(n755) );
  AOI221_X1 U1708 ( .B1(n1594), .B2(b[19]), .C1(n1595), .C2(b[18]), .A(n2001), 
        .ZN(n2000) );
  OAI22_X1 U1709 ( .A1(n1720), .A2(n1593), .B1(n1721), .B2(n1596), .ZN(n2001)
         );
  XNOR2_X1 U1710 ( .A(n1601), .B(n2002), .ZN(n754) );
  AOI221_X1 U1711 ( .B1(n1594), .B2(b[20]), .C1(n1595), .C2(b[19]), .A(n2003), 
        .ZN(n2002) );
  OAI22_X1 U1712 ( .A1(n1724), .A2(n1593), .B1(n1725), .B2(n1596), .ZN(n2003)
         );
  XNOR2_X1 U1713 ( .A(n1601), .B(n2004), .ZN(n753) );
  AOI221_X1 U1714 ( .B1(n1594), .B2(b[21]), .C1(n1595), .C2(b[20]), .A(n2005), 
        .ZN(n2004) );
  OAI22_X1 U1715 ( .A1(n1728), .A2(n1593), .B1(n1729), .B2(n1596), .ZN(n2005)
         );
  XNOR2_X1 U1716 ( .A(n1601), .B(n2006), .ZN(n752) );
  AOI221_X1 U1717 ( .B1(n1594), .B2(b[22]), .C1(n1545), .C2(n1376), .A(n2007), 
        .ZN(n2006) );
  OAI22_X1 U1718 ( .A1(n1640), .A2(n1597), .B1(n1643), .B2(n1547), .ZN(n2007)
         );
  XNOR2_X1 U1719 ( .A(n1601), .B(n2008), .ZN(n751) );
  AOI221_X1 U1720 ( .B1(n1595), .B2(b[22]), .C1(n1545), .C2(n1375), .A(n2009), 
        .ZN(n2008) );
  OAI22_X1 U1721 ( .A1(n1617), .A2(n1539), .B1(n1643), .B2(n1596), .ZN(n2009)
         );
  XNOR2_X1 U1722 ( .A(n1601), .B(n2010), .ZN(n750) );
  AOI221_X1 U1723 ( .B1(n1594), .B2(n1612), .C1(n1595), .C2(n1614), .A(n2011), 
        .ZN(n2010) );
  OAI22_X1 U1724 ( .A1(n1633), .A2(n1593), .B1(n1634), .B2(n1596), .ZN(n2011)
         );
  INV_X1 U1725 ( .A(b[22]), .ZN(n1634) );
  INV_X1 U1726 ( .A(n1374), .ZN(n1633) );
  XNOR2_X1 U1727 ( .A(n1600), .B(n2012), .ZN(n749) );
  OAI221_X1 U1728 ( .B1(n1617), .B2(n1597), .C1(n1619), .C2(n1593), .A(n2013), 
        .ZN(n2012) );
  OAI21_X1 U1729 ( .B1(n1594), .B2(n1595), .A(n1614), .ZN(n2013) );
  INV_X1 U1730 ( .A(n2017), .ZN(n2014) );
  NAND3_X1 U1731 ( .A1(n2017), .A2(n2016), .A3(n2015), .ZN(n1967) );
  XNOR2_X1 U1732 ( .A(a[18]), .B(a[19]), .ZN(n2015) );
  XOR2_X1 U1733 ( .A(a[19]), .B(n1600), .Z(n2016) );
  XOR2_X1 U1734 ( .A(a[18]), .B(n1603), .Z(n2017) );
  XNOR2_X1 U1735 ( .A(n2018), .B(n1599), .ZN(n748) );
  OAI22_X1 U1736 ( .A1(n1538), .A2(n1567), .B1(n1558), .B2(n1567), .ZN(n2018)
         );
  XNOR2_X1 U1737 ( .A(n2019), .B(n1599), .ZN(n747) );
  OAI222_X1 U1738 ( .A1(n1538), .A2(n1649), .B1(n1546), .B2(n1566), .C1(n1558), 
        .C2(n1650), .ZN(n2019) );
  XNOR2_X1 U1739 ( .A(n1598), .B(n2020), .ZN(n746) );
  AOI221_X1 U1740 ( .B1(b[2]), .B2(n1559), .C1(b[1]), .C2(n1560), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1741 ( .A1(n1558), .A2(n1653), .B1(n1557), .B2(n1567), .ZN(n2021)
         );
  INV_X1 U1742 ( .A(b[0]), .ZN(n1647) );
  INV_X1 U1743 ( .A(n1396), .ZN(n1653) );
  XNOR2_X1 U1744 ( .A(n1598), .B(n2022), .ZN(n745) );
  AOI221_X1 U1745 ( .B1(b[3]), .B2(n1559), .C1(b[2]), .C2(n1560), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1746 ( .A1(n1558), .A2(n1657), .B1(n1557), .B2(n1649), .ZN(n2023)
         );
  XNOR2_X1 U1747 ( .A(n1598), .B(n2024), .ZN(n744) );
  AOI221_X1 U1748 ( .B1(b[4]), .B2(n1559), .C1(b[3]), .C2(n1560), .A(n2025), 
        .ZN(n2024) );
  OAI22_X1 U1749 ( .A1(n1558), .A2(n1660), .B1(n1557), .B2(n1661), .ZN(n2025)
         );
  XNOR2_X1 U1750 ( .A(n1598), .B(n2026), .ZN(n743) );
  AOI221_X1 U1751 ( .B1(b[5]), .B2(n1559), .C1(b[4]), .C2(n1560), .A(n2027), 
        .ZN(n2026) );
  OAI22_X1 U1752 ( .A1(n1558), .A2(n1664), .B1(n1557), .B2(n1665), .ZN(n2027)
         );
  XNOR2_X1 U1753 ( .A(n1598), .B(n2028), .ZN(n742) );
  AOI221_X1 U1754 ( .B1(b[6]), .B2(n1559), .C1(b[5]), .C2(n1560), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1755 ( .A1(n1558), .A2(n1668), .B1(n1557), .B2(n1669), .ZN(n2029)
         );
  XNOR2_X1 U1756 ( .A(n1598), .B(n2030), .ZN(n741) );
  AOI221_X1 U1757 ( .B1(b[7]), .B2(n1559), .C1(b[6]), .C2(n1560), .A(n2031), 
        .ZN(n2030) );
  OAI22_X1 U1758 ( .A1(n1558), .A2(n1672), .B1(n1557), .B2(n1673), .ZN(n2031)
         );
  XNOR2_X1 U1759 ( .A(n1598), .B(n2032), .ZN(n740) );
  AOI221_X1 U1760 ( .B1(b[9]), .B2(n1559), .C1(b[8]), .C2(n1560), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1761 ( .A1(n1558), .A2(n1680), .B1(n1557), .B2(n1681), .ZN(n2033)
         );
  XNOR2_X1 U1762 ( .A(n1598), .B(n2034), .ZN(n739) );
  AOI221_X1 U1763 ( .B1(b[10]), .B2(n1559), .C1(b[9]), .C2(n1560), .A(n2035), 
        .ZN(n2034) );
  OAI22_X1 U1764 ( .A1(n1558), .A2(n1684), .B1(n1557), .B2(n1685), .ZN(n2035)
         );
  XNOR2_X1 U1765 ( .A(n1598), .B(n2036), .ZN(n738) );
  AOI221_X1 U1766 ( .B1(b[12]), .B2(n1559), .C1(b[11]), .C2(n1560), .A(n2037), 
        .ZN(n2036) );
  OAI22_X1 U1767 ( .A1(n1558), .A2(n1692), .B1(n1557), .B2(n1693), .ZN(n2037)
         );
  XNOR2_X1 U1768 ( .A(n1598), .B(n2038), .ZN(n737) );
  AOI221_X1 U1769 ( .B1(b[13]), .B2(n1559), .C1(b[12]), .C2(n1560), .A(n2039), 
        .ZN(n2038) );
  OAI22_X1 U1770 ( .A1(n1558), .A2(n1696), .B1(n1557), .B2(n1697), .ZN(n2039)
         );
  XNOR2_X1 U1771 ( .A(n1598), .B(n2040), .ZN(n736) );
  AOI221_X1 U1772 ( .B1(b[14]), .B2(n1559), .C1(b[13]), .C2(n1560), .A(n2041), 
        .ZN(n2040) );
  OAI22_X1 U1773 ( .A1(n1558), .A2(n1700), .B1(n1556), .B2(n1701), .ZN(n2041)
         );
  XNOR2_X1 U1774 ( .A(n1598), .B(n2042), .ZN(n735) );
  AOI221_X1 U1775 ( .B1(b[15]), .B2(n1559), .C1(b[14]), .C2(n1560), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1776 ( .A1(n1558), .A2(n1704), .B1(n1556), .B2(n1705), .ZN(n2043)
         );
  XNOR2_X1 U1777 ( .A(n1598), .B(n2044), .ZN(n734) );
  AOI221_X1 U1778 ( .B1(b[16]), .B2(n1559), .C1(b[15]), .C2(n1560), .A(n2045), 
        .ZN(n2044) );
  OAI22_X1 U1779 ( .A1(n1558), .A2(n1708), .B1(n1556), .B2(n1709), .ZN(n2045)
         );
  XNOR2_X1 U1780 ( .A(n1598), .B(n2046), .ZN(n733) );
  AOI221_X1 U1781 ( .B1(b[18]), .B2(n1559), .C1(b[17]), .C2(n1560), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1782 ( .A1(n1558), .A2(n1716), .B1(n1556), .B2(n1717), .ZN(n2047)
         );
  XNOR2_X1 U1783 ( .A(n1598), .B(n2048), .ZN(n732) );
  AOI221_X1 U1784 ( .B1(b[19]), .B2(n1559), .C1(b[18]), .C2(n1560), .A(n2049), 
        .ZN(n2048) );
  OAI22_X1 U1785 ( .A1(n1558), .A2(n1720), .B1(n1556), .B2(n1721), .ZN(n2049)
         );
  XNOR2_X1 U1786 ( .A(n1598), .B(n2050), .ZN(n731) );
  AOI221_X1 U1787 ( .B1(b[20]), .B2(n1559), .C1(b[19]), .C2(n1560), .A(n2051), 
        .ZN(n2050) );
  OAI22_X1 U1788 ( .A1(n1558), .A2(n1724), .B1(n1556), .B2(n1725), .ZN(n2051)
         );
  XNOR2_X1 U1789 ( .A(a[23]), .B(n2052), .ZN(n730) );
  AOI221_X1 U1790 ( .B1(b[21]), .B2(n1559), .C1(b[20]), .C2(n1560), .A(n2053), 
        .ZN(n2052) );
  OAI22_X1 U1791 ( .A1(n1558), .A2(n1728), .B1(n1556), .B2(n1729), .ZN(n2053)
         );
  XNOR2_X1 U1792 ( .A(a[23]), .B(n2054), .ZN(n729) );
  AOI221_X1 U1793 ( .B1(b[22]), .B2(n1559), .C1(n1376), .C2(n1544), .A(n2055), 
        .ZN(n2054) );
  OAI22_X1 U1794 ( .A1(n1556), .A2(n1640), .B1(n1546), .B2(n1643), .ZN(n2055)
         );
  INV_X1 U1795 ( .A(b[20]), .ZN(n1640) );
  XNOR2_X1 U1796 ( .A(n519), .B(n2056), .ZN(n506) );
  INV_X1 U1797 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1798 ( .A1(n2056), .A2(n519), .ZN(n493) );
  XOR2_X1 U1799 ( .A(n2057), .B(n1742), .Z(n2056) );
  OAI221_X1 U1800 ( .B1(n1618), .B2(n1639), .C1(n1619), .C2(n1564), .A(n2058), 
        .ZN(n2057) );
  OAI21_X1 U1801 ( .B1(n1561), .B2(n1563), .A(n1614), .ZN(n2058) );
  INV_X1 U1802 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1803 ( .A(n1598), .B(n2059), .Z(n454) );
  AOI221_X1 U1804 ( .B1(b[8]), .B2(n1559), .C1(b[7]), .C2(n1560), .A(n2060), 
        .ZN(n2059) );
  OAI22_X1 U1805 ( .A1(n1558), .A2(n1676), .B1(n1556), .B2(n1677), .ZN(n2060)
         );
  INV_X1 U1806 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1807 ( .A(n1598), .B(n2061), .Z(n421) );
  AOI221_X1 U1808 ( .B1(b[11]), .B2(n1559), .C1(b[10]), .C2(n1560), .A(n2062), 
        .ZN(n2061) );
  OAI22_X1 U1809 ( .A1(n1558), .A2(n1688), .B1(n1556), .B2(n1689), .ZN(n2062)
         );
  INV_X1 U1810 ( .A(n387), .ZN(n395) );
  INV_X1 U1811 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1812 ( .A(n1598), .B(n2063), .Z(n374) );
  AOI221_X1 U1813 ( .B1(b[17]), .B2(n1559), .C1(b[16]), .C2(n1560), .A(n2064), 
        .ZN(n2063) );
  OAI22_X1 U1814 ( .A1(n1558), .A2(n1712), .B1(n1556), .B2(n1713), .ZN(n2064)
         );
  INV_X1 U1815 ( .A(n356), .ZN(n360) );
  INV_X1 U1816 ( .A(n1627), .ZN(n351) );
  XOR2_X1 U1817 ( .A(n1599), .B(n2065), .Z(n1627) );
  AOI221_X1 U1818 ( .B1(b[22]), .B2(n1560), .C1(n1375), .C2(n1544), .A(n2066), 
        .ZN(n2065) );
  OAI22_X1 U1819 ( .A1(n1538), .A2(n1618), .B1(n1556), .B2(n1643), .ZN(n2066)
         );
  INV_X1 U1820 ( .A(b[21]), .ZN(n1643) );
  NAND3_X1 U1821 ( .A1(n2067), .A2(n2068), .A3(n2069), .ZN(n1629) );
  XNOR2_X1 U1822 ( .A(a[22]), .B(n1599), .ZN(n2068) );
  XNOR2_X1 U1823 ( .A(a[21]), .B(a[22]), .ZN(n2069) );
  INV_X1 U1824 ( .A(n2067), .ZN(n2070) );
  XNOR2_X1 U1825 ( .A(a[21]), .B(n1600), .ZN(n2067) );
  OAI222_X1 U1826 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n2073), .C1(n2073), 
        .C2(n2072), .ZN(n326) );
  INV_X1 U1827 ( .A(n550), .ZN(n2073) );
  XNOR2_X1 U1828 ( .A(n1742), .B(n2074), .ZN(n2072) );
  AOI221_X1 U1829 ( .B1(n1561), .B2(b[21]), .C1(b[20]), .C2(n1562), .A(n2075), 
        .ZN(n2074) );
  OAI22_X1 U1830 ( .A1(n1564), .A2(n1728), .B1(n1639), .B2(n1729), .ZN(n2075)
         );
  INV_X1 U1831 ( .A(b[19]), .ZN(n1729) );
  INV_X1 U1832 ( .A(n1377), .ZN(n1728) );
  AOI222_X1 U1833 ( .A1(n2076), .A2(n2077), .B1(n2076), .B2(n564), .C1(n564), 
        .C2(n2077), .ZN(n2071) );
  XNOR2_X1 U1834 ( .A(a[2]), .B(n2078), .ZN(n2077) );
  AOI221_X1 U1835 ( .B1(b[20]), .B2(n1561), .C1(b[19]), .C2(n1562), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1836 ( .A1(n1564), .A2(n1724), .B1(n1639), .B2(n1725), .ZN(n2079)
         );
  INV_X1 U1837 ( .A(b[18]), .ZN(n1725) );
  INV_X1 U1838 ( .A(n1378), .ZN(n1724) );
  INV_X1 U1839 ( .A(n2080), .ZN(n2076) );
  AOI222_X1 U1840 ( .A1(n2081), .A2(n2082), .B1(n2081), .B2(n576), .C1(n576), 
        .C2(n2082), .ZN(n2080) );
  XNOR2_X1 U1841 ( .A(a[2]), .B(n2083), .ZN(n2082) );
  AOI221_X1 U1842 ( .B1(b[19]), .B2(n1561), .C1(b[18]), .C2(n1562), .A(n2084), 
        .ZN(n2083) );
  OAI22_X1 U1843 ( .A1(n1564), .A2(n1720), .B1(n1639), .B2(n1721), .ZN(n2084)
         );
  INV_X1 U1844 ( .A(b[17]), .ZN(n1721) );
  INV_X1 U1845 ( .A(n1379), .ZN(n1720) );
  OAI222_X1 U1846 ( .A1(n2085), .A2(n2086), .B1(n2085), .B2(n2087), .C1(n2087), 
        .C2(n2086), .ZN(n2081) );
  INV_X1 U1847 ( .A(n588), .ZN(n2087) );
  XNOR2_X1 U1848 ( .A(n1742), .B(n2088), .ZN(n2086) );
  AOI221_X1 U1849 ( .B1(b[18]), .B2(n1561), .C1(b[17]), .C2(n1562), .A(n2089), 
        .ZN(n2088) );
  OAI22_X1 U1850 ( .A1(n1564), .A2(n1716), .B1(n1639), .B2(n1717), .ZN(n2089)
         );
  INV_X1 U1851 ( .A(b[16]), .ZN(n1717) );
  INV_X1 U1852 ( .A(n1380), .ZN(n1716) );
  AOI222_X1 U1853 ( .A1(n2090), .A2(n2091), .B1(n2090), .B2(n600), .C1(n600), 
        .C2(n2091), .ZN(n2085) );
  XNOR2_X1 U1854 ( .A(a[2]), .B(n2092), .ZN(n2091) );
  AOI221_X1 U1855 ( .B1(b[17]), .B2(n1561), .C1(b[16]), .C2(n1562), .A(n2093), 
        .ZN(n2092) );
  OAI22_X1 U1856 ( .A1(n1564), .A2(n1712), .B1(n1639), .B2(n1713), .ZN(n2093)
         );
  INV_X1 U1857 ( .A(b[15]), .ZN(n1713) );
  INV_X1 U1858 ( .A(n1381), .ZN(n1712) );
  OAI222_X1 U1859 ( .A1(n2094), .A2(n2095), .B1(n2094), .B2(n2096), .C1(n2096), 
        .C2(n2095), .ZN(n2090) );
  INV_X1 U1860 ( .A(n610), .ZN(n2096) );
  XNOR2_X1 U1861 ( .A(n1742), .B(n2097), .ZN(n2095) );
  AOI221_X1 U1862 ( .B1(b[16]), .B2(n1561), .C1(b[15]), .C2(n1562), .A(n2098), 
        .ZN(n2097) );
  OAI22_X1 U1863 ( .A1(n1564), .A2(n1708), .B1(n1639), .B2(n1709), .ZN(n2098)
         );
  INV_X1 U1864 ( .A(b[14]), .ZN(n1709) );
  INV_X1 U1865 ( .A(n1382), .ZN(n1708) );
  AOI222_X1 U1866 ( .A1(n2099), .A2(n2100), .B1(n2099), .B2(n620), .C1(n620), 
        .C2(n2100), .ZN(n2094) );
  XNOR2_X1 U1867 ( .A(a[2]), .B(n2101), .ZN(n2100) );
  AOI221_X1 U1868 ( .B1(b[15]), .B2(n1561), .C1(b[14]), .C2(n1562), .A(n2102), 
        .ZN(n2101) );
  OAI22_X1 U1869 ( .A1(n1564), .A2(n1704), .B1(n1639), .B2(n1705), .ZN(n2102)
         );
  INV_X1 U1870 ( .A(b[13]), .ZN(n1705) );
  INV_X1 U1871 ( .A(n1383), .ZN(n1704) );
  OAI222_X1 U1872 ( .A1(n2103), .A2(n2104), .B1(n2103), .B2(n2105), .C1(n2105), 
        .C2(n2104), .ZN(n2099) );
  INV_X1 U1873 ( .A(n630), .ZN(n2105) );
  XNOR2_X1 U1874 ( .A(n1742), .B(n2106), .ZN(n2104) );
  AOI221_X1 U1875 ( .B1(b[14]), .B2(n1561), .C1(b[13]), .C2(n1562), .A(n2107), 
        .ZN(n2106) );
  OAI22_X1 U1876 ( .A1(n1564), .A2(n1700), .B1(n1639), .B2(n1701), .ZN(n2107)
         );
  INV_X1 U1877 ( .A(b[12]), .ZN(n1701) );
  INV_X1 U1878 ( .A(n1384), .ZN(n1700) );
  AOI222_X1 U1879 ( .A1(n2108), .A2(n2109), .B1(n2108), .B2(n638), .C1(n638), 
        .C2(n2109), .ZN(n2103) );
  XNOR2_X1 U1880 ( .A(a[2]), .B(n2110), .ZN(n2109) );
  AOI221_X1 U1881 ( .B1(b[13]), .B2(n1561), .C1(b[12]), .C2(n1562), .A(n2111), 
        .ZN(n2110) );
  OAI22_X1 U1882 ( .A1(n1564), .A2(n1696), .B1(n1639), .B2(n1697), .ZN(n2111)
         );
  INV_X1 U1883 ( .A(b[11]), .ZN(n1697) );
  INV_X1 U1884 ( .A(n1385), .ZN(n1696) );
  OAI222_X1 U1885 ( .A1(n2112), .A2(n2113), .B1(n2112), .B2(n2114), .C1(n2114), 
        .C2(n2113), .ZN(n2108) );
  INV_X1 U1886 ( .A(n646), .ZN(n2114) );
  XNOR2_X1 U1887 ( .A(n1742), .B(n2115), .ZN(n2113) );
  AOI221_X1 U1888 ( .B1(b[12]), .B2(n1561), .C1(b[11]), .C2(n1562), .A(n2116), 
        .ZN(n2115) );
  OAI22_X1 U1889 ( .A1(n1564), .A2(n1692), .B1(n1639), .B2(n1693), .ZN(n2116)
         );
  INV_X1 U1890 ( .A(b[10]), .ZN(n1693) );
  INV_X1 U1891 ( .A(n1386), .ZN(n1692) );
  AOI222_X1 U1892 ( .A1(n2117), .A2(n2118), .B1(n2117), .B2(n654), .C1(n654), 
        .C2(n2118), .ZN(n2112) );
  XNOR2_X1 U1893 ( .A(a[2]), .B(n2119), .ZN(n2118) );
  AOI221_X1 U1894 ( .B1(b[11]), .B2(n1561), .C1(b[10]), .C2(n1562), .A(n2120), 
        .ZN(n2119) );
  OAI22_X1 U1895 ( .A1(n1564), .A2(n1688), .B1(n1639), .B2(n1689), .ZN(n2120)
         );
  INV_X1 U1896 ( .A(b[9]), .ZN(n1689) );
  INV_X1 U1897 ( .A(n1387), .ZN(n1688) );
  OAI222_X1 U1898 ( .A1(n2121), .A2(n2122), .B1(n2121), .B2(n2123), .C1(n2123), 
        .C2(n2122), .ZN(n2117) );
  INV_X1 U1899 ( .A(n660), .ZN(n2123) );
  XNOR2_X1 U1900 ( .A(n1742), .B(n2124), .ZN(n2122) );
  AOI221_X1 U1901 ( .B1(b[10]), .B2(n1561), .C1(b[9]), .C2(n1563), .A(n2125), 
        .ZN(n2124) );
  OAI22_X1 U1902 ( .A1(n1564), .A2(n1684), .B1(n1639), .B2(n1685), .ZN(n2125)
         );
  INV_X1 U1903 ( .A(b[8]), .ZN(n1685) );
  INV_X1 U1904 ( .A(n1388), .ZN(n1684) );
  AOI222_X1 U1905 ( .A1(n2126), .A2(n2127), .B1(n2126), .B2(n666), .C1(n666), 
        .C2(n2127), .ZN(n2121) );
  XNOR2_X1 U1906 ( .A(a[2]), .B(n2128), .ZN(n2127) );
  AOI221_X1 U1907 ( .B1(b[9]), .B2(n1561), .C1(b[8]), .C2(n1563), .A(n2129), 
        .ZN(n2128) );
  OAI22_X1 U1908 ( .A1(n1564), .A2(n1680), .B1(n1639), .B2(n1681), .ZN(n2129)
         );
  INV_X1 U1909 ( .A(b[7]), .ZN(n1681) );
  INV_X1 U1910 ( .A(n1389), .ZN(n1680) );
  OAI222_X1 U1911 ( .A1(n2130), .A2(n2131), .B1(n2130), .B2(n2132), .C1(n2132), 
        .C2(n2131), .ZN(n2126) );
  INV_X1 U1912 ( .A(n672), .ZN(n2132) );
  XNOR2_X1 U1913 ( .A(n1742), .B(n2133), .ZN(n2131) );
  AOI221_X1 U1914 ( .B1(b[8]), .B2(n1561), .C1(b[7]), .C2(n1562), .A(n2134), 
        .ZN(n2133) );
  OAI22_X1 U1915 ( .A1(n1564), .A2(n1676), .B1(n1639), .B2(n1677), .ZN(n2134)
         );
  INV_X1 U1916 ( .A(b[6]), .ZN(n1677) );
  INV_X1 U1917 ( .A(n1390), .ZN(n1676) );
  AOI222_X1 U1918 ( .A1(n2135), .A2(n2136), .B1(n2135), .B2(n676), .C1(n676), 
        .C2(n2136), .ZN(n2130) );
  XNOR2_X1 U1919 ( .A(a[2]), .B(n2137), .ZN(n2136) );
  AOI221_X1 U1920 ( .B1(b[7]), .B2(n1561), .C1(b[6]), .C2(n1563), .A(n2138), 
        .ZN(n2137) );
  OAI22_X1 U1921 ( .A1(n1564), .A2(n1672), .B1(n1639), .B2(n1673), .ZN(n2138)
         );
  INV_X1 U1922 ( .A(b[5]), .ZN(n1673) );
  INV_X1 U1923 ( .A(n1391), .ZN(n1672) );
  OAI222_X1 U1924 ( .A1(n2139), .A2(n2140), .B1(n2139), .B2(n2141), .C1(n2141), 
        .C2(n2140), .ZN(n2135) );
  INV_X1 U1925 ( .A(n680), .ZN(n2141) );
  XNOR2_X1 U1926 ( .A(n1742), .B(n2142), .ZN(n2140) );
  AOI221_X1 U1927 ( .B1(b[6]), .B2(n1561), .C1(b[5]), .C2(n1563), .A(n2143), 
        .ZN(n2142) );
  OAI22_X1 U1928 ( .A1(n1564), .A2(n1668), .B1(n1639), .B2(n1669), .ZN(n2143)
         );
  INV_X1 U1929 ( .A(b[4]), .ZN(n1669) );
  INV_X1 U1930 ( .A(n1392), .ZN(n1668) );
  AOI222_X1 U1931 ( .A1(n2144), .A2(n2145), .B1(n2144), .B2(n684), .C1(n684), 
        .C2(n2145), .ZN(n2139) );
  XNOR2_X1 U1932 ( .A(a[2]), .B(n2146), .ZN(n2145) );
  AOI221_X1 U1933 ( .B1(b[5]), .B2(n1561), .C1(b[4]), .C2(n1563), .A(n2147), 
        .ZN(n2146) );
  OAI22_X1 U1934 ( .A1(n1564), .A2(n1664), .B1(n1639), .B2(n1665), .ZN(n2147)
         );
  INV_X1 U1935 ( .A(b[3]), .ZN(n1665) );
  INV_X1 U1936 ( .A(n1393), .ZN(n1664) );
  OAI222_X1 U1937 ( .A1(n2148), .A2(n2149), .B1(n2148), .B2(n2150), .C1(n2150), 
        .C2(n2149), .ZN(n2144) );
  INV_X1 U1938 ( .A(n686), .ZN(n2150) );
  XNOR2_X1 U1939 ( .A(n1742), .B(n2151), .ZN(n2149) );
  AOI221_X1 U1940 ( .B1(b[4]), .B2(n1561), .C1(b[3]), .C2(n1563), .A(n2152), 
        .ZN(n2151) );
  OAI22_X1 U1941 ( .A1(n1564), .A2(n1660), .B1(n1639), .B2(n1661), .ZN(n2152)
         );
  INV_X1 U1942 ( .A(n1394), .ZN(n1660) );
  AOI222_X1 U1943 ( .A1(n2153), .A2(n2154), .B1(n2153), .B2(n688), .C1(n688), 
        .C2(n2154), .ZN(n2148) );
  XNOR2_X1 U1944 ( .A(a[2]), .B(n2155), .ZN(n2154) );
  AOI221_X1 U1945 ( .B1(b[3]), .B2(n1561), .C1(b[2]), .C2(n1563), .A(n2156), 
        .ZN(n2155) );
  OAI22_X1 U1946 ( .A1(n1564), .A2(n1657), .B1(n1639), .B2(n1649), .ZN(n2156)
         );
  INV_X1 U1947 ( .A(b[1]), .ZN(n1649) );
  INV_X1 U1948 ( .A(n1395), .ZN(n1657) );
  AND2_X1 U1949 ( .A1(n2160), .A2(n2161), .ZN(n2153) );
  AOI211_X1 U1950 ( .C1(b[1]), .C2(n1561), .A(n2162), .B(b[0]), .ZN(n2161) );
  OAI22_X1 U1951 ( .A1(n1535), .A2(n1661), .B1(n1564), .B2(n1650), .ZN(n2162)
         );
  INV_X1 U1952 ( .A(n1397), .ZN(n1650) );
  INV_X1 U1953 ( .A(b[2]), .ZN(n1661) );
  INV_X1 U1954 ( .A(a[0]), .ZN(n2158) );
  AOI221_X1 U1955 ( .B1(b[1]), .B2(n1563), .C1(n1396), .C2(n1555), .A(n1742), 
        .ZN(n2160) );
  XNOR2_X1 U1956 ( .A(a[1]), .B(n1742), .ZN(n2157) );
  INV_X1 U1957 ( .A(a[2]), .ZN(n1742) );
  NOR2_X1 U1958 ( .A1(n2159), .A2(a[0]), .ZN(n1636) );
  INV_X1 U1959 ( .A(a[1]), .ZN(n2159) );
endmodule


module iir_filter_DW_mult_tc_4 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(product[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(product[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(product[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(product[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(product[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(product[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(product[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(product[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(product[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(product[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(product[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(product[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(product[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(product[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(product[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(product[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(product[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(product[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(product[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(product[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(product[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(product[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(product[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1598), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1600), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1602), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1604), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1606), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1608), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1610), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(b[22]), .B(n1615), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(b[21]), .B(b[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(b[20]), .B(b[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(b[19]), .B(b[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(b[18]), .B(b[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(b[17]), .B(b[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(b[16]), .B(b[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(b[15]), .B(b[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(b[14]), .B(b[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(b[13]), .B(b[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(b[12]), .B(b[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(b[11]), .B(b[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(b[10]), .B(b[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(b[9]), .B(b[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(b[8]), .B(b[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(b[7]), .B(b[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(b[6]), .B(b[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(b[5]), .B(b[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(b[4]), .B(b[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(b[3]), .B(b[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(b[2]), .B(b[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(b[1]), .B(b[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(b[0]), .B(b[1]), .CO(n727), .S(n1397) );
  INV_X1 U1137 ( .A(n1616), .ZN(n1615) );
  INV_X1 U1138 ( .A(n1533), .ZN(n1570) );
  INV_X1 U1139 ( .A(n1536), .ZN(n1568) );
  INV_X1 U1140 ( .A(n1535), .ZN(n1561) );
  INV_X1 U1141 ( .A(n1534), .ZN(n1569) );
  BUF_X1 U1142 ( .A(n1655), .Z(n1572) );
  INV_X1 U1143 ( .A(n1545), .ZN(n1560) );
  INV_X1 U1144 ( .A(n1543), .ZN(n1558) );
  INV_X1 U1145 ( .A(n1549), .ZN(n1580) );
  INV_X1 U1146 ( .A(n1550), .ZN(n1575) );
  INV_X1 U1147 ( .A(n1548), .ZN(n1585) );
  INV_X1 U1148 ( .A(n1546), .ZN(n1595) );
  INV_X1 U1149 ( .A(n1547), .ZN(n1590) );
  INV_X1 U1150 ( .A(n1537), .ZN(n1559) );
  INV_X1 U1151 ( .A(n1544), .ZN(n1593) );
  INV_X1 U1152 ( .A(n1552), .ZN(n1583) );
  INV_X1 U1153 ( .A(n1551), .ZN(n1588) );
  INV_X1 U1154 ( .A(n1553), .ZN(n1578) );
  INV_X1 U1155 ( .A(n1554), .ZN(n1573) );
  BUF_X1 U1156 ( .A(n1655), .Z(n1571) );
  BUF_X1 U1157 ( .A(n1630), .Z(n1557) );
  BUF_X1 U1158 ( .A(n1968), .Z(n1596) );
  BUF_X1 U1159 ( .A(n1913), .Z(n1591) );
  BUF_X1 U1160 ( .A(n1858), .Z(n1586) );
  BUF_X1 U1161 ( .A(n1803), .Z(n1581) );
  BUF_X1 U1162 ( .A(n1748), .Z(n1576) );
  BUF_X1 U1163 ( .A(n1913), .Z(n1592) );
  BUF_X1 U1164 ( .A(n1858), .Z(n1587) );
  BUF_X1 U1165 ( .A(n1803), .Z(n1582) );
  BUF_X1 U1166 ( .A(n1748), .Z(n1577) );
  BUF_X1 U1167 ( .A(n1968), .Z(n1597) );
  INV_X1 U1168 ( .A(n1539), .ZN(n1589) );
  INV_X1 U1169 ( .A(n1540), .ZN(n1584) );
  INV_X1 U1170 ( .A(n1541), .ZN(n1579) );
  INV_X1 U1171 ( .A(n1542), .ZN(n1574) );
  BUF_X1 U1172 ( .A(n1630), .Z(n1556) );
  INV_X1 U1173 ( .A(n1538), .ZN(n1594) );
  NAND3_X1 U1174 ( .A1(n2158), .A2(n2159), .A3(n2160), .ZN(n1640) );
  INV_X1 U1175 ( .A(n1555), .ZN(n1564) );
  OR2_X1 U1176 ( .A1(n1739), .A2(n1740), .ZN(n1533) );
  OR2_X1 U1177 ( .A1(n1741), .A2(n1742), .ZN(n1534) );
  OR2_X1 U1178 ( .A1(n2159), .A2(n2158), .ZN(n1535) );
  AND2_X1 U1179 ( .A1(n1739), .A2(n1741), .ZN(n1536) );
  INV_X1 U1180 ( .A(n1611), .ZN(n1610) );
  INV_X1 U1181 ( .A(n1607), .ZN(n1606) );
  INV_X1 U1182 ( .A(n1609), .ZN(n1608) );
  INV_X1 U1183 ( .A(n1605), .ZN(n1604) );
  INV_X1 U1184 ( .A(n1603), .ZN(n1602) );
  BUF_X1 U1185 ( .A(n1637), .Z(n1562) );
  BUF_X1 U1186 ( .A(n1637), .Z(n1563) );
  BUF_X1 U1187 ( .A(n1648), .Z(n1565) );
  BUF_X1 U1188 ( .A(n1648), .Z(n1566) );
  OR2_X1 U1189 ( .A1(n2069), .A2(n2068), .ZN(n1537) );
  OR2_X1 U1190 ( .A1(n2017), .A2(n2018), .ZN(n1538) );
  OR2_X1 U1191 ( .A1(n1962), .A2(n1963), .ZN(n1539) );
  OR2_X1 U1192 ( .A1(n1907), .A2(n1908), .ZN(n1540) );
  OR2_X1 U1193 ( .A1(n1852), .A2(n1853), .ZN(n1541) );
  OR2_X1 U1194 ( .A1(n1797), .A2(n1798), .ZN(n1542) );
  AND2_X1 U1195 ( .A1(n2071), .A2(n2069), .ZN(n1543) );
  AND2_X1 U1196 ( .A1(n2015), .A2(n2017), .ZN(n1544) );
  OR2_X1 U1197 ( .A1(n2071), .A2(n2070), .ZN(n1545) );
  OR2_X1 U1198 ( .A1(n2015), .A2(n2016), .ZN(n1546) );
  OR2_X1 U1199 ( .A1(n1960), .A2(n1961), .ZN(n1547) );
  OR2_X1 U1200 ( .A1(n1905), .A2(n1906), .ZN(n1548) );
  OR2_X1 U1201 ( .A1(n1850), .A2(n1851), .ZN(n1549) );
  OR2_X1 U1202 ( .A1(n1795), .A2(n1796), .ZN(n1550) );
  AND2_X1 U1203 ( .A1(n1960), .A2(n1962), .ZN(n1551) );
  AND2_X1 U1204 ( .A1(n1905), .A2(n1907), .ZN(n1552) );
  AND2_X1 U1205 ( .A1(n1850), .A2(n1852), .ZN(n1553) );
  AND2_X1 U1206 ( .A1(n1795), .A2(n1797), .ZN(n1554) );
  BUF_X1 U1207 ( .A(n1648), .Z(n1567) );
  INV_X1 U1208 ( .A(n1599), .ZN(n1598) );
  AND2_X1 U1209 ( .A1(a[0]), .A2(n2158), .ZN(n1555) );
  BUF_X1 U1210 ( .A(a[20]), .Z(n1600) );
  INV_X1 U1211 ( .A(a[23]), .ZN(n1599) );
  INV_X1 U1212 ( .A(a[5]), .ZN(n1611) );
  INV_X1 U1213 ( .A(a[11]), .ZN(n1607) );
  INV_X1 U1214 ( .A(a[8]), .ZN(n1609) );
  INV_X1 U1215 ( .A(a[14]), .ZN(n1605) );
  INV_X1 U1216 ( .A(a[17]), .ZN(n1603) );
  BUF_X1 U1217 ( .A(a[20]), .Z(n1601) );
  CLKBUF_X1 U1218 ( .A(b[23]), .Z(n1612) );
  CLKBUF_X1 U1219 ( .A(b[23]), .Z(n1613) );
  CLKBUF_X1 U1220 ( .A(b[23]), .Z(n1614) );
  INV_X1 U1221 ( .A(n1612), .ZN(n1616) );
  INV_X1 U1222 ( .A(n1612), .ZN(n1617) );
  INV_X1 U1223 ( .A(n1613), .ZN(n1618) );
  INV_X1 U1224 ( .A(n1613), .ZN(n1619) );
  INV_X1 U1225 ( .A(n1614), .ZN(n1620) );
  INV_X1 U1226 ( .A(n1614), .ZN(n1621) );
  AOI21_X1 U1227 ( .B1(n1622), .B2(n1623), .A(n1624), .ZN(product[47]) );
  OAI22_X1 U1228 ( .A1(n1625), .A2(n1626), .B1(n1625), .B2(n1627), .ZN(n1624)
         );
  INV_X1 U1229 ( .A(n1623), .ZN(n1627) );
  AOI222_X1 U1230 ( .A1(n1628), .A2(n303), .B1(n1626), .B2(n303), .C1(n1628), 
        .C2(n1626), .ZN(n1625) );
  XOR2_X1 U1231 ( .A(n1629), .B(n1599), .Z(n1623) );
  OAI221_X1 U1232 ( .B1(n1617), .B2(n1557), .C1(n1621), .C2(n1558), .A(n1631), 
        .ZN(n1629) );
  OAI21_X1 U1233 ( .B1(n1559), .B2(n1560), .A(n1615), .ZN(n1631) );
  INV_X1 U1234 ( .A(n1626), .ZN(n1622) );
  XOR2_X1 U1235 ( .A(a[23]), .B(n1632), .Z(n1626) );
  AOI221_X1 U1236 ( .B1(n1614), .B2(n1559), .C1(n1560), .C2(n1615), .A(n1633), 
        .ZN(n1632) );
  OAI22_X1 U1237 ( .A1(n1558), .A2(n1634), .B1(n1557), .B2(n1635), .ZN(n1633)
         );
  XNOR2_X1 U1238 ( .A(a[2]), .B(n1636), .ZN(n908) );
  AOI221_X1 U1239 ( .B1(n1561), .B2(b[22]), .C1(n1563), .C2(b[21]), .A(n1638), 
        .ZN(n1636) );
  OAI22_X1 U1240 ( .A1(n1564), .A2(n1639), .B1(n1640), .B2(n1641), .ZN(n1638)
         );
  INV_X1 U1241 ( .A(n1376), .ZN(n1639) );
  XNOR2_X1 U1242 ( .A(a[2]), .B(n1642), .ZN(n907) );
  AOI221_X1 U1243 ( .B1(n1563), .B2(b[22]), .C1(n1555), .C2(n1375), .A(n1643), 
        .ZN(n1642) );
  OAI22_X1 U1244 ( .A1(n1644), .A2(n1640), .B1(n1617), .B2(n1535), .ZN(n1643)
         );
  XNOR2_X1 U1245 ( .A(a[2]), .B(n1645), .ZN(n906) );
  AOI221_X1 U1246 ( .B1(n1561), .B2(n1614), .C1(n1563), .C2(n1615), .A(n1646), 
        .ZN(n1645) );
  OAI22_X1 U1247 ( .A1(n1634), .A2(n1564), .B1(n1635), .B2(n1640), .ZN(n1646)
         );
  XNOR2_X1 U1248 ( .A(n1647), .B(n1611), .ZN(n904) );
  OAI22_X1 U1249 ( .A1(n1565), .A2(n1534), .B1(n1568), .B2(n1567), .ZN(n1647)
         );
  XNOR2_X1 U1250 ( .A(n1649), .B(n1611), .ZN(n903) );
  OAI222_X1 U1251 ( .A1(n1534), .A2(n1650), .B1(n1566), .B2(n1533), .C1(n1568), 
        .C2(n1651), .ZN(n1649) );
  XNOR2_X1 U1252 ( .A(n1610), .B(n1652), .ZN(n902) );
  AOI221_X1 U1253 ( .B1(b[2]), .B2(n1569), .C1(b[1]), .C2(n1570), .A(n1653), 
        .ZN(n1652) );
  OAI22_X1 U1254 ( .A1(n1568), .A2(n1654), .B1(n1565), .B2(n1572), .ZN(n1653)
         );
  XNOR2_X1 U1255 ( .A(n1610), .B(n1656), .ZN(n901) );
  AOI221_X1 U1256 ( .B1(b[3]), .B2(n1569), .C1(b[2]), .C2(n1570), .A(n1657), 
        .ZN(n1656) );
  OAI22_X1 U1257 ( .A1(n1568), .A2(n1658), .B1(n1650), .B2(n1572), .ZN(n1657)
         );
  XNOR2_X1 U1258 ( .A(n1610), .B(n1659), .ZN(n900) );
  AOI221_X1 U1259 ( .B1(b[4]), .B2(n1569), .C1(b[3]), .C2(n1570), .A(n1660), 
        .ZN(n1659) );
  OAI22_X1 U1260 ( .A1(n1568), .A2(n1661), .B1(n1662), .B2(n1572), .ZN(n1660)
         );
  XNOR2_X1 U1261 ( .A(n1610), .B(n1663), .ZN(n899) );
  AOI221_X1 U1262 ( .B1(b[5]), .B2(n1569), .C1(b[4]), .C2(n1570), .A(n1664), 
        .ZN(n1663) );
  OAI22_X1 U1263 ( .A1(n1568), .A2(n1665), .B1(n1572), .B2(n1666), .ZN(n1664)
         );
  XNOR2_X1 U1264 ( .A(n1610), .B(n1667), .ZN(n898) );
  AOI221_X1 U1265 ( .B1(b[6]), .B2(n1569), .C1(b[5]), .C2(n1570), .A(n1668), 
        .ZN(n1667) );
  OAI22_X1 U1266 ( .A1(n1568), .A2(n1669), .B1(n1572), .B2(n1670), .ZN(n1668)
         );
  XNOR2_X1 U1267 ( .A(n1610), .B(n1671), .ZN(n897) );
  AOI221_X1 U1268 ( .B1(b[7]), .B2(n1569), .C1(b[6]), .C2(n1570), .A(n1672), 
        .ZN(n1671) );
  OAI22_X1 U1269 ( .A1(n1568), .A2(n1673), .B1(n1572), .B2(n1674), .ZN(n1672)
         );
  XNOR2_X1 U1270 ( .A(n1610), .B(n1675), .ZN(n896) );
  AOI221_X1 U1271 ( .B1(b[8]), .B2(n1569), .C1(b[7]), .C2(n1570), .A(n1676), 
        .ZN(n1675) );
  OAI22_X1 U1272 ( .A1(n1568), .A2(n1677), .B1(n1571), .B2(n1678), .ZN(n1676)
         );
  XNOR2_X1 U1273 ( .A(n1610), .B(n1679), .ZN(n895) );
  AOI221_X1 U1274 ( .B1(b[9]), .B2(n1569), .C1(b[8]), .C2(n1570), .A(n1680), 
        .ZN(n1679) );
  OAI22_X1 U1275 ( .A1(n1568), .A2(n1681), .B1(n1572), .B2(n1682), .ZN(n1680)
         );
  XNOR2_X1 U1276 ( .A(n1610), .B(n1683), .ZN(n894) );
  AOI221_X1 U1277 ( .B1(b[10]), .B2(n1569), .C1(b[9]), .C2(n1570), .A(n1684), 
        .ZN(n1683) );
  OAI22_X1 U1278 ( .A1(n1568), .A2(n1685), .B1(n1572), .B2(n1686), .ZN(n1684)
         );
  XNOR2_X1 U1279 ( .A(n1610), .B(n1687), .ZN(n893) );
  AOI221_X1 U1280 ( .B1(b[11]), .B2(n1569), .C1(b[10]), .C2(n1570), .A(n1688), 
        .ZN(n1687) );
  OAI22_X1 U1281 ( .A1(n1568), .A2(n1689), .B1(n1571), .B2(n1690), .ZN(n1688)
         );
  XNOR2_X1 U1282 ( .A(n1610), .B(n1691), .ZN(n892) );
  AOI221_X1 U1283 ( .B1(b[12]), .B2(n1569), .C1(b[11]), .C2(n1570), .A(n1692), 
        .ZN(n1691) );
  OAI22_X1 U1284 ( .A1(n1568), .A2(n1693), .B1(n1571), .B2(n1694), .ZN(n1692)
         );
  XNOR2_X1 U1285 ( .A(n1610), .B(n1695), .ZN(n891) );
  AOI221_X1 U1286 ( .B1(b[13]), .B2(n1569), .C1(b[12]), .C2(n1570), .A(n1696), 
        .ZN(n1695) );
  OAI22_X1 U1287 ( .A1(n1568), .A2(n1697), .B1(n1571), .B2(n1698), .ZN(n1696)
         );
  XNOR2_X1 U1288 ( .A(n1610), .B(n1699), .ZN(n890) );
  AOI221_X1 U1289 ( .B1(b[14]), .B2(n1569), .C1(b[13]), .C2(n1570), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U1290 ( .A1(n1568), .A2(n1701), .B1(n1571), .B2(n1702), .ZN(n1700)
         );
  XNOR2_X1 U1291 ( .A(n1610), .B(n1703), .ZN(n889) );
  AOI221_X1 U1292 ( .B1(b[15]), .B2(n1569), .C1(b[14]), .C2(n1570), .A(n1704), 
        .ZN(n1703) );
  OAI22_X1 U1293 ( .A1(n1568), .A2(n1705), .B1(n1571), .B2(n1706), .ZN(n1704)
         );
  XNOR2_X1 U1294 ( .A(n1610), .B(n1707), .ZN(n888) );
  AOI221_X1 U1295 ( .B1(b[16]), .B2(n1569), .C1(b[15]), .C2(n1570), .A(n1708), 
        .ZN(n1707) );
  OAI22_X1 U1296 ( .A1(n1568), .A2(n1709), .B1(n1571), .B2(n1710), .ZN(n1708)
         );
  XNOR2_X1 U1297 ( .A(n1610), .B(n1711), .ZN(n887) );
  AOI221_X1 U1298 ( .B1(b[17]), .B2(n1569), .C1(b[16]), .C2(n1570), .A(n1712), 
        .ZN(n1711) );
  OAI22_X1 U1299 ( .A1(n1568), .A2(n1713), .B1(n1571), .B2(n1714), .ZN(n1712)
         );
  XNOR2_X1 U1300 ( .A(n1610), .B(n1715), .ZN(n886) );
  AOI221_X1 U1301 ( .B1(b[18]), .B2(n1569), .C1(b[17]), .C2(n1570), .A(n1716), 
        .ZN(n1715) );
  OAI22_X1 U1302 ( .A1(n1568), .A2(n1717), .B1(n1571), .B2(n1718), .ZN(n1716)
         );
  XNOR2_X1 U1303 ( .A(n1610), .B(n1719), .ZN(n885) );
  AOI221_X1 U1304 ( .B1(b[19]), .B2(n1569), .C1(b[18]), .C2(n1570), .A(n1720), 
        .ZN(n1719) );
  OAI22_X1 U1305 ( .A1(n1568), .A2(n1721), .B1(n1571), .B2(n1722), .ZN(n1720)
         );
  XNOR2_X1 U1306 ( .A(a[5]), .B(n1723), .ZN(n884) );
  AOI221_X1 U1307 ( .B1(n1569), .B2(b[20]), .C1(b[19]), .C2(n1570), .A(n1724), 
        .ZN(n1723) );
  OAI22_X1 U1308 ( .A1(n1568), .A2(n1725), .B1(n1571), .B2(n1726), .ZN(n1724)
         );
  XNOR2_X1 U1309 ( .A(a[5]), .B(n1727), .ZN(n883) );
  AOI221_X1 U1310 ( .B1(n1569), .B2(b[21]), .C1(n1570), .C2(b[20]), .A(n1728), 
        .ZN(n1727) );
  OAI22_X1 U1311 ( .A1(n1568), .A2(n1729), .B1(n1571), .B2(n1730), .ZN(n1728)
         );
  XNOR2_X1 U1312 ( .A(a[5]), .B(n1731), .ZN(n882) );
  AOI221_X1 U1313 ( .B1(n1569), .B2(b[22]), .C1(n1536), .C2(n1376), .A(n1732), 
        .ZN(n1731) );
  OAI22_X1 U1314 ( .A1(n1641), .A2(n1572), .B1(n1644), .B2(n1533), .ZN(n1732)
         );
  XNOR2_X1 U1315 ( .A(a[5]), .B(n1733), .ZN(n881) );
  AOI221_X1 U1316 ( .B1(n1570), .B2(b[22]), .C1(n1536), .C2(n1375), .A(n1734), 
        .ZN(n1733) );
  OAI22_X1 U1317 ( .A1(n1616), .A2(n1534), .B1(n1644), .B2(n1572), .ZN(n1734)
         );
  XNOR2_X1 U1318 ( .A(a[5]), .B(n1735), .ZN(n880) );
  AOI221_X1 U1319 ( .B1(n1569), .B2(n1614), .C1(n1570), .C2(n1615), .A(n1736), 
        .ZN(n1735) );
  OAI22_X1 U1320 ( .A1(n1634), .A2(n1568), .B1(n1635), .B2(n1572), .ZN(n1736)
         );
  XNOR2_X1 U1321 ( .A(n1610), .B(n1737), .ZN(n879) );
  OAI221_X1 U1322 ( .B1(n1618), .B2(n1572), .C1(n1621), .C2(n1568), .A(n1738), 
        .ZN(n1737) );
  OAI21_X1 U1323 ( .B1(n1569), .B2(n1570), .A(n1615), .ZN(n1738) );
  INV_X1 U1324 ( .A(n1742), .ZN(n1739) );
  NAND3_X1 U1325 ( .A1(n1742), .A2(n1741), .A3(n1740), .ZN(n1655) );
  XNOR2_X1 U1326 ( .A(a[3]), .B(a[4]), .ZN(n1740) );
  XNOR2_X1 U1327 ( .A(a[4]), .B(n1611), .ZN(n1741) );
  XOR2_X1 U1328 ( .A(a[3]), .B(n1743), .Z(n1742) );
  XNOR2_X1 U1329 ( .A(n1744), .B(n1609), .ZN(n878) );
  OAI22_X1 U1330 ( .A1(n1565), .A2(n1542), .B1(n1565), .B2(n1573), .ZN(n1744)
         );
  XNOR2_X1 U1331 ( .A(n1745), .B(n1609), .ZN(n877) );
  OAI222_X1 U1332 ( .A1(n1650), .A2(n1542), .B1(n1566), .B2(n1550), .C1(n1651), 
        .C2(n1573), .ZN(n1745) );
  XNOR2_X1 U1333 ( .A(n1608), .B(n1746), .ZN(n876) );
  AOI221_X1 U1334 ( .B1(n1574), .B2(b[2]), .C1(n1575), .C2(b[1]), .A(n1747), 
        .ZN(n1746) );
  OAI22_X1 U1335 ( .A1(n1654), .A2(n1573), .B1(n1565), .B2(n1576), .ZN(n1747)
         );
  XNOR2_X1 U1336 ( .A(n1608), .B(n1749), .ZN(n875) );
  AOI221_X1 U1337 ( .B1(n1574), .B2(b[3]), .C1(n1575), .C2(b[2]), .A(n1750), 
        .ZN(n1749) );
  OAI22_X1 U1338 ( .A1(n1658), .A2(n1573), .B1(n1650), .B2(n1577), .ZN(n1750)
         );
  XNOR2_X1 U1339 ( .A(n1608), .B(n1751), .ZN(n874) );
  AOI221_X1 U1340 ( .B1(n1574), .B2(b[4]), .C1(n1575), .C2(b[3]), .A(n1752), 
        .ZN(n1751) );
  OAI22_X1 U1341 ( .A1(n1661), .A2(n1573), .B1(n1662), .B2(n1577), .ZN(n1752)
         );
  XNOR2_X1 U1342 ( .A(n1608), .B(n1753), .ZN(n873) );
  AOI221_X1 U1343 ( .B1(n1574), .B2(b[5]), .C1(n1575), .C2(b[4]), .A(n1754), 
        .ZN(n1753) );
  OAI22_X1 U1344 ( .A1(n1665), .A2(n1573), .B1(n1666), .B2(n1577), .ZN(n1754)
         );
  XNOR2_X1 U1345 ( .A(n1608), .B(n1755), .ZN(n872) );
  AOI221_X1 U1346 ( .B1(n1574), .B2(b[6]), .C1(n1575), .C2(b[5]), .A(n1756), 
        .ZN(n1755) );
  OAI22_X1 U1347 ( .A1(n1669), .A2(n1573), .B1(n1670), .B2(n1577), .ZN(n1756)
         );
  XNOR2_X1 U1348 ( .A(n1608), .B(n1757), .ZN(n871) );
  AOI221_X1 U1349 ( .B1(n1574), .B2(b[7]), .C1(n1575), .C2(b[6]), .A(n1758), 
        .ZN(n1757) );
  OAI22_X1 U1350 ( .A1(n1673), .A2(n1573), .B1(n1674), .B2(n1577), .ZN(n1758)
         );
  XNOR2_X1 U1351 ( .A(n1608), .B(n1759), .ZN(n870) );
  AOI221_X1 U1352 ( .B1(n1574), .B2(b[8]), .C1(n1575), .C2(b[7]), .A(n1760), 
        .ZN(n1759) );
  OAI22_X1 U1353 ( .A1(n1677), .A2(n1573), .B1(n1678), .B2(n1577), .ZN(n1760)
         );
  XNOR2_X1 U1354 ( .A(n1608), .B(n1761), .ZN(n869) );
  AOI221_X1 U1355 ( .B1(n1574), .B2(b[9]), .C1(n1575), .C2(b[8]), .A(n1762), 
        .ZN(n1761) );
  OAI22_X1 U1356 ( .A1(n1681), .A2(n1573), .B1(n1682), .B2(n1577), .ZN(n1762)
         );
  XNOR2_X1 U1357 ( .A(n1608), .B(n1763), .ZN(n868) );
  AOI221_X1 U1358 ( .B1(n1574), .B2(b[10]), .C1(n1575), .C2(b[9]), .A(n1764), 
        .ZN(n1763) );
  OAI22_X1 U1359 ( .A1(n1685), .A2(n1573), .B1(n1686), .B2(n1577), .ZN(n1764)
         );
  XNOR2_X1 U1360 ( .A(n1608), .B(n1765), .ZN(n867) );
  AOI221_X1 U1361 ( .B1(n1574), .B2(b[11]), .C1(n1575), .C2(b[10]), .A(n1766), 
        .ZN(n1765) );
  OAI22_X1 U1362 ( .A1(n1689), .A2(n1573), .B1(n1690), .B2(n1577), .ZN(n1766)
         );
  XNOR2_X1 U1363 ( .A(n1608), .B(n1767), .ZN(n866) );
  AOI221_X1 U1364 ( .B1(n1574), .B2(b[12]), .C1(n1575), .C2(b[11]), .A(n1768), 
        .ZN(n1767) );
  OAI22_X1 U1365 ( .A1(n1693), .A2(n1573), .B1(n1694), .B2(n1577), .ZN(n1768)
         );
  XNOR2_X1 U1366 ( .A(n1608), .B(n1769), .ZN(n865) );
  AOI221_X1 U1367 ( .B1(n1574), .B2(b[13]), .C1(n1575), .C2(b[12]), .A(n1770), 
        .ZN(n1769) );
  OAI22_X1 U1368 ( .A1(n1697), .A2(n1573), .B1(n1698), .B2(n1576), .ZN(n1770)
         );
  XNOR2_X1 U1369 ( .A(n1608), .B(n1771), .ZN(n864) );
  AOI221_X1 U1370 ( .B1(n1574), .B2(b[14]), .C1(n1575), .C2(b[13]), .A(n1772), 
        .ZN(n1771) );
  OAI22_X1 U1371 ( .A1(n1701), .A2(n1573), .B1(n1702), .B2(n1576), .ZN(n1772)
         );
  XNOR2_X1 U1372 ( .A(n1608), .B(n1773), .ZN(n863) );
  AOI221_X1 U1373 ( .B1(n1574), .B2(b[15]), .C1(n1575), .C2(b[14]), .A(n1774), 
        .ZN(n1773) );
  OAI22_X1 U1374 ( .A1(n1705), .A2(n1573), .B1(n1706), .B2(n1576), .ZN(n1774)
         );
  XNOR2_X1 U1375 ( .A(n1608), .B(n1775), .ZN(n862) );
  AOI221_X1 U1376 ( .B1(n1574), .B2(b[16]), .C1(n1575), .C2(b[15]), .A(n1776), 
        .ZN(n1775) );
  OAI22_X1 U1377 ( .A1(n1709), .A2(n1573), .B1(n1710), .B2(n1576), .ZN(n1776)
         );
  XNOR2_X1 U1378 ( .A(n1608), .B(n1777), .ZN(n861) );
  AOI221_X1 U1379 ( .B1(n1574), .B2(b[17]), .C1(n1575), .C2(b[16]), .A(n1778), 
        .ZN(n1777) );
  OAI22_X1 U1380 ( .A1(n1713), .A2(n1573), .B1(n1714), .B2(n1576), .ZN(n1778)
         );
  XNOR2_X1 U1381 ( .A(n1608), .B(n1779), .ZN(n860) );
  AOI221_X1 U1382 ( .B1(n1574), .B2(b[18]), .C1(n1575), .C2(b[17]), .A(n1780), 
        .ZN(n1779) );
  OAI22_X1 U1383 ( .A1(n1717), .A2(n1573), .B1(n1718), .B2(n1576), .ZN(n1780)
         );
  XNOR2_X1 U1384 ( .A(n1608), .B(n1781), .ZN(n859) );
  AOI221_X1 U1385 ( .B1(n1574), .B2(b[19]), .C1(n1575), .C2(b[18]), .A(n1782), 
        .ZN(n1781) );
  OAI22_X1 U1386 ( .A1(n1721), .A2(n1573), .B1(n1722), .B2(n1576), .ZN(n1782)
         );
  XNOR2_X1 U1387 ( .A(a[8]), .B(n1783), .ZN(n858) );
  AOI221_X1 U1388 ( .B1(n1574), .B2(b[20]), .C1(n1575), .C2(b[19]), .A(n1784), 
        .ZN(n1783) );
  OAI22_X1 U1389 ( .A1(n1725), .A2(n1573), .B1(n1726), .B2(n1576), .ZN(n1784)
         );
  XNOR2_X1 U1390 ( .A(a[8]), .B(n1785), .ZN(n857) );
  AOI221_X1 U1391 ( .B1(n1574), .B2(b[21]), .C1(n1575), .C2(b[20]), .A(n1786), 
        .ZN(n1785) );
  OAI22_X1 U1392 ( .A1(n1729), .A2(n1573), .B1(n1730), .B2(n1576), .ZN(n1786)
         );
  XNOR2_X1 U1393 ( .A(a[8]), .B(n1787), .ZN(n856) );
  AOI221_X1 U1394 ( .B1(n1574), .B2(b[22]), .C1(n1554), .C2(n1376), .A(n1788), 
        .ZN(n1787) );
  OAI22_X1 U1395 ( .A1(n1641), .A2(n1577), .B1(n1644), .B2(n1550), .ZN(n1788)
         );
  XNOR2_X1 U1396 ( .A(a[8]), .B(n1789), .ZN(n855) );
  AOI221_X1 U1397 ( .B1(n1575), .B2(b[22]), .C1(n1554), .C2(n1375), .A(n1790), 
        .ZN(n1789) );
  OAI22_X1 U1398 ( .A1(n1617), .A2(n1542), .B1(n1644), .B2(n1576), .ZN(n1790)
         );
  XNOR2_X1 U1399 ( .A(a[8]), .B(n1791), .ZN(n854) );
  AOI221_X1 U1400 ( .B1(n1574), .B2(n1614), .C1(n1575), .C2(n1615), .A(n1792), 
        .ZN(n1791) );
  OAI22_X1 U1401 ( .A1(n1634), .A2(n1573), .B1(n1635), .B2(n1576), .ZN(n1792)
         );
  XNOR2_X1 U1402 ( .A(n1608), .B(n1793), .ZN(n853) );
  OAI221_X1 U1403 ( .B1(n1618), .B2(n1577), .C1(n1617), .C2(n1573), .A(n1794), 
        .ZN(n1793) );
  OAI21_X1 U1404 ( .B1(n1574), .B2(n1575), .A(n1615), .ZN(n1794) );
  INV_X1 U1405 ( .A(n1798), .ZN(n1795) );
  NAND3_X1 U1406 ( .A1(n1798), .A2(n1797), .A3(n1796), .ZN(n1748) );
  XNOR2_X1 U1407 ( .A(a[6]), .B(a[7]), .ZN(n1796) );
  XNOR2_X1 U1408 ( .A(a[7]), .B(n1609), .ZN(n1797) );
  XOR2_X1 U1409 ( .A(a[6]), .B(n1611), .Z(n1798) );
  XNOR2_X1 U1410 ( .A(n1799), .B(n1607), .ZN(n852) );
  OAI22_X1 U1411 ( .A1(n1565), .A2(n1541), .B1(n1565), .B2(n1578), .ZN(n1799)
         );
  XNOR2_X1 U1412 ( .A(n1800), .B(n1607), .ZN(n851) );
  OAI222_X1 U1413 ( .A1(n1650), .A2(n1541), .B1(n1566), .B2(n1549), .C1(n1651), 
        .C2(n1578), .ZN(n1800) );
  XNOR2_X1 U1414 ( .A(n1606), .B(n1801), .ZN(n850) );
  AOI221_X1 U1415 ( .B1(n1579), .B2(b[2]), .C1(n1580), .C2(b[1]), .A(n1802), 
        .ZN(n1801) );
  OAI22_X1 U1416 ( .A1(n1654), .A2(n1578), .B1(n1566), .B2(n1581), .ZN(n1802)
         );
  XNOR2_X1 U1417 ( .A(n1606), .B(n1804), .ZN(n849) );
  AOI221_X1 U1418 ( .B1(n1579), .B2(b[3]), .C1(n1580), .C2(b[2]), .A(n1805), 
        .ZN(n1804) );
  OAI22_X1 U1419 ( .A1(n1658), .A2(n1578), .B1(n1650), .B2(n1582), .ZN(n1805)
         );
  XNOR2_X1 U1420 ( .A(n1606), .B(n1806), .ZN(n848) );
  AOI221_X1 U1421 ( .B1(n1579), .B2(b[4]), .C1(n1580), .C2(b[3]), .A(n1807), 
        .ZN(n1806) );
  OAI22_X1 U1422 ( .A1(n1661), .A2(n1578), .B1(n1662), .B2(n1582), .ZN(n1807)
         );
  XNOR2_X1 U1423 ( .A(n1606), .B(n1808), .ZN(n847) );
  AOI221_X1 U1424 ( .B1(n1579), .B2(b[5]), .C1(n1580), .C2(b[4]), .A(n1809), 
        .ZN(n1808) );
  OAI22_X1 U1425 ( .A1(n1665), .A2(n1578), .B1(n1666), .B2(n1582), .ZN(n1809)
         );
  XNOR2_X1 U1426 ( .A(n1606), .B(n1810), .ZN(n846) );
  AOI221_X1 U1427 ( .B1(n1579), .B2(b[6]), .C1(n1580), .C2(b[5]), .A(n1811), 
        .ZN(n1810) );
  OAI22_X1 U1428 ( .A1(n1669), .A2(n1578), .B1(n1670), .B2(n1582), .ZN(n1811)
         );
  XNOR2_X1 U1429 ( .A(n1606), .B(n1812), .ZN(n845) );
  AOI221_X1 U1430 ( .B1(n1579), .B2(b[7]), .C1(n1580), .C2(b[6]), .A(n1813), 
        .ZN(n1812) );
  OAI22_X1 U1431 ( .A1(n1673), .A2(n1578), .B1(n1674), .B2(n1582), .ZN(n1813)
         );
  XNOR2_X1 U1432 ( .A(n1606), .B(n1814), .ZN(n844) );
  AOI221_X1 U1433 ( .B1(n1579), .B2(b[8]), .C1(n1580), .C2(b[7]), .A(n1815), 
        .ZN(n1814) );
  OAI22_X1 U1434 ( .A1(n1677), .A2(n1578), .B1(n1678), .B2(n1582), .ZN(n1815)
         );
  XNOR2_X1 U1435 ( .A(n1606), .B(n1816), .ZN(n843) );
  AOI221_X1 U1436 ( .B1(n1579), .B2(b[9]), .C1(n1580), .C2(b[8]), .A(n1817), 
        .ZN(n1816) );
  OAI22_X1 U1437 ( .A1(n1681), .A2(n1578), .B1(n1682), .B2(n1582), .ZN(n1817)
         );
  XNOR2_X1 U1438 ( .A(n1606), .B(n1818), .ZN(n842) );
  AOI221_X1 U1439 ( .B1(n1579), .B2(b[10]), .C1(n1580), .C2(b[9]), .A(n1819), 
        .ZN(n1818) );
  OAI22_X1 U1440 ( .A1(n1685), .A2(n1578), .B1(n1686), .B2(n1582), .ZN(n1819)
         );
  XNOR2_X1 U1441 ( .A(n1606), .B(n1820), .ZN(n841) );
  AOI221_X1 U1442 ( .B1(n1579), .B2(b[11]), .C1(n1580), .C2(b[10]), .A(n1821), 
        .ZN(n1820) );
  OAI22_X1 U1443 ( .A1(n1689), .A2(n1578), .B1(n1690), .B2(n1582), .ZN(n1821)
         );
  XNOR2_X1 U1444 ( .A(n1606), .B(n1822), .ZN(n840) );
  AOI221_X1 U1445 ( .B1(n1579), .B2(b[12]), .C1(n1580), .C2(b[11]), .A(n1823), 
        .ZN(n1822) );
  OAI22_X1 U1446 ( .A1(n1693), .A2(n1578), .B1(n1694), .B2(n1582), .ZN(n1823)
         );
  XNOR2_X1 U1447 ( .A(n1606), .B(n1824), .ZN(n839) );
  AOI221_X1 U1448 ( .B1(n1579), .B2(b[13]), .C1(n1580), .C2(b[12]), .A(n1825), 
        .ZN(n1824) );
  OAI22_X1 U1449 ( .A1(n1697), .A2(n1578), .B1(n1698), .B2(n1581), .ZN(n1825)
         );
  XNOR2_X1 U1450 ( .A(n1606), .B(n1826), .ZN(n838) );
  AOI221_X1 U1451 ( .B1(n1579), .B2(b[14]), .C1(n1580), .C2(b[13]), .A(n1827), 
        .ZN(n1826) );
  OAI22_X1 U1452 ( .A1(n1701), .A2(n1578), .B1(n1702), .B2(n1581), .ZN(n1827)
         );
  XNOR2_X1 U1453 ( .A(n1606), .B(n1828), .ZN(n837) );
  AOI221_X1 U1454 ( .B1(n1579), .B2(b[15]), .C1(n1580), .C2(b[14]), .A(n1829), 
        .ZN(n1828) );
  OAI22_X1 U1455 ( .A1(n1705), .A2(n1578), .B1(n1706), .B2(n1581), .ZN(n1829)
         );
  XNOR2_X1 U1456 ( .A(n1606), .B(n1830), .ZN(n836) );
  AOI221_X1 U1457 ( .B1(n1579), .B2(b[16]), .C1(n1580), .C2(b[15]), .A(n1831), 
        .ZN(n1830) );
  OAI22_X1 U1458 ( .A1(n1709), .A2(n1578), .B1(n1710), .B2(n1581), .ZN(n1831)
         );
  XNOR2_X1 U1459 ( .A(n1606), .B(n1832), .ZN(n835) );
  AOI221_X1 U1460 ( .B1(n1579), .B2(b[17]), .C1(n1580), .C2(b[16]), .A(n1833), 
        .ZN(n1832) );
  OAI22_X1 U1461 ( .A1(n1713), .A2(n1578), .B1(n1714), .B2(n1581), .ZN(n1833)
         );
  XNOR2_X1 U1462 ( .A(n1606), .B(n1834), .ZN(n834) );
  AOI221_X1 U1463 ( .B1(n1579), .B2(b[18]), .C1(n1580), .C2(b[17]), .A(n1835), 
        .ZN(n1834) );
  OAI22_X1 U1464 ( .A1(n1717), .A2(n1578), .B1(n1718), .B2(n1581), .ZN(n1835)
         );
  XNOR2_X1 U1465 ( .A(n1606), .B(n1836), .ZN(n833) );
  AOI221_X1 U1466 ( .B1(n1579), .B2(b[19]), .C1(n1580), .C2(b[18]), .A(n1837), 
        .ZN(n1836) );
  OAI22_X1 U1467 ( .A1(n1721), .A2(n1578), .B1(n1722), .B2(n1581), .ZN(n1837)
         );
  XNOR2_X1 U1468 ( .A(n1606), .B(n1838), .ZN(n832) );
  AOI221_X1 U1469 ( .B1(n1579), .B2(b[20]), .C1(n1580), .C2(b[19]), .A(n1839), 
        .ZN(n1838) );
  OAI22_X1 U1470 ( .A1(n1725), .A2(n1578), .B1(n1726), .B2(n1581), .ZN(n1839)
         );
  XNOR2_X1 U1471 ( .A(a[11]), .B(n1840), .ZN(n831) );
  AOI221_X1 U1472 ( .B1(n1579), .B2(b[21]), .C1(n1580), .C2(b[20]), .A(n1841), 
        .ZN(n1840) );
  OAI22_X1 U1473 ( .A1(n1729), .A2(n1578), .B1(n1730), .B2(n1581), .ZN(n1841)
         );
  XNOR2_X1 U1474 ( .A(a[11]), .B(n1842), .ZN(n830) );
  AOI221_X1 U1475 ( .B1(n1579), .B2(b[22]), .C1(n1553), .C2(n1376), .A(n1843), 
        .ZN(n1842) );
  OAI22_X1 U1476 ( .A1(n1641), .A2(n1582), .B1(n1644), .B2(n1549), .ZN(n1843)
         );
  XNOR2_X1 U1477 ( .A(a[11]), .B(n1844), .ZN(n829) );
  AOI221_X1 U1478 ( .B1(n1580), .B2(b[22]), .C1(n1553), .C2(n1375), .A(n1845), 
        .ZN(n1844) );
  OAI22_X1 U1479 ( .A1(n1617), .A2(n1541), .B1(n1644), .B2(n1581), .ZN(n1845)
         );
  XNOR2_X1 U1480 ( .A(a[11]), .B(n1846), .ZN(n828) );
  AOI221_X1 U1481 ( .B1(n1579), .B2(n1615), .C1(n1580), .C2(n1615), .A(n1847), 
        .ZN(n1846) );
  OAI22_X1 U1482 ( .A1(n1634), .A2(n1578), .B1(n1635), .B2(n1581), .ZN(n1847)
         );
  XNOR2_X1 U1483 ( .A(a[11]), .B(n1848), .ZN(n827) );
  OAI221_X1 U1484 ( .B1(n1618), .B2(n1582), .C1(n1617), .C2(n1578), .A(n1849), 
        .ZN(n1848) );
  OAI21_X1 U1485 ( .B1(n1579), .B2(n1580), .A(n1615), .ZN(n1849) );
  INV_X1 U1486 ( .A(n1853), .ZN(n1850) );
  NAND3_X1 U1487 ( .A1(n1853), .A2(n1852), .A3(n1851), .ZN(n1803) );
  XNOR2_X1 U1488 ( .A(a[10]), .B(a[9]), .ZN(n1851) );
  XNOR2_X1 U1489 ( .A(a[10]), .B(n1607), .ZN(n1852) );
  XOR2_X1 U1490 ( .A(a[9]), .B(n1609), .Z(n1853) );
  XNOR2_X1 U1491 ( .A(n1854), .B(n1605), .ZN(n826) );
  OAI22_X1 U1492 ( .A1(n1565), .A2(n1540), .B1(n1565), .B2(n1583), .ZN(n1854)
         );
  XNOR2_X1 U1493 ( .A(n1855), .B(n1605), .ZN(n825) );
  OAI222_X1 U1494 ( .A1(n1650), .A2(n1540), .B1(n1566), .B2(n1548), .C1(n1651), 
        .C2(n1583), .ZN(n1855) );
  XNOR2_X1 U1495 ( .A(n1604), .B(n1856), .ZN(n824) );
  AOI221_X1 U1496 ( .B1(n1584), .B2(b[2]), .C1(n1585), .C2(b[1]), .A(n1857), 
        .ZN(n1856) );
  OAI22_X1 U1497 ( .A1(n1654), .A2(n1583), .B1(n1565), .B2(n1586), .ZN(n1857)
         );
  XNOR2_X1 U1498 ( .A(n1604), .B(n1859), .ZN(n823) );
  AOI221_X1 U1499 ( .B1(n1584), .B2(b[3]), .C1(n1585), .C2(b[2]), .A(n1860), 
        .ZN(n1859) );
  OAI22_X1 U1500 ( .A1(n1658), .A2(n1583), .B1(n1650), .B2(n1587), .ZN(n1860)
         );
  XNOR2_X1 U1501 ( .A(n1604), .B(n1861), .ZN(n822) );
  AOI221_X1 U1502 ( .B1(n1584), .B2(b[4]), .C1(n1585), .C2(b[3]), .A(n1862), 
        .ZN(n1861) );
  OAI22_X1 U1503 ( .A1(n1661), .A2(n1583), .B1(n1662), .B2(n1587), .ZN(n1862)
         );
  XNOR2_X1 U1504 ( .A(n1604), .B(n1863), .ZN(n821) );
  AOI221_X1 U1505 ( .B1(n1584), .B2(b[5]), .C1(n1585), .C2(b[4]), .A(n1864), 
        .ZN(n1863) );
  OAI22_X1 U1506 ( .A1(n1665), .A2(n1583), .B1(n1666), .B2(n1587), .ZN(n1864)
         );
  XNOR2_X1 U1507 ( .A(n1604), .B(n1865), .ZN(n820) );
  AOI221_X1 U1508 ( .B1(n1584), .B2(b[6]), .C1(n1585), .C2(b[5]), .A(n1866), 
        .ZN(n1865) );
  OAI22_X1 U1509 ( .A1(n1669), .A2(n1583), .B1(n1670), .B2(n1587), .ZN(n1866)
         );
  XNOR2_X1 U1510 ( .A(n1604), .B(n1867), .ZN(n819) );
  AOI221_X1 U1511 ( .B1(n1584), .B2(b[7]), .C1(n1585), .C2(b[6]), .A(n1868), 
        .ZN(n1867) );
  OAI22_X1 U1512 ( .A1(n1673), .A2(n1583), .B1(n1674), .B2(n1587), .ZN(n1868)
         );
  XNOR2_X1 U1513 ( .A(n1604), .B(n1869), .ZN(n818) );
  AOI221_X1 U1514 ( .B1(n1584), .B2(b[8]), .C1(n1585), .C2(b[7]), .A(n1870), 
        .ZN(n1869) );
  OAI22_X1 U1515 ( .A1(n1677), .A2(n1583), .B1(n1678), .B2(n1587), .ZN(n1870)
         );
  XNOR2_X1 U1516 ( .A(n1604), .B(n1871), .ZN(n817) );
  AOI221_X1 U1517 ( .B1(n1584), .B2(b[9]), .C1(n1585), .C2(b[8]), .A(n1872), 
        .ZN(n1871) );
  OAI22_X1 U1518 ( .A1(n1681), .A2(n1583), .B1(n1682), .B2(n1587), .ZN(n1872)
         );
  XNOR2_X1 U1519 ( .A(n1604), .B(n1873), .ZN(n816) );
  AOI221_X1 U1520 ( .B1(n1584), .B2(b[10]), .C1(n1585), .C2(b[9]), .A(n1874), 
        .ZN(n1873) );
  OAI22_X1 U1521 ( .A1(n1685), .A2(n1583), .B1(n1686), .B2(n1587), .ZN(n1874)
         );
  XNOR2_X1 U1522 ( .A(n1604), .B(n1875), .ZN(n815) );
  AOI221_X1 U1523 ( .B1(n1584), .B2(b[11]), .C1(n1585), .C2(b[10]), .A(n1876), 
        .ZN(n1875) );
  OAI22_X1 U1524 ( .A1(n1689), .A2(n1583), .B1(n1690), .B2(n1587), .ZN(n1876)
         );
  XNOR2_X1 U1525 ( .A(n1604), .B(n1877), .ZN(n814) );
  AOI221_X1 U1526 ( .B1(n1584), .B2(b[12]), .C1(n1585), .C2(b[11]), .A(n1878), 
        .ZN(n1877) );
  OAI22_X1 U1527 ( .A1(n1693), .A2(n1583), .B1(n1694), .B2(n1587), .ZN(n1878)
         );
  XNOR2_X1 U1528 ( .A(n1604), .B(n1879), .ZN(n813) );
  AOI221_X1 U1529 ( .B1(n1584), .B2(b[13]), .C1(n1585), .C2(b[12]), .A(n1880), 
        .ZN(n1879) );
  OAI22_X1 U1530 ( .A1(n1697), .A2(n1583), .B1(n1698), .B2(n1586), .ZN(n1880)
         );
  XNOR2_X1 U1531 ( .A(n1604), .B(n1881), .ZN(n812) );
  AOI221_X1 U1532 ( .B1(n1584), .B2(b[14]), .C1(n1585), .C2(b[13]), .A(n1882), 
        .ZN(n1881) );
  OAI22_X1 U1533 ( .A1(n1701), .A2(n1583), .B1(n1702), .B2(n1586), .ZN(n1882)
         );
  XNOR2_X1 U1534 ( .A(n1604), .B(n1883), .ZN(n811) );
  AOI221_X1 U1535 ( .B1(n1584), .B2(b[15]), .C1(n1585), .C2(b[14]), .A(n1884), 
        .ZN(n1883) );
  OAI22_X1 U1536 ( .A1(n1705), .A2(n1583), .B1(n1706), .B2(n1586), .ZN(n1884)
         );
  XNOR2_X1 U1537 ( .A(n1604), .B(n1885), .ZN(n810) );
  AOI221_X1 U1538 ( .B1(n1584), .B2(b[16]), .C1(n1585), .C2(b[15]), .A(n1886), 
        .ZN(n1885) );
  OAI22_X1 U1539 ( .A1(n1709), .A2(n1583), .B1(n1710), .B2(n1586), .ZN(n1886)
         );
  XNOR2_X1 U1540 ( .A(n1604), .B(n1887), .ZN(n809) );
  AOI221_X1 U1541 ( .B1(n1584), .B2(b[17]), .C1(n1585), .C2(b[16]), .A(n1888), 
        .ZN(n1887) );
  OAI22_X1 U1542 ( .A1(n1713), .A2(n1583), .B1(n1714), .B2(n1586), .ZN(n1888)
         );
  XNOR2_X1 U1543 ( .A(n1604), .B(n1889), .ZN(n808) );
  AOI221_X1 U1544 ( .B1(n1584), .B2(b[18]), .C1(n1585), .C2(b[17]), .A(n1890), 
        .ZN(n1889) );
  OAI22_X1 U1545 ( .A1(n1717), .A2(n1583), .B1(n1718), .B2(n1586), .ZN(n1890)
         );
  XNOR2_X1 U1546 ( .A(n1604), .B(n1891), .ZN(n807) );
  AOI221_X1 U1547 ( .B1(n1584), .B2(b[19]), .C1(n1585), .C2(b[18]), .A(n1892), 
        .ZN(n1891) );
  OAI22_X1 U1548 ( .A1(n1721), .A2(n1583), .B1(n1722), .B2(n1586), .ZN(n1892)
         );
  XNOR2_X1 U1549 ( .A(n1604), .B(n1893), .ZN(n806) );
  AOI221_X1 U1550 ( .B1(n1584), .B2(b[20]), .C1(n1585), .C2(b[19]), .A(n1894), 
        .ZN(n1893) );
  OAI22_X1 U1551 ( .A1(n1725), .A2(n1583), .B1(n1726), .B2(n1586), .ZN(n1894)
         );
  XNOR2_X1 U1552 ( .A(a[14]), .B(n1895), .ZN(n805) );
  AOI221_X1 U1553 ( .B1(n1584), .B2(b[21]), .C1(n1585), .C2(b[20]), .A(n1896), 
        .ZN(n1895) );
  OAI22_X1 U1554 ( .A1(n1729), .A2(n1583), .B1(n1730), .B2(n1586), .ZN(n1896)
         );
  XNOR2_X1 U1555 ( .A(a[14]), .B(n1897), .ZN(n804) );
  AOI221_X1 U1556 ( .B1(n1584), .B2(b[22]), .C1(n1552), .C2(n1376), .A(n1898), 
        .ZN(n1897) );
  OAI22_X1 U1557 ( .A1(n1641), .A2(n1587), .B1(n1644), .B2(n1548), .ZN(n1898)
         );
  XNOR2_X1 U1558 ( .A(a[14]), .B(n1899), .ZN(n803) );
  AOI221_X1 U1559 ( .B1(n1585), .B2(b[22]), .C1(n1552), .C2(n1375), .A(n1900), 
        .ZN(n1899) );
  OAI22_X1 U1560 ( .A1(n1617), .A2(n1540), .B1(n1644), .B2(n1586), .ZN(n1900)
         );
  XNOR2_X1 U1561 ( .A(a[14]), .B(n1901), .ZN(n802) );
  AOI221_X1 U1562 ( .B1(n1584), .B2(n1615), .C1(n1585), .C2(n1615), .A(n1902), 
        .ZN(n1901) );
  OAI22_X1 U1563 ( .A1(n1634), .A2(n1583), .B1(n1635), .B2(n1586), .ZN(n1902)
         );
  XNOR2_X1 U1564 ( .A(a[14]), .B(n1903), .ZN(n801) );
  OAI221_X1 U1565 ( .B1(n1617), .B2(n1587), .C1(n1620), .C2(n1583), .A(n1904), 
        .ZN(n1903) );
  OAI21_X1 U1566 ( .B1(n1584), .B2(n1585), .A(n1615), .ZN(n1904) );
  INV_X1 U1567 ( .A(n1908), .ZN(n1905) );
  NAND3_X1 U1568 ( .A1(n1908), .A2(n1907), .A3(n1906), .ZN(n1858) );
  XNOR2_X1 U1569 ( .A(a[12]), .B(a[13]), .ZN(n1906) );
  XNOR2_X1 U1570 ( .A(a[13]), .B(n1605), .ZN(n1907) );
  XOR2_X1 U1571 ( .A(a[12]), .B(n1607), .Z(n1908) );
  XNOR2_X1 U1572 ( .A(n1909), .B(n1603), .ZN(n800) );
  OAI22_X1 U1573 ( .A1(n1565), .A2(n1539), .B1(n1566), .B2(n1588), .ZN(n1909)
         );
  XNOR2_X1 U1574 ( .A(n1910), .B(n1603), .ZN(n799) );
  OAI222_X1 U1575 ( .A1(n1650), .A2(n1539), .B1(n1566), .B2(n1547), .C1(n1651), 
        .C2(n1588), .ZN(n1910) );
  XNOR2_X1 U1576 ( .A(n1602), .B(n1911), .ZN(n798) );
  AOI221_X1 U1577 ( .B1(n1589), .B2(b[2]), .C1(n1590), .C2(b[1]), .A(n1912), 
        .ZN(n1911) );
  OAI22_X1 U1578 ( .A1(n1654), .A2(n1588), .B1(n1566), .B2(n1591), .ZN(n1912)
         );
  XNOR2_X1 U1579 ( .A(n1602), .B(n1914), .ZN(n797) );
  AOI221_X1 U1580 ( .B1(n1589), .B2(b[3]), .C1(n1590), .C2(b[2]), .A(n1915), 
        .ZN(n1914) );
  OAI22_X1 U1581 ( .A1(n1658), .A2(n1588), .B1(n1650), .B2(n1592), .ZN(n1915)
         );
  XNOR2_X1 U1582 ( .A(n1602), .B(n1916), .ZN(n796) );
  AOI221_X1 U1583 ( .B1(n1589), .B2(b[4]), .C1(n1590), .C2(b[3]), .A(n1917), 
        .ZN(n1916) );
  OAI22_X1 U1584 ( .A1(n1661), .A2(n1588), .B1(n1662), .B2(n1592), .ZN(n1917)
         );
  XNOR2_X1 U1585 ( .A(n1602), .B(n1918), .ZN(n795) );
  AOI221_X1 U1586 ( .B1(n1589), .B2(b[5]), .C1(n1590), .C2(b[4]), .A(n1919), 
        .ZN(n1918) );
  OAI22_X1 U1587 ( .A1(n1665), .A2(n1588), .B1(n1666), .B2(n1592), .ZN(n1919)
         );
  XNOR2_X1 U1588 ( .A(n1602), .B(n1920), .ZN(n794) );
  AOI221_X1 U1589 ( .B1(n1589), .B2(b[6]), .C1(n1590), .C2(b[5]), .A(n1921), 
        .ZN(n1920) );
  OAI22_X1 U1590 ( .A1(n1669), .A2(n1588), .B1(n1670), .B2(n1592), .ZN(n1921)
         );
  XNOR2_X1 U1591 ( .A(n1602), .B(n1922), .ZN(n793) );
  AOI221_X1 U1592 ( .B1(n1589), .B2(b[7]), .C1(n1590), .C2(b[6]), .A(n1923), 
        .ZN(n1922) );
  OAI22_X1 U1593 ( .A1(n1673), .A2(n1588), .B1(n1674), .B2(n1592), .ZN(n1923)
         );
  XNOR2_X1 U1594 ( .A(n1602), .B(n1924), .ZN(n792) );
  AOI221_X1 U1595 ( .B1(n1589), .B2(b[8]), .C1(n1590), .C2(b[7]), .A(n1925), 
        .ZN(n1924) );
  OAI22_X1 U1596 ( .A1(n1677), .A2(n1588), .B1(n1678), .B2(n1592), .ZN(n1925)
         );
  XNOR2_X1 U1597 ( .A(n1602), .B(n1926), .ZN(n791) );
  AOI221_X1 U1598 ( .B1(n1589), .B2(b[9]), .C1(n1590), .C2(b[8]), .A(n1927), 
        .ZN(n1926) );
  OAI22_X1 U1599 ( .A1(n1681), .A2(n1588), .B1(n1682), .B2(n1592), .ZN(n1927)
         );
  XNOR2_X1 U1600 ( .A(n1602), .B(n1928), .ZN(n790) );
  AOI221_X1 U1601 ( .B1(n1589), .B2(b[10]), .C1(n1590), .C2(b[9]), .A(n1929), 
        .ZN(n1928) );
  OAI22_X1 U1602 ( .A1(n1685), .A2(n1588), .B1(n1686), .B2(n1592), .ZN(n1929)
         );
  XNOR2_X1 U1603 ( .A(n1602), .B(n1930), .ZN(n789) );
  AOI221_X1 U1604 ( .B1(n1589), .B2(b[11]), .C1(n1590), .C2(b[10]), .A(n1931), 
        .ZN(n1930) );
  OAI22_X1 U1605 ( .A1(n1689), .A2(n1588), .B1(n1690), .B2(n1592), .ZN(n1931)
         );
  XNOR2_X1 U1606 ( .A(n1602), .B(n1932), .ZN(n788) );
  AOI221_X1 U1607 ( .B1(n1589), .B2(b[12]), .C1(n1590), .C2(b[11]), .A(n1933), 
        .ZN(n1932) );
  OAI22_X1 U1608 ( .A1(n1693), .A2(n1588), .B1(n1694), .B2(n1592), .ZN(n1933)
         );
  XNOR2_X1 U1609 ( .A(n1602), .B(n1934), .ZN(n787) );
  AOI221_X1 U1610 ( .B1(n1589), .B2(b[13]), .C1(n1590), .C2(b[12]), .A(n1935), 
        .ZN(n1934) );
  OAI22_X1 U1611 ( .A1(n1697), .A2(n1588), .B1(n1698), .B2(n1591), .ZN(n1935)
         );
  XNOR2_X1 U1612 ( .A(n1602), .B(n1936), .ZN(n786) );
  AOI221_X1 U1613 ( .B1(n1589), .B2(b[14]), .C1(n1590), .C2(b[13]), .A(n1937), 
        .ZN(n1936) );
  OAI22_X1 U1614 ( .A1(n1701), .A2(n1588), .B1(n1702), .B2(n1591), .ZN(n1937)
         );
  XNOR2_X1 U1615 ( .A(n1602), .B(n1938), .ZN(n785) );
  AOI221_X1 U1616 ( .B1(n1589), .B2(b[15]), .C1(n1590), .C2(b[14]), .A(n1939), 
        .ZN(n1938) );
  OAI22_X1 U1617 ( .A1(n1705), .A2(n1588), .B1(n1706), .B2(n1591), .ZN(n1939)
         );
  XNOR2_X1 U1618 ( .A(n1602), .B(n1940), .ZN(n784) );
  AOI221_X1 U1619 ( .B1(n1589), .B2(b[16]), .C1(n1590), .C2(b[15]), .A(n1941), 
        .ZN(n1940) );
  OAI22_X1 U1620 ( .A1(n1709), .A2(n1588), .B1(n1710), .B2(n1591), .ZN(n1941)
         );
  XNOR2_X1 U1621 ( .A(n1602), .B(n1942), .ZN(n783) );
  AOI221_X1 U1622 ( .B1(n1589), .B2(b[17]), .C1(n1590), .C2(b[16]), .A(n1943), 
        .ZN(n1942) );
  OAI22_X1 U1623 ( .A1(n1713), .A2(n1588), .B1(n1714), .B2(n1591), .ZN(n1943)
         );
  XNOR2_X1 U1624 ( .A(n1602), .B(n1944), .ZN(n782) );
  AOI221_X1 U1625 ( .B1(n1589), .B2(b[18]), .C1(n1590), .C2(b[17]), .A(n1945), 
        .ZN(n1944) );
  OAI22_X1 U1626 ( .A1(n1717), .A2(n1588), .B1(n1718), .B2(n1591), .ZN(n1945)
         );
  XNOR2_X1 U1627 ( .A(n1602), .B(n1946), .ZN(n781) );
  AOI221_X1 U1628 ( .B1(n1589), .B2(b[19]), .C1(n1590), .C2(b[18]), .A(n1947), 
        .ZN(n1946) );
  OAI22_X1 U1629 ( .A1(n1721), .A2(n1588), .B1(n1722), .B2(n1591), .ZN(n1947)
         );
  XNOR2_X1 U1630 ( .A(n1602), .B(n1948), .ZN(n780) );
  AOI221_X1 U1631 ( .B1(n1589), .B2(b[20]), .C1(n1590), .C2(b[19]), .A(n1949), 
        .ZN(n1948) );
  OAI22_X1 U1632 ( .A1(n1725), .A2(n1588), .B1(n1726), .B2(n1591), .ZN(n1949)
         );
  XNOR2_X1 U1633 ( .A(a[17]), .B(n1950), .ZN(n779) );
  AOI221_X1 U1634 ( .B1(n1589), .B2(b[21]), .C1(n1590), .C2(b[20]), .A(n1951), 
        .ZN(n1950) );
  OAI22_X1 U1635 ( .A1(n1729), .A2(n1588), .B1(n1730), .B2(n1591), .ZN(n1951)
         );
  XNOR2_X1 U1636 ( .A(a[17]), .B(n1952), .ZN(n778) );
  AOI221_X1 U1637 ( .B1(n1589), .B2(b[22]), .C1(n1551), .C2(n1376), .A(n1953), 
        .ZN(n1952) );
  OAI22_X1 U1638 ( .A1(n1641), .A2(n1592), .B1(n1644), .B2(n1547), .ZN(n1953)
         );
  XNOR2_X1 U1639 ( .A(a[17]), .B(n1954), .ZN(n777) );
  AOI221_X1 U1640 ( .B1(n1590), .B2(b[22]), .C1(n1551), .C2(n1375), .A(n1955), 
        .ZN(n1954) );
  OAI22_X1 U1641 ( .A1(n1617), .A2(n1539), .B1(n1644), .B2(n1591), .ZN(n1955)
         );
  XNOR2_X1 U1642 ( .A(a[17]), .B(n1956), .ZN(n776) );
  AOI221_X1 U1643 ( .B1(n1589), .B2(n1614), .C1(n1590), .C2(n1615), .A(n1957), 
        .ZN(n1956) );
  OAI22_X1 U1644 ( .A1(n1634), .A2(n1588), .B1(n1635), .B2(n1591), .ZN(n1957)
         );
  XNOR2_X1 U1645 ( .A(a[17]), .B(n1958), .ZN(n775) );
  OAI221_X1 U1646 ( .B1(n1619), .B2(n1592), .C1(n1617), .C2(n1588), .A(n1959), 
        .ZN(n1958) );
  OAI21_X1 U1647 ( .B1(n1589), .B2(n1590), .A(n1615), .ZN(n1959) );
  INV_X1 U1648 ( .A(n1963), .ZN(n1960) );
  NAND3_X1 U1649 ( .A1(n1963), .A2(n1962), .A3(n1961), .ZN(n1913) );
  XNOR2_X1 U1650 ( .A(a[15]), .B(a[16]), .ZN(n1961) );
  XNOR2_X1 U1651 ( .A(a[16]), .B(n1603), .ZN(n1962) );
  XOR2_X1 U1652 ( .A(a[15]), .B(n1605), .Z(n1963) );
  XOR2_X1 U1653 ( .A(n1964), .B(n1600), .Z(n774) );
  OAI22_X1 U1654 ( .A1(n1565), .A2(n1538), .B1(n1566), .B2(n1593), .ZN(n1964)
         );
  XOR2_X1 U1655 ( .A(n1965), .B(n1600), .Z(n773) );
  OAI222_X1 U1656 ( .A1(n1650), .A2(n1538), .B1(n1566), .B2(n1546), .C1(n1651), 
        .C2(n1593), .ZN(n1965) );
  XNOR2_X1 U1657 ( .A(n1600), .B(n1966), .ZN(n772) );
  AOI221_X1 U1658 ( .B1(n1594), .B2(b[2]), .C1(n1595), .C2(b[1]), .A(n1967), 
        .ZN(n1966) );
  OAI22_X1 U1659 ( .A1(n1654), .A2(n1593), .B1(n1566), .B2(n1596), .ZN(n1967)
         );
  XNOR2_X1 U1660 ( .A(n1600), .B(n1969), .ZN(n771) );
  AOI221_X1 U1661 ( .B1(n1594), .B2(b[3]), .C1(n1595), .C2(b[2]), .A(n1970), 
        .ZN(n1969) );
  OAI22_X1 U1662 ( .A1(n1658), .A2(n1593), .B1(n1650), .B2(n1597), .ZN(n1970)
         );
  XNOR2_X1 U1663 ( .A(n1600), .B(n1971), .ZN(n770) );
  AOI221_X1 U1664 ( .B1(n1594), .B2(b[4]), .C1(n1595), .C2(b[3]), .A(n1972), 
        .ZN(n1971) );
  OAI22_X1 U1665 ( .A1(n1661), .A2(n1593), .B1(n1662), .B2(n1597), .ZN(n1972)
         );
  XNOR2_X1 U1666 ( .A(n1600), .B(n1973), .ZN(n769) );
  AOI221_X1 U1667 ( .B1(n1594), .B2(b[5]), .C1(n1595), .C2(b[4]), .A(n1974), 
        .ZN(n1973) );
  OAI22_X1 U1668 ( .A1(n1665), .A2(n1593), .B1(n1666), .B2(n1597), .ZN(n1974)
         );
  XNOR2_X1 U1669 ( .A(n1600), .B(n1975), .ZN(n768) );
  AOI221_X1 U1670 ( .B1(n1594), .B2(b[6]), .C1(n1595), .C2(b[5]), .A(n1976), 
        .ZN(n1975) );
  OAI22_X1 U1671 ( .A1(n1669), .A2(n1593), .B1(n1670), .B2(n1597), .ZN(n1976)
         );
  XNOR2_X1 U1672 ( .A(n1600), .B(n1977), .ZN(n767) );
  AOI221_X1 U1673 ( .B1(n1594), .B2(b[7]), .C1(n1595), .C2(b[6]), .A(n1978), 
        .ZN(n1977) );
  OAI22_X1 U1674 ( .A1(n1673), .A2(n1593), .B1(n1674), .B2(n1597), .ZN(n1978)
         );
  XNOR2_X1 U1675 ( .A(n1600), .B(n1979), .ZN(n766) );
  AOI221_X1 U1676 ( .B1(n1594), .B2(b[8]), .C1(n1595), .C2(b[7]), .A(n1980), 
        .ZN(n1979) );
  OAI22_X1 U1677 ( .A1(n1677), .A2(n1593), .B1(n1678), .B2(n1597), .ZN(n1980)
         );
  XNOR2_X1 U1678 ( .A(n1600), .B(n1981), .ZN(n765) );
  AOI221_X1 U1679 ( .B1(n1594), .B2(b[9]), .C1(n1595), .C2(b[8]), .A(n1982), 
        .ZN(n1981) );
  OAI22_X1 U1680 ( .A1(n1681), .A2(n1593), .B1(n1682), .B2(n1597), .ZN(n1982)
         );
  XNOR2_X1 U1681 ( .A(n1600), .B(n1983), .ZN(n764) );
  AOI221_X1 U1682 ( .B1(n1594), .B2(b[10]), .C1(n1595), .C2(b[9]), .A(n1984), 
        .ZN(n1983) );
  OAI22_X1 U1683 ( .A1(n1685), .A2(n1593), .B1(n1686), .B2(n1597), .ZN(n1984)
         );
  XNOR2_X1 U1684 ( .A(n1600), .B(n1985), .ZN(n763) );
  AOI221_X1 U1685 ( .B1(n1594), .B2(b[11]), .C1(n1595), .C2(b[10]), .A(n1986), 
        .ZN(n1985) );
  OAI22_X1 U1686 ( .A1(n1689), .A2(n1593), .B1(n1690), .B2(n1597), .ZN(n1986)
         );
  XNOR2_X1 U1687 ( .A(n1601), .B(n1987), .ZN(n762) );
  AOI221_X1 U1688 ( .B1(n1594), .B2(b[12]), .C1(n1595), .C2(b[11]), .A(n1988), 
        .ZN(n1987) );
  OAI22_X1 U1689 ( .A1(n1693), .A2(n1593), .B1(n1694), .B2(n1597), .ZN(n1988)
         );
  XNOR2_X1 U1690 ( .A(n1601), .B(n1989), .ZN(n761) );
  AOI221_X1 U1691 ( .B1(n1594), .B2(b[13]), .C1(n1595), .C2(b[12]), .A(n1990), 
        .ZN(n1989) );
  OAI22_X1 U1692 ( .A1(n1697), .A2(n1593), .B1(n1698), .B2(n1596), .ZN(n1990)
         );
  XNOR2_X1 U1693 ( .A(n1601), .B(n1991), .ZN(n760) );
  AOI221_X1 U1694 ( .B1(n1594), .B2(b[14]), .C1(n1595), .C2(b[13]), .A(n1992), 
        .ZN(n1991) );
  OAI22_X1 U1695 ( .A1(n1701), .A2(n1593), .B1(n1702), .B2(n1596), .ZN(n1992)
         );
  XNOR2_X1 U1696 ( .A(n1601), .B(n1993), .ZN(n759) );
  AOI221_X1 U1697 ( .B1(n1594), .B2(b[15]), .C1(n1595), .C2(b[14]), .A(n1994), 
        .ZN(n1993) );
  OAI22_X1 U1698 ( .A1(n1705), .A2(n1593), .B1(n1706), .B2(n1596), .ZN(n1994)
         );
  XNOR2_X1 U1699 ( .A(n1601), .B(n1995), .ZN(n758) );
  AOI221_X1 U1700 ( .B1(n1594), .B2(b[16]), .C1(n1595), .C2(b[15]), .A(n1996), 
        .ZN(n1995) );
  OAI22_X1 U1701 ( .A1(n1709), .A2(n1593), .B1(n1710), .B2(n1596), .ZN(n1996)
         );
  XNOR2_X1 U1702 ( .A(n1601), .B(n1997), .ZN(n757) );
  AOI221_X1 U1703 ( .B1(n1594), .B2(b[17]), .C1(n1595), .C2(b[16]), .A(n1998), 
        .ZN(n1997) );
  OAI22_X1 U1704 ( .A1(n1713), .A2(n1593), .B1(n1714), .B2(n1596), .ZN(n1998)
         );
  XNOR2_X1 U1705 ( .A(n1601), .B(n1999), .ZN(n756) );
  AOI221_X1 U1706 ( .B1(n1594), .B2(b[18]), .C1(n1595), .C2(b[17]), .A(n2000), 
        .ZN(n1999) );
  OAI22_X1 U1707 ( .A1(n1717), .A2(n1593), .B1(n1718), .B2(n1596), .ZN(n2000)
         );
  XNOR2_X1 U1708 ( .A(n1601), .B(n2001), .ZN(n755) );
  AOI221_X1 U1709 ( .B1(n1594), .B2(b[19]), .C1(n1595), .C2(b[18]), .A(n2002), 
        .ZN(n2001) );
  OAI22_X1 U1710 ( .A1(n1721), .A2(n1593), .B1(n1722), .B2(n1596), .ZN(n2002)
         );
  XNOR2_X1 U1711 ( .A(n1601), .B(n2003), .ZN(n754) );
  AOI221_X1 U1712 ( .B1(n1594), .B2(b[20]), .C1(n1595), .C2(b[19]), .A(n2004), 
        .ZN(n2003) );
  OAI22_X1 U1713 ( .A1(n1725), .A2(n1593), .B1(n1726), .B2(n1596), .ZN(n2004)
         );
  XNOR2_X1 U1714 ( .A(n1601), .B(n2005), .ZN(n753) );
  AOI221_X1 U1715 ( .B1(n1594), .B2(b[21]), .C1(n1595), .C2(b[20]), .A(n2006), 
        .ZN(n2005) );
  OAI22_X1 U1716 ( .A1(n1729), .A2(n1593), .B1(n1730), .B2(n1596), .ZN(n2006)
         );
  XNOR2_X1 U1717 ( .A(n1601), .B(n2007), .ZN(n752) );
  AOI221_X1 U1718 ( .B1(n1594), .B2(b[22]), .C1(n1544), .C2(n1376), .A(n2008), 
        .ZN(n2007) );
  OAI22_X1 U1719 ( .A1(n1641), .A2(n1597), .B1(n1644), .B2(n1546), .ZN(n2008)
         );
  XNOR2_X1 U1720 ( .A(n1601), .B(n2009), .ZN(n751) );
  AOI221_X1 U1721 ( .B1(n1595), .B2(b[22]), .C1(n1544), .C2(n1375), .A(n2010), 
        .ZN(n2009) );
  OAI22_X1 U1722 ( .A1(n1617), .A2(n1538), .B1(n1644), .B2(n1596), .ZN(n2010)
         );
  XNOR2_X1 U1723 ( .A(n1601), .B(n2011), .ZN(n750) );
  AOI221_X1 U1724 ( .B1(n1594), .B2(n1613), .C1(n1595), .C2(n1615), .A(n2012), 
        .ZN(n2011) );
  OAI22_X1 U1725 ( .A1(n1634), .A2(n1593), .B1(n1635), .B2(n1596), .ZN(n2012)
         );
  INV_X1 U1726 ( .A(b[22]), .ZN(n1635) );
  INV_X1 U1727 ( .A(n1374), .ZN(n1634) );
  XNOR2_X1 U1728 ( .A(n1600), .B(n2013), .ZN(n749) );
  OAI221_X1 U1729 ( .B1(n1617), .B2(n1597), .C1(n1620), .C2(n1593), .A(n2014), 
        .ZN(n2013) );
  OAI21_X1 U1730 ( .B1(n1594), .B2(n1595), .A(n1615), .ZN(n2014) );
  INV_X1 U1731 ( .A(n2018), .ZN(n2015) );
  NAND3_X1 U1732 ( .A1(n2018), .A2(n2017), .A3(n2016), .ZN(n1968) );
  XNOR2_X1 U1733 ( .A(a[18]), .B(a[19]), .ZN(n2016) );
  XOR2_X1 U1734 ( .A(a[19]), .B(n1600), .Z(n2017) );
  XOR2_X1 U1735 ( .A(a[18]), .B(n1603), .Z(n2018) );
  XNOR2_X1 U1736 ( .A(n2019), .B(n1599), .ZN(n748) );
  OAI22_X1 U1737 ( .A1(n1537), .A2(n1567), .B1(n1558), .B2(n1567), .ZN(n2019)
         );
  XNOR2_X1 U1738 ( .A(n2020), .B(n1599), .ZN(n747) );
  OAI222_X1 U1739 ( .A1(n1537), .A2(n1650), .B1(n1545), .B2(n1566), .C1(n1558), 
        .C2(n1651), .ZN(n2020) );
  XNOR2_X1 U1740 ( .A(n1598), .B(n2021), .ZN(n746) );
  AOI221_X1 U1741 ( .B1(b[2]), .B2(n1559), .C1(b[1]), .C2(n1560), .A(n2022), 
        .ZN(n2021) );
  OAI22_X1 U1742 ( .A1(n1558), .A2(n1654), .B1(n1557), .B2(n1567), .ZN(n2022)
         );
  INV_X1 U1743 ( .A(b[0]), .ZN(n1648) );
  INV_X1 U1744 ( .A(n1396), .ZN(n1654) );
  XNOR2_X1 U1745 ( .A(n1598), .B(n2023), .ZN(n745) );
  AOI221_X1 U1746 ( .B1(b[3]), .B2(n1559), .C1(b[2]), .C2(n1560), .A(n2024), 
        .ZN(n2023) );
  OAI22_X1 U1747 ( .A1(n1558), .A2(n1658), .B1(n1557), .B2(n1650), .ZN(n2024)
         );
  XNOR2_X1 U1748 ( .A(n1598), .B(n2025), .ZN(n744) );
  AOI221_X1 U1749 ( .B1(b[4]), .B2(n1559), .C1(b[3]), .C2(n1560), .A(n2026), 
        .ZN(n2025) );
  OAI22_X1 U1750 ( .A1(n1558), .A2(n1661), .B1(n1557), .B2(n1662), .ZN(n2026)
         );
  XNOR2_X1 U1751 ( .A(n1598), .B(n2027), .ZN(n743) );
  AOI221_X1 U1752 ( .B1(b[5]), .B2(n1559), .C1(b[4]), .C2(n1560), .A(n2028), 
        .ZN(n2027) );
  OAI22_X1 U1753 ( .A1(n1558), .A2(n1665), .B1(n1557), .B2(n1666), .ZN(n2028)
         );
  XNOR2_X1 U1754 ( .A(n1598), .B(n2029), .ZN(n742) );
  AOI221_X1 U1755 ( .B1(b[6]), .B2(n1559), .C1(b[5]), .C2(n1560), .A(n2030), 
        .ZN(n2029) );
  OAI22_X1 U1756 ( .A1(n1558), .A2(n1669), .B1(n1557), .B2(n1670), .ZN(n2030)
         );
  XNOR2_X1 U1757 ( .A(n1598), .B(n2031), .ZN(n741) );
  AOI221_X1 U1758 ( .B1(b[7]), .B2(n1559), .C1(b[6]), .C2(n1560), .A(n2032), 
        .ZN(n2031) );
  OAI22_X1 U1759 ( .A1(n1558), .A2(n1673), .B1(n1557), .B2(n1674), .ZN(n2032)
         );
  XNOR2_X1 U1760 ( .A(n1598), .B(n2033), .ZN(n740) );
  AOI221_X1 U1761 ( .B1(b[9]), .B2(n1559), .C1(b[8]), .C2(n1560), .A(n2034), 
        .ZN(n2033) );
  OAI22_X1 U1762 ( .A1(n1558), .A2(n1681), .B1(n1557), .B2(n1682), .ZN(n2034)
         );
  XNOR2_X1 U1763 ( .A(n1598), .B(n2035), .ZN(n739) );
  AOI221_X1 U1764 ( .B1(b[10]), .B2(n1559), .C1(b[9]), .C2(n1560), .A(n2036), 
        .ZN(n2035) );
  OAI22_X1 U1765 ( .A1(n1558), .A2(n1685), .B1(n1557), .B2(n1686), .ZN(n2036)
         );
  XNOR2_X1 U1766 ( .A(n1598), .B(n2037), .ZN(n738) );
  AOI221_X1 U1767 ( .B1(b[12]), .B2(n1559), .C1(b[11]), .C2(n1560), .A(n2038), 
        .ZN(n2037) );
  OAI22_X1 U1768 ( .A1(n1558), .A2(n1693), .B1(n1557), .B2(n1694), .ZN(n2038)
         );
  XNOR2_X1 U1769 ( .A(n1598), .B(n2039), .ZN(n737) );
  AOI221_X1 U1770 ( .B1(b[13]), .B2(n1559), .C1(b[12]), .C2(n1560), .A(n2040), 
        .ZN(n2039) );
  OAI22_X1 U1771 ( .A1(n1558), .A2(n1697), .B1(n1557), .B2(n1698), .ZN(n2040)
         );
  XNOR2_X1 U1772 ( .A(n1598), .B(n2041), .ZN(n736) );
  AOI221_X1 U1773 ( .B1(b[14]), .B2(n1559), .C1(b[13]), .C2(n1560), .A(n2042), 
        .ZN(n2041) );
  OAI22_X1 U1774 ( .A1(n1558), .A2(n1701), .B1(n1556), .B2(n1702), .ZN(n2042)
         );
  XNOR2_X1 U1775 ( .A(n1598), .B(n2043), .ZN(n735) );
  AOI221_X1 U1776 ( .B1(b[15]), .B2(n1559), .C1(b[14]), .C2(n1560), .A(n2044), 
        .ZN(n2043) );
  OAI22_X1 U1777 ( .A1(n1558), .A2(n1705), .B1(n1556), .B2(n1706), .ZN(n2044)
         );
  XNOR2_X1 U1778 ( .A(n1598), .B(n2045), .ZN(n734) );
  AOI221_X1 U1779 ( .B1(b[16]), .B2(n1559), .C1(b[15]), .C2(n1560), .A(n2046), 
        .ZN(n2045) );
  OAI22_X1 U1780 ( .A1(n1558), .A2(n1709), .B1(n1556), .B2(n1710), .ZN(n2046)
         );
  XNOR2_X1 U1781 ( .A(n1598), .B(n2047), .ZN(n733) );
  AOI221_X1 U1782 ( .B1(b[18]), .B2(n1559), .C1(b[17]), .C2(n1560), .A(n2048), 
        .ZN(n2047) );
  OAI22_X1 U1783 ( .A1(n1558), .A2(n1717), .B1(n1556), .B2(n1718), .ZN(n2048)
         );
  XNOR2_X1 U1784 ( .A(n1598), .B(n2049), .ZN(n732) );
  AOI221_X1 U1785 ( .B1(b[19]), .B2(n1559), .C1(b[18]), .C2(n1560), .A(n2050), 
        .ZN(n2049) );
  OAI22_X1 U1786 ( .A1(n1558), .A2(n1721), .B1(n1556), .B2(n1722), .ZN(n2050)
         );
  XNOR2_X1 U1787 ( .A(n1598), .B(n2051), .ZN(n731) );
  AOI221_X1 U1788 ( .B1(b[20]), .B2(n1559), .C1(b[19]), .C2(n1560), .A(n2052), 
        .ZN(n2051) );
  OAI22_X1 U1789 ( .A1(n1558), .A2(n1725), .B1(n1556), .B2(n1726), .ZN(n2052)
         );
  XNOR2_X1 U1790 ( .A(a[23]), .B(n2053), .ZN(n730) );
  AOI221_X1 U1791 ( .B1(b[21]), .B2(n1559), .C1(b[20]), .C2(n1560), .A(n2054), 
        .ZN(n2053) );
  OAI22_X1 U1792 ( .A1(n1558), .A2(n1729), .B1(n1556), .B2(n1730), .ZN(n2054)
         );
  XNOR2_X1 U1793 ( .A(a[23]), .B(n2055), .ZN(n729) );
  AOI221_X1 U1794 ( .B1(b[22]), .B2(n1559), .C1(n1376), .C2(n1543), .A(n2056), 
        .ZN(n2055) );
  OAI22_X1 U1795 ( .A1(n1556), .A2(n1641), .B1(n1545), .B2(n1644), .ZN(n2056)
         );
  INV_X1 U1796 ( .A(b[20]), .ZN(n1641) );
  XNOR2_X1 U1797 ( .A(n519), .B(n2057), .ZN(n506) );
  INV_X1 U1798 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1799 ( .A1(n2057), .A2(n519), .ZN(n493) );
  XOR2_X1 U1800 ( .A(n2058), .B(n1743), .Z(n2057) );
  OAI221_X1 U1801 ( .B1(n1619), .B2(n1640), .C1(n1620), .C2(n1564), .A(n2059), 
        .ZN(n2058) );
  OAI21_X1 U1802 ( .B1(n1561), .B2(n1563), .A(n1615), .ZN(n2059) );
  INV_X1 U1803 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1804 ( .A(n1598), .B(n2060), .Z(n454) );
  AOI221_X1 U1805 ( .B1(b[8]), .B2(n1559), .C1(b[7]), .C2(n1560), .A(n2061), 
        .ZN(n2060) );
  OAI22_X1 U1806 ( .A1(n1558), .A2(n1677), .B1(n1556), .B2(n1678), .ZN(n2061)
         );
  INV_X1 U1807 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1808 ( .A(n1598), .B(n2062), .Z(n421) );
  AOI221_X1 U1809 ( .B1(b[11]), .B2(n1559), .C1(b[10]), .C2(n1560), .A(n2063), 
        .ZN(n2062) );
  OAI22_X1 U1810 ( .A1(n1558), .A2(n1689), .B1(n1556), .B2(n1690), .ZN(n2063)
         );
  INV_X1 U1811 ( .A(n387), .ZN(n395) );
  INV_X1 U1812 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1813 ( .A(n1598), .B(n2064), .Z(n374) );
  AOI221_X1 U1814 ( .B1(b[17]), .B2(n1559), .C1(b[16]), .C2(n1560), .A(n2065), 
        .ZN(n2064) );
  OAI22_X1 U1815 ( .A1(n1558), .A2(n1713), .B1(n1556), .B2(n1714), .ZN(n2065)
         );
  INV_X1 U1816 ( .A(n356), .ZN(n360) );
  INV_X1 U1817 ( .A(n1628), .ZN(n351) );
  XOR2_X1 U1818 ( .A(n1599), .B(n2066), .Z(n1628) );
  AOI221_X1 U1819 ( .B1(b[22]), .B2(n1560), .C1(n1375), .C2(n1543), .A(n2067), 
        .ZN(n2066) );
  OAI22_X1 U1820 ( .A1(n1537), .A2(n1619), .B1(n1556), .B2(n1644), .ZN(n2067)
         );
  INV_X1 U1821 ( .A(b[21]), .ZN(n1644) );
  NAND3_X1 U1822 ( .A1(n2068), .A2(n2069), .A3(n2070), .ZN(n1630) );
  XNOR2_X1 U1823 ( .A(a[22]), .B(n1599), .ZN(n2069) );
  XNOR2_X1 U1824 ( .A(a[21]), .B(a[22]), .ZN(n2070) );
  INV_X1 U1825 ( .A(n2068), .ZN(n2071) );
  XNOR2_X1 U1826 ( .A(a[21]), .B(n1600), .ZN(n2068) );
  OAI222_X1 U1827 ( .A1(n2072), .A2(n2073), .B1(n2072), .B2(n2074), .C1(n2074), 
        .C2(n2073), .ZN(n326) );
  INV_X1 U1828 ( .A(n550), .ZN(n2074) );
  XNOR2_X1 U1829 ( .A(n1743), .B(n2075), .ZN(n2073) );
  AOI221_X1 U1830 ( .B1(n1561), .B2(b[21]), .C1(b[20]), .C2(n1562), .A(n2076), 
        .ZN(n2075) );
  OAI22_X1 U1831 ( .A1(n1564), .A2(n1729), .B1(n1640), .B2(n1730), .ZN(n2076)
         );
  INV_X1 U1832 ( .A(b[19]), .ZN(n1730) );
  INV_X1 U1833 ( .A(n1377), .ZN(n1729) );
  AOI222_X1 U1834 ( .A1(n2077), .A2(n2078), .B1(n2077), .B2(n564), .C1(n564), 
        .C2(n2078), .ZN(n2072) );
  XNOR2_X1 U1835 ( .A(a[2]), .B(n2079), .ZN(n2078) );
  AOI221_X1 U1836 ( .B1(b[20]), .B2(n1561), .C1(b[19]), .C2(n1562), .A(n2080), 
        .ZN(n2079) );
  OAI22_X1 U1837 ( .A1(n1564), .A2(n1725), .B1(n1640), .B2(n1726), .ZN(n2080)
         );
  INV_X1 U1838 ( .A(b[18]), .ZN(n1726) );
  INV_X1 U1839 ( .A(n1378), .ZN(n1725) );
  INV_X1 U1840 ( .A(n2081), .ZN(n2077) );
  AOI222_X1 U1841 ( .A1(n2082), .A2(n2083), .B1(n2082), .B2(n576), .C1(n576), 
        .C2(n2083), .ZN(n2081) );
  XNOR2_X1 U1842 ( .A(a[2]), .B(n2084), .ZN(n2083) );
  AOI221_X1 U1843 ( .B1(b[19]), .B2(n1561), .C1(b[18]), .C2(n1562), .A(n2085), 
        .ZN(n2084) );
  OAI22_X1 U1844 ( .A1(n1564), .A2(n1721), .B1(n1640), .B2(n1722), .ZN(n2085)
         );
  INV_X1 U1845 ( .A(b[17]), .ZN(n1722) );
  INV_X1 U1846 ( .A(n1379), .ZN(n1721) );
  OAI222_X1 U1847 ( .A1(n2086), .A2(n2087), .B1(n2086), .B2(n2088), .C1(n2088), 
        .C2(n2087), .ZN(n2082) );
  INV_X1 U1848 ( .A(n588), .ZN(n2088) );
  XNOR2_X1 U1849 ( .A(n1743), .B(n2089), .ZN(n2087) );
  AOI221_X1 U1850 ( .B1(b[18]), .B2(n1561), .C1(b[17]), .C2(n1562), .A(n2090), 
        .ZN(n2089) );
  OAI22_X1 U1851 ( .A1(n1564), .A2(n1717), .B1(n1640), .B2(n1718), .ZN(n2090)
         );
  INV_X1 U1852 ( .A(b[16]), .ZN(n1718) );
  INV_X1 U1853 ( .A(n1380), .ZN(n1717) );
  AOI222_X1 U1854 ( .A1(n2091), .A2(n2092), .B1(n2091), .B2(n600), .C1(n600), 
        .C2(n2092), .ZN(n2086) );
  XNOR2_X1 U1855 ( .A(a[2]), .B(n2093), .ZN(n2092) );
  AOI221_X1 U1856 ( .B1(b[17]), .B2(n1561), .C1(b[16]), .C2(n1562), .A(n2094), 
        .ZN(n2093) );
  OAI22_X1 U1857 ( .A1(n1564), .A2(n1713), .B1(n1640), .B2(n1714), .ZN(n2094)
         );
  INV_X1 U1858 ( .A(b[15]), .ZN(n1714) );
  INV_X1 U1859 ( .A(n1381), .ZN(n1713) );
  OAI222_X1 U1860 ( .A1(n2095), .A2(n2096), .B1(n2095), .B2(n2097), .C1(n2097), 
        .C2(n2096), .ZN(n2091) );
  INV_X1 U1861 ( .A(n610), .ZN(n2097) );
  XNOR2_X1 U1862 ( .A(n1743), .B(n2098), .ZN(n2096) );
  AOI221_X1 U1863 ( .B1(b[16]), .B2(n1561), .C1(b[15]), .C2(n1562), .A(n2099), 
        .ZN(n2098) );
  OAI22_X1 U1864 ( .A1(n1564), .A2(n1709), .B1(n1640), .B2(n1710), .ZN(n2099)
         );
  INV_X1 U1865 ( .A(b[14]), .ZN(n1710) );
  INV_X1 U1866 ( .A(n1382), .ZN(n1709) );
  AOI222_X1 U1867 ( .A1(n2100), .A2(n2101), .B1(n2100), .B2(n620), .C1(n620), 
        .C2(n2101), .ZN(n2095) );
  XNOR2_X1 U1868 ( .A(a[2]), .B(n2102), .ZN(n2101) );
  AOI221_X1 U1869 ( .B1(b[15]), .B2(n1561), .C1(b[14]), .C2(n1562), .A(n2103), 
        .ZN(n2102) );
  OAI22_X1 U1870 ( .A1(n1564), .A2(n1705), .B1(n1640), .B2(n1706), .ZN(n2103)
         );
  INV_X1 U1871 ( .A(b[13]), .ZN(n1706) );
  INV_X1 U1872 ( .A(n1383), .ZN(n1705) );
  OAI222_X1 U1873 ( .A1(n2104), .A2(n2105), .B1(n2104), .B2(n2106), .C1(n2106), 
        .C2(n2105), .ZN(n2100) );
  INV_X1 U1874 ( .A(n630), .ZN(n2106) );
  XNOR2_X1 U1875 ( .A(n1743), .B(n2107), .ZN(n2105) );
  AOI221_X1 U1876 ( .B1(b[14]), .B2(n1561), .C1(b[13]), .C2(n1562), .A(n2108), 
        .ZN(n2107) );
  OAI22_X1 U1877 ( .A1(n1564), .A2(n1701), .B1(n1640), .B2(n1702), .ZN(n2108)
         );
  INV_X1 U1878 ( .A(b[12]), .ZN(n1702) );
  INV_X1 U1879 ( .A(n1384), .ZN(n1701) );
  AOI222_X1 U1880 ( .A1(n2109), .A2(n2110), .B1(n2109), .B2(n638), .C1(n638), 
        .C2(n2110), .ZN(n2104) );
  XNOR2_X1 U1881 ( .A(a[2]), .B(n2111), .ZN(n2110) );
  AOI221_X1 U1882 ( .B1(b[13]), .B2(n1561), .C1(b[12]), .C2(n1562), .A(n2112), 
        .ZN(n2111) );
  OAI22_X1 U1883 ( .A1(n1564), .A2(n1697), .B1(n1640), .B2(n1698), .ZN(n2112)
         );
  INV_X1 U1884 ( .A(b[11]), .ZN(n1698) );
  INV_X1 U1885 ( .A(n1385), .ZN(n1697) );
  OAI222_X1 U1886 ( .A1(n2113), .A2(n2114), .B1(n2113), .B2(n2115), .C1(n2115), 
        .C2(n2114), .ZN(n2109) );
  INV_X1 U1887 ( .A(n646), .ZN(n2115) );
  XNOR2_X1 U1888 ( .A(n1743), .B(n2116), .ZN(n2114) );
  AOI221_X1 U1889 ( .B1(b[12]), .B2(n1561), .C1(b[11]), .C2(n1562), .A(n2117), 
        .ZN(n2116) );
  OAI22_X1 U1890 ( .A1(n1564), .A2(n1693), .B1(n1640), .B2(n1694), .ZN(n2117)
         );
  INV_X1 U1891 ( .A(b[10]), .ZN(n1694) );
  INV_X1 U1892 ( .A(n1386), .ZN(n1693) );
  AOI222_X1 U1893 ( .A1(n2118), .A2(n2119), .B1(n2118), .B2(n654), .C1(n654), 
        .C2(n2119), .ZN(n2113) );
  XNOR2_X1 U1894 ( .A(a[2]), .B(n2120), .ZN(n2119) );
  AOI221_X1 U1895 ( .B1(b[11]), .B2(n1561), .C1(b[10]), .C2(n1562), .A(n2121), 
        .ZN(n2120) );
  OAI22_X1 U1896 ( .A1(n1564), .A2(n1689), .B1(n1640), .B2(n1690), .ZN(n2121)
         );
  INV_X1 U1897 ( .A(b[9]), .ZN(n1690) );
  INV_X1 U1898 ( .A(n1387), .ZN(n1689) );
  OAI222_X1 U1899 ( .A1(n2122), .A2(n2123), .B1(n2122), .B2(n2124), .C1(n2124), 
        .C2(n2123), .ZN(n2118) );
  INV_X1 U1900 ( .A(n660), .ZN(n2124) );
  XNOR2_X1 U1901 ( .A(n1743), .B(n2125), .ZN(n2123) );
  AOI221_X1 U1902 ( .B1(b[10]), .B2(n1561), .C1(b[9]), .C2(n1563), .A(n2126), 
        .ZN(n2125) );
  OAI22_X1 U1903 ( .A1(n1564), .A2(n1685), .B1(n1640), .B2(n1686), .ZN(n2126)
         );
  INV_X1 U1904 ( .A(b[8]), .ZN(n1686) );
  INV_X1 U1905 ( .A(n1388), .ZN(n1685) );
  AOI222_X1 U1906 ( .A1(n2127), .A2(n2128), .B1(n2127), .B2(n666), .C1(n666), 
        .C2(n2128), .ZN(n2122) );
  XNOR2_X1 U1907 ( .A(a[2]), .B(n2129), .ZN(n2128) );
  AOI221_X1 U1908 ( .B1(b[9]), .B2(n1561), .C1(b[8]), .C2(n1563), .A(n2130), 
        .ZN(n2129) );
  OAI22_X1 U1909 ( .A1(n1564), .A2(n1681), .B1(n1640), .B2(n1682), .ZN(n2130)
         );
  INV_X1 U1910 ( .A(b[7]), .ZN(n1682) );
  INV_X1 U1911 ( .A(n1389), .ZN(n1681) );
  OAI222_X1 U1912 ( .A1(n2131), .A2(n2132), .B1(n2131), .B2(n2133), .C1(n2133), 
        .C2(n2132), .ZN(n2127) );
  INV_X1 U1913 ( .A(n672), .ZN(n2133) );
  XNOR2_X1 U1914 ( .A(n1743), .B(n2134), .ZN(n2132) );
  AOI221_X1 U1915 ( .B1(b[8]), .B2(n1561), .C1(b[7]), .C2(n1562), .A(n2135), 
        .ZN(n2134) );
  OAI22_X1 U1916 ( .A1(n1564), .A2(n1677), .B1(n1640), .B2(n1678), .ZN(n2135)
         );
  INV_X1 U1917 ( .A(b[6]), .ZN(n1678) );
  INV_X1 U1918 ( .A(n1390), .ZN(n1677) );
  AOI222_X1 U1919 ( .A1(n2136), .A2(n2137), .B1(n2136), .B2(n676), .C1(n676), 
        .C2(n2137), .ZN(n2131) );
  XNOR2_X1 U1920 ( .A(a[2]), .B(n2138), .ZN(n2137) );
  AOI221_X1 U1921 ( .B1(b[7]), .B2(n1561), .C1(b[6]), .C2(n1563), .A(n2139), 
        .ZN(n2138) );
  OAI22_X1 U1922 ( .A1(n1564), .A2(n1673), .B1(n1640), .B2(n1674), .ZN(n2139)
         );
  INV_X1 U1923 ( .A(b[5]), .ZN(n1674) );
  INV_X1 U1924 ( .A(n1391), .ZN(n1673) );
  OAI222_X1 U1925 ( .A1(n2140), .A2(n2141), .B1(n2140), .B2(n2142), .C1(n2142), 
        .C2(n2141), .ZN(n2136) );
  INV_X1 U1926 ( .A(n680), .ZN(n2142) );
  XNOR2_X1 U1927 ( .A(n1743), .B(n2143), .ZN(n2141) );
  AOI221_X1 U1928 ( .B1(b[6]), .B2(n1561), .C1(b[5]), .C2(n1563), .A(n2144), 
        .ZN(n2143) );
  OAI22_X1 U1929 ( .A1(n1564), .A2(n1669), .B1(n1640), .B2(n1670), .ZN(n2144)
         );
  INV_X1 U1930 ( .A(b[4]), .ZN(n1670) );
  INV_X1 U1931 ( .A(n1392), .ZN(n1669) );
  AOI222_X1 U1932 ( .A1(n2145), .A2(n2146), .B1(n2145), .B2(n684), .C1(n684), 
        .C2(n2146), .ZN(n2140) );
  XNOR2_X1 U1933 ( .A(a[2]), .B(n2147), .ZN(n2146) );
  AOI221_X1 U1934 ( .B1(b[5]), .B2(n1561), .C1(b[4]), .C2(n1563), .A(n2148), 
        .ZN(n2147) );
  OAI22_X1 U1935 ( .A1(n1564), .A2(n1665), .B1(n1640), .B2(n1666), .ZN(n2148)
         );
  INV_X1 U1936 ( .A(b[3]), .ZN(n1666) );
  INV_X1 U1937 ( .A(n1393), .ZN(n1665) );
  OAI222_X1 U1938 ( .A1(n2149), .A2(n2150), .B1(n2149), .B2(n2151), .C1(n2151), 
        .C2(n2150), .ZN(n2145) );
  INV_X1 U1939 ( .A(n686), .ZN(n2151) );
  XNOR2_X1 U1940 ( .A(n1743), .B(n2152), .ZN(n2150) );
  AOI221_X1 U1941 ( .B1(b[4]), .B2(n1561), .C1(b[3]), .C2(n1563), .A(n2153), 
        .ZN(n2152) );
  OAI22_X1 U1942 ( .A1(n1564), .A2(n1661), .B1(n1640), .B2(n1662), .ZN(n2153)
         );
  INV_X1 U1943 ( .A(n1394), .ZN(n1661) );
  AOI222_X1 U1944 ( .A1(n2154), .A2(n2155), .B1(n2154), .B2(n688), .C1(n688), 
        .C2(n2155), .ZN(n2149) );
  XNOR2_X1 U1945 ( .A(a[2]), .B(n2156), .ZN(n2155) );
  AOI221_X1 U1946 ( .B1(b[3]), .B2(n1561), .C1(b[2]), .C2(n1563), .A(n2157), 
        .ZN(n2156) );
  OAI22_X1 U1947 ( .A1(n1564), .A2(n1658), .B1(n1640), .B2(n1650), .ZN(n2157)
         );
  INV_X1 U1948 ( .A(b[1]), .ZN(n1650) );
  INV_X1 U1949 ( .A(n1395), .ZN(n1658) );
  AND2_X1 U1950 ( .A1(n2161), .A2(n2162), .ZN(n2154) );
  AOI211_X1 U1951 ( .C1(b[1]), .C2(n1561), .A(n2163), .B(b[0]), .ZN(n2162) );
  OAI22_X1 U1952 ( .A1(n1535), .A2(n1662), .B1(n1564), .B2(n1651), .ZN(n2163)
         );
  INV_X1 U1953 ( .A(n1397), .ZN(n1651) );
  INV_X1 U1954 ( .A(b[2]), .ZN(n1662) );
  INV_X1 U1955 ( .A(a[0]), .ZN(n2159) );
  AOI221_X1 U1956 ( .B1(b[1]), .B2(n1563), .C1(n1396), .C2(n1555), .A(n1743), 
        .ZN(n2161) );
  XNOR2_X1 U1957 ( .A(a[1]), .B(n1743), .ZN(n2158) );
  INV_X1 U1958 ( .A(a[2]), .ZN(n1743) );
  NOR2_X1 U1959 ( .A1(n2160), .A2(a[0]), .ZN(n1637) );
  INV_X1 U1960 ( .A(a[1]), .ZN(n2160) );
endmodule


module iir_filter_DW_mult_tc_3 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(product[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(product[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(product[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(product[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(product[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(product[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(product[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(product[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(product[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(product[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(product[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(product[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(product[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(product[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(product[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(product[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(product[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(product[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(product[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(product[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(product[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(product[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(product[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1598), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1600), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1602), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1604), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1606), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1608), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1610), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(b[22]), .B(n1614), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(b[21]), .B(b[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(b[20]), .B(b[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(b[19]), .B(b[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(b[18]), .B(b[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(b[17]), .B(b[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(b[16]), .B(b[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(b[15]), .B(b[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(b[14]), .B(b[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(b[13]), .B(b[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(b[12]), .B(b[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(b[11]), .B(b[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(b[10]), .B(b[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(b[9]), .B(b[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(b[8]), .B(b[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(b[7]), .B(b[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(b[6]), .B(b[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(b[5]), .B(b[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(b[4]), .B(b[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(b[3]), .B(b[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(b[2]), .B(b[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(b[1]), .B(b[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(b[0]), .B(b[1]), .CO(n727), .S(n1397) );
  INV_X1 U1137 ( .A(n1533), .ZN(n1570) );
  INV_X1 U1138 ( .A(n1536), .ZN(n1568) );
  INV_X1 U1139 ( .A(n1535), .ZN(n1561) );
  INV_X1 U1140 ( .A(n1534), .ZN(n1569) );
  BUF_X1 U1141 ( .A(n1654), .Z(n1572) );
  INV_X1 U1142 ( .A(n1547), .ZN(n1560) );
  INV_X1 U1143 ( .A(n1544), .ZN(n1558) );
  INV_X1 U1144 ( .A(n1537), .ZN(n1580) );
  INV_X1 U1145 ( .A(n1551), .ZN(n1575) );
  INV_X1 U1146 ( .A(n1550), .ZN(n1585) );
  INV_X1 U1147 ( .A(n1548), .ZN(n1595) );
  INV_X1 U1148 ( .A(n1549), .ZN(n1590) );
  INV_X1 U1149 ( .A(n1538), .ZN(n1559) );
  INV_X1 U1150 ( .A(n1545), .ZN(n1593) );
  INV_X1 U1151 ( .A(n1553), .ZN(n1583) );
  INV_X1 U1152 ( .A(n1552), .ZN(n1588) );
  INV_X1 U1153 ( .A(n1546), .ZN(n1578) );
  INV_X1 U1154 ( .A(n1554), .ZN(n1573) );
  BUF_X1 U1155 ( .A(n1654), .Z(n1571) );
  BUF_X1 U1156 ( .A(n1629), .Z(n1557) );
  BUF_X1 U1157 ( .A(n1967), .Z(n1596) );
  BUF_X1 U1158 ( .A(n1912), .Z(n1591) );
  BUF_X1 U1159 ( .A(n1857), .Z(n1586) );
  BUF_X1 U1160 ( .A(n1802), .Z(n1581) );
  BUF_X1 U1161 ( .A(n1747), .Z(n1576) );
  BUF_X1 U1162 ( .A(n1912), .Z(n1592) );
  BUF_X1 U1163 ( .A(n1857), .Z(n1587) );
  BUF_X1 U1164 ( .A(n1802), .Z(n1582) );
  BUF_X1 U1165 ( .A(n1747), .Z(n1577) );
  BUF_X1 U1166 ( .A(n1967), .Z(n1597) );
  INV_X1 U1167 ( .A(n1615), .ZN(n1614) );
  INV_X1 U1168 ( .A(n1540), .ZN(n1589) );
  INV_X1 U1169 ( .A(n1541), .ZN(n1584) );
  INV_X1 U1170 ( .A(n1542), .ZN(n1579) );
  INV_X1 U1171 ( .A(n1543), .ZN(n1574) );
  BUF_X1 U1172 ( .A(n1629), .Z(n1556) );
  INV_X1 U1173 ( .A(n1539), .ZN(n1594) );
  NAND3_X1 U1174 ( .A1(n2157), .A2(n2158), .A3(n2159), .ZN(n1639) );
  INV_X1 U1175 ( .A(n1555), .ZN(n1564) );
  OR2_X1 U1176 ( .A1(n1738), .A2(n1739), .ZN(n1533) );
  OR2_X1 U1177 ( .A1(n1740), .A2(n1741), .ZN(n1534) );
  OR2_X1 U1178 ( .A1(n2158), .A2(n2157), .ZN(n1535) );
  AND2_X1 U1179 ( .A1(n1738), .A2(n1740), .ZN(n1536) );
  INV_X1 U1180 ( .A(n1611), .ZN(n1610) );
  INV_X1 U1181 ( .A(n1607), .ZN(n1606) );
  INV_X1 U1182 ( .A(n1609), .ZN(n1608) );
  INV_X1 U1183 ( .A(n1603), .ZN(n1602) );
  INV_X1 U1184 ( .A(n1605), .ZN(n1604) );
  OR2_X1 U1185 ( .A1(n1849), .A2(n1850), .ZN(n1537) );
  BUF_X1 U1186 ( .A(n1636), .Z(n1562) );
  BUF_X1 U1187 ( .A(n1636), .Z(n1563) );
  BUF_X1 U1188 ( .A(n1647), .Z(n1565) );
  BUF_X1 U1189 ( .A(n1647), .Z(n1566) );
  OR2_X1 U1190 ( .A1(n2068), .A2(n2067), .ZN(n1538) );
  OR2_X1 U1191 ( .A1(n2016), .A2(n2017), .ZN(n1539) );
  OR2_X1 U1192 ( .A1(n1961), .A2(n1962), .ZN(n1540) );
  OR2_X1 U1193 ( .A1(n1906), .A2(n1907), .ZN(n1541) );
  OR2_X1 U1194 ( .A1(n1851), .A2(n1852), .ZN(n1542) );
  OR2_X1 U1195 ( .A1(n1796), .A2(n1797), .ZN(n1543) );
  AND2_X1 U1196 ( .A1(n2070), .A2(n2068), .ZN(n1544) );
  AND2_X1 U1197 ( .A1(n2014), .A2(n2016), .ZN(n1545) );
  AND2_X1 U1198 ( .A1(n1849), .A2(n1851), .ZN(n1546) );
  OR2_X1 U1199 ( .A1(n2070), .A2(n2069), .ZN(n1547) );
  OR2_X1 U1200 ( .A1(n2014), .A2(n2015), .ZN(n1548) );
  OR2_X1 U1201 ( .A1(n1959), .A2(n1960), .ZN(n1549) );
  OR2_X1 U1202 ( .A1(n1904), .A2(n1905), .ZN(n1550) );
  OR2_X1 U1203 ( .A1(n1794), .A2(n1795), .ZN(n1551) );
  AND2_X1 U1204 ( .A1(n1959), .A2(n1961), .ZN(n1552) );
  AND2_X1 U1205 ( .A1(n1904), .A2(n1906), .ZN(n1553) );
  AND2_X1 U1206 ( .A1(n1794), .A2(n1796), .ZN(n1554) );
  BUF_X1 U1207 ( .A(n1647), .Z(n1567) );
  INV_X1 U1208 ( .A(n1599), .ZN(n1598) );
  AND2_X1 U1209 ( .A1(a[0]), .A2(n2157), .ZN(n1555) );
  BUF_X1 U1210 ( .A(a[20]), .Z(n1600) );
  INV_X1 U1211 ( .A(a[23]), .ZN(n1599) );
  INV_X1 U1212 ( .A(a[5]), .ZN(n1611) );
  INV_X1 U1213 ( .A(a[11]), .ZN(n1607) );
  INV_X1 U1214 ( .A(a[8]), .ZN(n1609) );
  INV_X1 U1215 ( .A(a[17]), .ZN(n1603) );
  INV_X1 U1216 ( .A(a[14]), .ZN(n1605) );
  BUF_X1 U1217 ( .A(a[20]), .Z(n1601) );
  CLKBUF_X1 U1218 ( .A(b[23]), .Z(n1612) );
  CLKBUF_X1 U1219 ( .A(b[23]), .Z(n1613) );
  INV_X1 U1220 ( .A(b[23]), .ZN(n1615) );
  INV_X1 U1221 ( .A(n1612), .ZN(n1616) );
  INV_X1 U1222 ( .A(n1612), .ZN(n1617) );
  INV_X1 U1223 ( .A(n1612), .ZN(n1618) );
  INV_X1 U1224 ( .A(n1613), .ZN(n1619) );
  INV_X1 U1225 ( .A(n1613), .ZN(n1620) );
  AOI21_X1 U1226 ( .B1(n1621), .B2(n1622), .A(n1623), .ZN(product[47]) );
  OAI22_X1 U1227 ( .A1(n1624), .A2(n1625), .B1(n1624), .B2(n1626), .ZN(n1623)
         );
  INV_X1 U1228 ( .A(n1622), .ZN(n1626) );
  AOI222_X1 U1229 ( .A1(n1627), .A2(n303), .B1(n1625), .B2(n303), .C1(n1627), 
        .C2(n1625), .ZN(n1624) );
  XOR2_X1 U1230 ( .A(n1628), .B(n1599), .Z(n1622) );
  OAI221_X1 U1231 ( .B1(n1617), .B2(n1557), .C1(n1620), .C2(n1558), .A(n1630), 
        .ZN(n1628) );
  OAI21_X1 U1232 ( .B1(n1559), .B2(n1560), .A(n1614), .ZN(n1630) );
  INV_X1 U1233 ( .A(n1625), .ZN(n1621) );
  XOR2_X1 U1234 ( .A(a[23]), .B(n1631), .Z(n1625) );
  AOI221_X1 U1235 ( .B1(n1613), .B2(n1559), .C1(n1560), .C2(n1614), .A(n1632), 
        .ZN(n1631) );
  OAI22_X1 U1236 ( .A1(n1558), .A2(n1633), .B1(n1557), .B2(n1634), .ZN(n1632)
         );
  XNOR2_X1 U1237 ( .A(a[2]), .B(n1635), .ZN(n908) );
  AOI221_X1 U1238 ( .B1(n1561), .B2(b[22]), .C1(n1563), .C2(b[21]), .A(n1637), 
        .ZN(n1635) );
  OAI22_X1 U1239 ( .A1(n1564), .A2(n1638), .B1(n1639), .B2(n1640), .ZN(n1637)
         );
  INV_X1 U1240 ( .A(n1376), .ZN(n1638) );
  XNOR2_X1 U1241 ( .A(a[2]), .B(n1641), .ZN(n907) );
  AOI221_X1 U1242 ( .B1(n1563), .B2(b[22]), .C1(n1555), .C2(n1375), .A(n1642), 
        .ZN(n1641) );
  OAI22_X1 U1243 ( .A1(n1643), .A2(n1639), .B1(n1617), .B2(n1535), .ZN(n1642)
         );
  XNOR2_X1 U1244 ( .A(a[2]), .B(n1644), .ZN(n906) );
  AOI221_X1 U1245 ( .B1(n1561), .B2(n1613), .C1(n1563), .C2(n1614), .A(n1645), 
        .ZN(n1644) );
  OAI22_X1 U1246 ( .A1(n1633), .A2(n1564), .B1(n1634), .B2(n1639), .ZN(n1645)
         );
  XNOR2_X1 U1247 ( .A(n1646), .B(n1611), .ZN(n904) );
  OAI22_X1 U1248 ( .A1(n1565), .A2(n1534), .B1(n1568), .B2(n1567), .ZN(n1646)
         );
  XNOR2_X1 U1249 ( .A(n1648), .B(n1611), .ZN(n903) );
  OAI222_X1 U1250 ( .A1(n1534), .A2(n1649), .B1(n1566), .B2(n1533), .C1(n1568), 
        .C2(n1650), .ZN(n1648) );
  XNOR2_X1 U1251 ( .A(n1610), .B(n1651), .ZN(n902) );
  AOI221_X1 U1252 ( .B1(b[2]), .B2(n1569), .C1(b[1]), .C2(n1570), .A(n1652), 
        .ZN(n1651) );
  OAI22_X1 U1253 ( .A1(n1568), .A2(n1653), .B1(n1565), .B2(n1572), .ZN(n1652)
         );
  XNOR2_X1 U1254 ( .A(n1610), .B(n1655), .ZN(n901) );
  AOI221_X1 U1255 ( .B1(b[3]), .B2(n1569), .C1(b[2]), .C2(n1570), .A(n1656), 
        .ZN(n1655) );
  OAI22_X1 U1256 ( .A1(n1568), .A2(n1657), .B1(n1649), .B2(n1572), .ZN(n1656)
         );
  XNOR2_X1 U1257 ( .A(n1610), .B(n1658), .ZN(n900) );
  AOI221_X1 U1258 ( .B1(b[4]), .B2(n1569), .C1(b[3]), .C2(n1570), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1259 ( .A1(n1568), .A2(n1660), .B1(n1661), .B2(n1572), .ZN(n1659)
         );
  XNOR2_X1 U1260 ( .A(n1610), .B(n1662), .ZN(n899) );
  AOI221_X1 U1261 ( .B1(b[5]), .B2(n1569), .C1(b[4]), .C2(n1570), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1262 ( .A1(n1568), .A2(n1664), .B1(n1572), .B2(n1665), .ZN(n1663)
         );
  XNOR2_X1 U1263 ( .A(n1610), .B(n1666), .ZN(n898) );
  AOI221_X1 U1264 ( .B1(b[6]), .B2(n1569), .C1(b[5]), .C2(n1570), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1265 ( .A1(n1568), .A2(n1668), .B1(n1572), .B2(n1669), .ZN(n1667)
         );
  XNOR2_X1 U1266 ( .A(n1610), .B(n1670), .ZN(n897) );
  AOI221_X1 U1267 ( .B1(b[7]), .B2(n1569), .C1(b[6]), .C2(n1570), .A(n1671), 
        .ZN(n1670) );
  OAI22_X1 U1268 ( .A1(n1568), .A2(n1672), .B1(n1572), .B2(n1673), .ZN(n1671)
         );
  XNOR2_X1 U1269 ( .A(n1610), .B(n1674), .ZN(n896) );
  AOI221_X1 U1270 ( .B1(b[8]), .B2(n1569), .C1(b[7]), .C2(n1570), .A(n1675), 
        .ZN(n1674) );
  OAI22_X1 U1271 ( .A1(n1568), .A2(n1676), .B1(n1571), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1272 ( .A(n1610), .B(n1678), .ZN(n895) );
  AOI221_X1 U1273 ( .B1(b[9]), .B2(n1569), .C1(b[8]), .C2(n1570), .A(n1679), 
        .ZN(n1678) );
  OAI22_X1 U1274 ( .A1(n1568), .A2(n1680), .B1(n1572), .B2(n1681), .ZN(n1679)
         );
  XNOR2_X1 U1275 ( .A(n1610), .B(n1682), .ZN(n894) );
  AOI221_X1 U1276 ( .B1(b[10]), .B2(n1569), .C1(b[9]), .C2(n1570), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1277 ( .A1(n1568), .A2(n1684), .B1(n1572), .B2(n1685), .ZN(n1683)
         );
  XNOR2_X1 U1278 ( .A(n1610), .B(n1686), .ZN(n893) );
  AOI221_X1 U1279 ( .B1(b[11]), .B2(n1569), .C1(b[10]), .C2(n1570), .A(n1687), 
        .ZN(n1686) );
  OAI22_X1 U1280 ( .A1(n1568), .A2(n1688), .B1(n1571), .B2(n1689), .ZN(n1687)
         );
  XNOR2_X1 U1281 ( .A(n1610), .B(n1690), .ZN(n892) );
  AOI221_X1 U1282 ( .B1(b[12]), .B2(n1569), .C1(b[11]), .C2(n1570), .A(n1691), 
        .ZN(n1690) );
  OAI22_X1 U1283 ( .A1(n1568), .A2(n1692), .B1(n1571), .B2(n1693), .ZN(n1691)
         );
  XNOR2_X1 U1284 ( .A(n1610), .B(n1694), .ZN(n891) );
  AOI221_X1 U1285 ( .B1(b[13]), .B2(n1569), .C1(b[12]), .C2(n1570), .A(n1695), 
        .ZN(n1694) );
  OAI22_X1 U1286 ( .A1(n1568), .A2(n1696), .B1(n1571), .B2(n1697), .ZN(n1695)
         );
  XNOR2_X1 U1287 ( .A(n1610), .B(n1698), .ZN(n890) );
  AOI221_X1 U1288 ( .B1(b[14]), .B2(n1569), .C1(b[13]), .C2(n1570), .A(n1699), 
        .ZN(n1698) );
  OAI22_X1 U1289 ( .A1(n1568), .A2(n1700), .B1(n1571), .B2(n1701), .ZN(n1699)
         );
  XNOR2_X1 U1290 ( .A(n1610), .B(n1702), .ZN(n889) );
  AOI221_X1 U1291 ( .B1(b[15]), .B2(n1569), .C1(b[14]), .C2(n1570), .A(n1703), 
        .ZN(n1702) );
  OAI22_X1 U1292 ( .A1(n1568), .A2(n1704), .B1(n1571), .B2(n1705), .ZN(n1703)
         );
  XNOR2_X1 U1293 ( .A(n1610), .B(n1706), .ZN(n888) );
  AOI221_X1 U1294 ( .B1(b[16]), .B2(n1569), .C1(b[15]), .C2(n1570), .A(n1707), 
        .ZN(n1706) );
  OAI22_X1 U1295 ( .A1(n1568), .A2(n1708), .B1(n1571), .B2(n1709), .ZN(n1707)
         );
  XNOR2_X1 U1296 ( .A(n1610), .B(n1710), .ZN(n887) );
  AOI221_X1 U1297 ( .B1(b[17]), .B2(n1569), .C1(b[16]), .C2(n1570), .A(n1711), 
        .ZN(n1710) );
  OAI22_X1 U1298 ( .A1(n1568), .A2(n1712), .B1(n1571), .B2(n1713), .ZN(n1711)
         );
  XNOR2_X1 U1299 ( .A(n1610), .B(n1714), .ZN(n886) );
  AOI221_X1 U1300 ( .B1(b[18]), .B2(n1569), .C1(b[17]), .C2(n1570), .A(n1715), 
        .ZN(n1714) );
  OAI22_X1 U1301 ( .A1(n1568), .A2(n1716), .B1(n1571), .B2(n1717), .ZN(n1715)
         );
  XNOR2_X1 U1302 ( .A(n1610), .B(n1718), .ZN(n885) );
  AOI221_X1 U1303 ( .B1(b[19]), .B2(n1569), .C1(b[18]), .C2(n1570), .A(n1719), 
        .ZN(n1718) );
  OAI22_X1 U1304 ( .A1(n1568), .A2(n1720), .B1(n1571), .B2(n1721), .ZN(n1719)
         );
  XNOR2_X1 U1305 ( .A(a[5]), .B(n1722), .ZN(n884) );
  AOI221_X1 U1306 ( .B1(n1569), .B2(b[20]), .C1(b[19]), .C2(n1570), .A(n1723), 
        .ZN(n1722) );
  OAI22_X1 U1307 ( .A1(n1568), .A2(n1724), .B1(n1571), .B2(n1725), .ZN(n1723)
         );
  XNOR2_X1 U1308 ( .A(a[5]), .B(n1726), .ZN(n883) );
  AOI221_X1 U1309 ( .B1(n1569), .B2(b[21]), .C1(n1570), .C2(b[20]), .A(n1727), 
        .ZN(n1726) );
  OAI22_X1 U1310 ( .A1(n1568), .A2(n1728), .B1(n1571), .B2(n1729), .ZN(n1727)
         );
  XNOR2_X1 U1311 ( .A(a[5]), .B(n1730), .ZN(n882) );
  AOI221_X1 U1312 ( .B1(n1569), .B2(b[22]), .C1(n1536), .C2(n1376), .A(n1731), 
        .ZN(n1730) );
  OAI22_X1 U1313 ( .A1(n1640), .A2(n1572), .B1(n1643), .B2(n1533), .ZN(n1731)
         );
  XNOR2_X1 U1314 ( .A(a[5]), .B(n1732), .ZN(n881) );
  AOI221_X1 U1315 ( .B1(n1570), .B2(b[22]), .C1(n1536), .C2(n1375), .A(n1733), 
        .ZN(n1732) );
  OAI22_X1 U1316 ( .A1(n1615), .A2(n1534), .B1(n1643), .B2(n1572), .ZN(n1733)
         );
  XNOR2_X1 U1317 ( .A(a[5]), .B(n1734), .ZN(n880) );
  AOI221_X1 U1318 ( .B1(n1569), .B2(n1613), .C1(n1570), .C2(n1614), .A(n1735), 
        .ZN(n1734) );
  OAI22_X1 U1319 ( .A1(n1633), .A2(n1568), .B1(n1634), .B2(n1572), .ZN(n1735)
         );
  XNOR2_X1 U1320 ( .A(n1610), .B(n1736), .ZN(n879) );
  OAI221_X1 U1321 ( .B1(n1616), .B2(n1572), .C1(n1620), .C2(n1568), .A(n1737), 
        .ZN(n1736) );
  OAI21_X1 U1322 ( .B1(n1569), .B2(n1570), .A(n1614), .ZN(n1737) );
  INV_X1 U1323 ( .A(n1741), .ZN(n1738) );
  NAND3_X1 U1324 ( .A1(n1741), .A2(n1740), .A3(n1739), .ZN(n1654) );
  XNOR2_X1 U1325 ( .A(a[3]), .B(a[4]), .ZN(n1739) );
  XNOR2_X1 U1326 ( .A(a[4]), .B(n1611), .ZN(n1740) );
  XOR2_X1 U1327 ( .A(a[3]), .B(n1742), .Z(n1741) );
  XNOR2_X1 U1328 ( .A(n1743), .B(n1609), .ZN(n878) );
  OAI22_X1 U1329 ( .A1(n1565), .A2(n1543), .B1(n1565), .B2(n1573), .ZN(n1743)
         );
  XNOR2_X1 U1330 ( .A(n1744), .B(n1609), .ZN(n877) );
  OAI222_X1 U1331 ( .A1(n1649), .A2(n1543), .B1(n1566), .B2(n1551), .C1(n1650), 
        .C2(n1573), .ZN(n1744) );
  XNOR2_X1 U1332 ( .A(n1608), .B(n1745), .ZN(n876) );
  AOI221_X1 U1333 ( .B1(n1574), .B2(b[2]), .C1(n1575), .C2(b[1]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1334 ( .A1(n1653), .A2(n1573), .B1(n1565), .B2(n1576), .ZN(n1746)
         );
  XNOR2_X1 U1335 ( .A(n1608), .B(n1748), .ZN(n875) );
  AOI221_X1 U1336 ( .B1(n1574), .B2(b[3]), .C1(n1575), .C2(b[2]), .A(n1749), 
        .ZN(n1748) );
  OAI22_X1 U1337 ( .A1(n1657), .A2(n1573), .B1(n1649), .B2(n1577), .ZN(n1749)
         );
  XNOR2_X1 U1338 ( .A(n1608), .B(n1750), .ZN(n874) );
  AOI221_X1 U1339 ( .B1(n1574), .B2(b[4]), .C1(n1575), .C2(b[3]), .A(n1751), 
        .ZN(n1750) );
  OAI22_X1 U1340 ( .A1(n1660), .A2(n1573), .B1(n1661), .B2(n1577), .ZN(n1751)
         );
  XNOR2_X1 U1341 ( .A(n1608), .B(n1752), .ZN(n873) );
  AOI221_X1 U1342 ( .B1(n1574), .B2(b[5]), .C1(n1575), .C2(b[4]), .A(n1753), 
        .ZN(n1752) );
  OAI22_X1 U1343 ( .A1(n1664), .A2(n1573), .B1(n1665), .B2(n1577), .ZN(n1753)
         );
  XNOR2_X1 U1344 ( .A(n1608), .B(n1754), .ZN(n872) );
  AOI221_X1 U1345 ( .B1(n1574), .B2(b[6]), .C1(n1575), .C2(b[5]), .A(n1755), 
        .ZN(n1754) );
  OAI22_X1 U1346 ( .A1(n1668), .A2(n1573), .B1(n1669), .B2(n1577), .ZN(n1755)
         );
  XNOR2_X1 U1347 ( .A(n1608), .B(n1756), .ZN(n871) );
  AOI221_X1 U1348 ( .B1(n1574), .B2(b[7]), .C1(n1575), .C2(b[6]), .A(n1757), 
        .ZN(n1756) );
  OAI22_X1 U1349 ( .A1(n1672), .A2(n1573), .B1(n1673), .B2(n1577), .ZN(n1757)
         );
  XNOR2_X1 U1350 ( .A(n1608), .B(n1758), .ZN(n870) );
  AOI221_X1 U1351 ( .B1(n1574), .B2(b[8]), .C1(n1575), .C2(b[7]), .A(n1759), 
        .ZN(n1758) );
  OAI22_X1 U1352 ( .A1(n1676), .A2(n1573), .B1(n1677), .B2(n1577), .ZN(n1759)
         );
  XNOR2_X1 U1353 ( .A(n1608), .B(n1760), .ZN(n869) );
  AOI221_X1 U1354 ( .B1(n1574), .B2(b[9]), .C1(n1575), .C2(b[8]), .A(n1761), 
        .ZN(n1760) );
  OAI22_X1 U1355 ( .A1(n1680), .A2(n1573), .B1(n1681), .B2(n1577), .ZN(n1761)
         );
  XNOR2_X1 U1356 ( .A(n1608), .B(n1762), .ZN(n868) );
  AOI221_X1 U1357 ( .B1(n1574), .B2(b[10]), .C1(n1575), .C2(b[9]), .A(n1763), 
        .ZN(n1762) );
  OAI22_X1 U1358 ( .A1(n1684), .A2(n1573), .B1(n1685), .B2(n1577), .ZN(n1763)
         );
  XNOR2_X1 U1359 ( .A(n1608), .B(n1764), .ZN(n867) );
  AOI221_X1 U1360 ( .B1(n1574), .B2(b[11]), .C1(n1575), .C2(b[10]), .A(n1765), 
        .ZN(n1764) );
  OAI22_X1 U1361 ( .A1(n1688), .A2(n1573), .B1(n1689), .B2(n1577), .ZN(n1765)
         );
  XNOR2_X1 U1362 ( .A(n1608), .B(n1766), .ZN(n866) );
  AOI221_X1 U1363 ( .B1(n1574), .B2(b[12]), .C1(n1575), .C2(b[11]), .A(n1767), 
        .ZN(n1766) );
  OAI22_X1 U1364 ( .A1(n1692), .A2(n1573), .B1(n1693), .B2(n1577), .ZN(n1767)
         );
  XNOR2_X1 U1365 ( .A(n1608), .B(n1768), .ZN(n865) );
  AOI221_X1 U1366 ( .B1(n1574), .B2(b[13]), .C1(n1575), .C2(b[12]), .A(n1769), 
        .ZN(n1768) );
  OAI22_X1 U1367 ( .A1(n1696), .A2(n1573), .B1(n1697), .B2(n1576), .ZN(n1769)
         );
  XNOR2_X1 U1368 ( .A(n1608), .B(n1770), .ZN(n864) );
  AOI221_X1 U1369 ( .B1(n1574), .B2(b[14]), .C1(n1575), .C2(b[13]), .A(n1771), 
        .ZN(n1770) );
  OAI22_X1 U1370 ( .A1(n1700), .A2(n1573), .B1(n1701), .B2(n1576), .ZN(n1771)
         );
  XNOR2_X1 U1371 ( .A(n1608), .B(n1772), .ZN(n863) );
  AOI221_X1 U1372 ( .B1(n1574), .B2(b[15]), .C1(n1575), .C2(b[14]), .A(n1773), 
        .ZN(n1772) );
  OAI22_X1 U1373 ( .A1(n1704), .A2(n1573), .B1(n1705), .B2(n1576), .ZN(n1773)
         );
  XNOR2_X1 U1374 ( .A(n1608), .B(n1774), .ZN(n862) );
  AOI221_X1 U1375 ( .B1(n1574), .B2(b[16]), .C1(n1575), .C2(b[15]), .A(n1775), 
        .ZN(n1774) );
  OAI22_X1 U1376 ( .A1(n1708), .A2(n1573), .B1(n1709), .B2(n1576), .ZN(n1775)
         );
  XNOR2_X1 U1377 ( .A(n1608), .B(n1776), .ZN(n861) );
  AOI221_X1 U1378 ( .B1(n1574), .B2(b[17]), .C1(n1575), .C2(b[16]), .A(n1777), 
        .ZN(n1776) );
  OAI22_X1 U1379 ( .A1(n1712), .A2(n1573), .B1(n1713), .B2(n1576), .ZN(n1777)
         );
  XNOR2_X1 U1380 ( .A(n1608), .B(n1778), .ZN(n860) );
  AOI221_X1 U1381 ( .B1(n1574), .B2(b[18]), .C1(n1575), .C2(b[17]), .A(n1779), 
        .ZN(n1778) );
  OAI22_X1 U1382 ( .A1(n1716), .A2(n1573), .B1(n1717), .B2(n1576), .ZN(n1779)
         );
  XNOR2_X1 U1383 ( .A(n1608), .B(n1780), .ZN(n859) );
  AOI221_X1 U1384 ( .B1(n1574), .B2(b[19]), .C1(n1575), .C2(b[18]), .A(n1781), 
        .ZN(n1780) );
  OAI22_X1 U1385 ( .A1(n1720), .A2(n1573), .B1(n1721), .B2(n1576), .ZN(n1781)
         );
  XNOR2_X1 U1386 ( .A(a[8]), .B(n1782), .ZN(n858) );
  AOI221_X1 U1387 ( .B1(n1574), .B2(b[20]), .C1(n1575), .C2(b[19]), .A(n1783), 
        .ZN(n1782) );
  OAI22_X1 U1388 ( .A1(n1724), .A2(n1573), .B1(n1725), .B2(n1576), .ZN(n1783)
         );
  XNOR2_X1 U1389 ( .A(a[8]), .B(n1784), .ZN(n857) );
  AOI221_X1 U1390 ( .B1(n1574), .B2(b[21]), .C1(n1575), .C2(b[20]), .A(n1785), 
        .ZN(n1784) );
  OAI22_X1 U1391 ( .A1(n1728), .A2(n1573), .B1(n1729), .B2(n1576), .ZN(n1785)
         );
  XNOR2_X1 U1392 ( .A(a[8]), .B(n1786), .ZN(n856) );
  AOI221_X1 U1393 ( .B1(n1574), .B2(b[22]), .C1(n1554), .C2(n1376), .A(n1787), 
        .ZN(n1786) );
  OAI22_X1 U1394 ( .A1(n1640), .A2(n1577), .B1(n1643), .B2(n1551), .ZN(n1787)
         );
  XNOR2_X1 U1395 ( .A(a[8]), .B(n1788), .ZN(n855) );
  AOI221_X1 U1396 ( .B1(n1575), .B2(b[22]), .C1(n1554), .C2(n1375), .A(n1789), 
        .ZN(n1788) );
  OAI22_X1 U1397 ( .A1(n1617), .A2(n1543), .B1(n1643), .B2(n1576), .ZN(n1789)
         );
  XNOR2_X1 U1398 ( .A(a[8]), .B(n1790), .ZN(n854) );
  AOI221_X1 U1399 ( .B1(n1574), .B2(n1613), .C1(n1575), .C2(n1614), .A(n1791), 
        .ZN(n1790) );
  OAI22_X1 U1400 ( .A1(n1633), .A2(n1573), .B1(n1634), .B2(n1576), .ZN(n1791)
         );
  XNOR2_X1 U1401 ( .A(n1608), .B(n1792), .ZN(n853) );
  OAI221_X1 U1402 ( .B1(n1616), .B2(n1577), .C1(n1617), .C2(n1573), .A(n1793), 
        .ZN(n1792) );
  OAI21_X1 U1403 ( .B1(n1574), .B2(n1575), .A(n1614), .ZN(n1793) );
  INV_X1 U1404 ( .A(n1797), .ZN(n1794) );
  NAND3_X1 U1405 ( .A1(n1797), .A2(n1796), .A3(n1795), .ZN(n1747) );
  XNOR2_X1 U1406 ( .A(a[6]), .B(a[7]), .ZN(n1795) );
  XNOR2_X1 U1407 ( .A(a[7]), .B(n1609), .ZN(n1796) );
  XOR2_X1 U1408 ( .A(a[6]), .B(n1611), .Z(n1797) );
  XNOR2_X1 U1409 ( .A(n1798), .B(n1607), .ZN(n852) );
  OAI22_X1 U1410 ( .A1(n1565), .A2(n1542), .B1(n1565), .B2(n1578), .ZN(n1798)
         );
  XNOR2_X1 U1411 ( .A(n1799), .B(n1607), .ZN(n851) );
  OAI222_X1 U1412 ( .A1(n1649), .A2(n1542), .B1(n1566), .B2(n1537), .C1(n1650), 
        .C2(n1578), .ZN(n1799) );
  XNOR2_X1 U1413 ( .A(n1606), .B(n1800), .ZN(n850) );
  AOI221_X1 U1414 ( .B1(n1579), .B2(b[2]), .C1(n1580), .C2(b[1]), .A(n1801), 
        .ZN(n1800) );
  OAI22_X1 U1415 ( .A1(n1653), .A2(n1578), .B1(n1566), .B2(n1581), .ZN(n1801)
         );
  XNOR2_X1 U1416 ( .A(n1606), .B(n1803), .ZN(n849) );
  AOI221_X1 U1417 ( .B1(n1579), .B2(b[3]), .C1(n1580), .C2(b[2]), .A(n1804), 
        .ZN(n1803) );
  OAI22_X1 U1418 ( .A1(n1657), .A2(n1578), .B1(n1649), .B2(n1582), .ZN(n1804)
         );
  XNOR2_X1 U1419 ( .A(n1606), .B(n1805), .ZN(n848) );
  AOI221_X1 U1420 ( .B1(n1579), .B2(b[4]), .C1(n1580), .C2(b[3]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1421 ( .A1(n1660), .A2(n1578), .B1(n1661), .B2(n1582), .ZN(n1806)
         );
  XNOR2_X1 U1422 ( .A(n1606), .B(n1807), .ZN(n847) );
  AOI221_X1 U1423 ( .B1(n1579), .B2(b[5]), .C1(n1580), .C2(b[4]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1424 ( .A1(n1664), .A2(n1578), .B1(n1665), .B2(n1582), .ZN(n1808)
         );
  XNOR2_X1 U1425 ( .A(n1606), .B(n1809), .ZN(n846) );
  AOI221_X1 U1426 ( .B1(n1579), .B2(b[6]), .C1(n1580), .C2(b[5]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1427 ( .A1(n1668), .A2(n1578), .B1(n1669), .B2(n1582), .ZN(n1810)
         );
  XNOR2_X1 U1428 ( .A(n1606), .B(n1811), .ZN(n845) );
  AOI221_X1 U1429 ( .B1(n1579), .B2(b[7]), .C1(n1580), .C2(b[6]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1430 ( .A1(n1672), .A2(n1578), .B1(n1673), .B2(n1582), .ZN(n1812)
         );
  XNOR2_X1 U1431 ( .A(n1606), .B(n1813), .ZN(n844) );
  AOI221_X1 U1432 ( .B1(n1579), .B2(b[8]), .C1(n1580), .C2(b[7]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1433 ( .A1(n1676), .A2(n1578), .B1(n1677), .B2(n1582), .ZN(n1814)
         );
  XNOR2_X1 U1434 ( .A(n1606), .B(n1815), .ZN(n843) );
  AOI221_X1 U1435 ( .B1(n1579), .B2(b[9]), .C1(n1580), .C2(b[8]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1436 ( .A1(n1680), .A2(n1578), .B1(n1681), .B2(n1582), .ZN(n1816)
         );
  XNOR2_X1 U1437 ( .A(n1606), .B(n1817), .ZN(n842) );
  AOI221_X1 U1438 ( .B1(n1579), .B2(b[10]), .C1(n1580), .C2(b[9]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1439 ( .A1(n1684), .A2(n1578), .B1(n1685), .B2(n1582), .ZN(n1818)
         );
  XNOR2_X1 U1440 ( .A(n1606), .B(n1819), .ZN(n841) );
  AOI221_X1 U1441 ( .B1(n1579), .B2(b[11]), .C1(n1580), .C2(b[10]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1442 ( .A1(n1688), .A2(n1578), .B1(n1689), .B2(n1582), .ZN(n1820)
         );
  XNOR2_X1 U1443 ( .A(n1606), .B(n1821), .ZN(n840) );
  AOI221_X1 U1444 ( .B1(n1579), .B2(b[12]), .C1(n1580), .C2(b[11]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1445 ( .A1(n1692), .A2(n1578), .B1(n1693), .B2(n1582), .ZN(n1822)
         );
  XNOR2_X1 U1446 ( .A(n1606), .B(n1823), .ZN(n839) );
  AOI221_X1 U1447 ( .B1(n1579), .B2(b[13]), .C1(n1580), .C2(b[12]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1448 ( .A1(n1696), .A2(n1578), .B1(n1697), .B2(n1581), .ZN(n1824)
         );
  XNOR2_X1 U1449 ( .A(n1606), .B(n1825), .ZN(n838) );
  AOI221_X1 U1450 ( .B1(n1579), .B2(b[14]), .C1(n1580), .C2(b[13]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1451 ( .A1(n1700), .A2(n1578), .B1(n1701), .B2(n1581), .ZN(n1826)
         );
  XNOR2_X1 U1452 ( .A(n1606), .B(n1827), .ZN(n837) );
  AOI221_X1 U1453 ( .B1(n1579), .B2(b[15]), .C1(n1580), .C2(b[14]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1454 ( .A1(n1704), .A2(n1578), .B1(n1705), .B2(n1581), .ZN(n1828)
         );
  XNOR2_X1 U1455 ( .A(n1606), .B(n1829), .ZN(n836) );
  AOI221_X1 U1456 ( .B1(n1579), .B2(b[16]), .C1(n1580), .C2(b[15]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1457 ( .A1(n1708), .A2(n1578), .B1(n1709), .B2(n1581), .ZN(n1830)
         );
  XNOR2_X1 U1458 ( .A(n1606), .B(n1831), .ZN(n835) );
  AOI221_X1 U1459 ( .B1(n1579), .B2(b[17]), .C1(n1580), .C2(b[16]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1460 ( .A1(n1712), .A2(n1578), .B1(n1713), .B2(n1581), .ZN(n1832)
         );
  XNOR2_X1 U1461 ( .A(n1606), .B(n1833), .ZN(n834) );
  AOI221_X1 U1462 ( .B1(n1579), .B2(b[18]), .C1(n1580), .C2(b[17]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1463 ( .A1(n1716), .A2(n1578), .B1(n1717), .B2(n1581), .ZN(n1834)
         );
  XNOR2_X1 U1464 ( .A(n1606), .B(n1835), .ZN(n833) );
  AOI221_X1 U1465 ( .B1(n1579), .B2(b[19]), .C1(n1580), .C2(b[18]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1466 ( .A1(n1720), .A2(n1578), .B1(n1721), .B2(n1581), .ZN(n1836)
         );
  XNOR2_X1 U1467 ( .A(n1606), .B(n1837), .ZN(n832) );
  AOI221_X1 U1468 ( .B1(n1579), .B2(b[20]), .C1(n1580), .C2(b[19]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1469 ( .A1(n1724), .A2(n1578), .B1(n1725), .B2(n1581), .ZN(n1838)
         );
  XNOR2_X1 U1470 ( .A(a[11]), .B(n1839), .ZN(n831) );
  AOI221_X1 U1471 ( .B1(n1579), .B2(b[21]), .C1(n1580), .C2(b[20]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1472 ( .A1(n1728), .A2(n1578), .B1(n1729), .B2(n1581), .ZN(n1840)
         );
  XNOR2_X1 U1473 ( .A(a[11]), .B(n1841), .ZN(n830) );
  AOI221_X1 U1474 ( .B1(n1579), .B2(b[22]), .C1(n1546), .C2(n1376), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1475 ( .A1(n1640), .A2(n1582), .B1(n1643), .B2(n1537), .ZN(n1842)
         );
  XNOR2_X1 U1476 ( .A(a[11]), .B(n1843), .ZN(n829) );
  AOI221_X1 U1477 ( .B1(n1580), .B2(b[22]), .C1(n1546), .C2(n1375), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1478 ( .A1(n1617), .A2(n1542), .B1(n1643), .B2(n1581), .ZN(n1844)
         );
  XNOR2_X1 U1479 ( .A(a[11]), .B(n1845), .ZN(n828) );
  AOI221_X1 U1480 ( .B1(n1579), .B2(n1614), .C1(n1580), .C2(n1614), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1481 ( .A1(n1633), .A2(n1578), .B1(n1634), .B2(n1581), .ZN(n1846)
         );
  XNOR2_X1 U1482 ( .A(a[11]), .B(n1847), .ZN(n827) );
  OAI221_X1 U1483 ( .B1(n1616), .B2(n1582), .C1(n1617), .C2(n1578), .A(n1848), 
        .ZN(n1847) );
  OAI21_X1 U1484 ( .B1(n1579), .B2(n1580), .A(n1614), .ZN(n1848) );
  INV_X1 U1485 ( .A(n1852), .ZN(n1849) );
  NAND3_X1 U1486 ( .A1(n1852), .A2(n1851), .A3(n1850), .ZN(n1802) );
  XNOR2_X1 U1487 ( .A(a[10]), .B(a[9]), .ZN(n1850) );
  XNOR2_X1 U1488 ( .A(a[10]), .B(n1607), .ZN(n1851) );
  XOR2_X1 U1489 ( .A(a[9]), .B(n1609), .Z(n1852) );
  XNOR2_X1 U1490 ( .A(n1853), .B(n1605), .ZN(n826) );
  OAI22_X1 U1491 ( .A1(n1565), .A2(n1541), .B1(n1565), .B2(n1583), .ZN(n1853)
         );
  XNOR2_X1 U1492 ( .A(n1854), .B(n1605), .ZN(n825) );
  OAI222_X1 U1493 ( .A1(n1649), .A2(n1541), .B1(n1566), .B2(n1550), .C1(n1650), 
        .C2(n1583), .ZN(n1854) );
  XNOR2_X1 U1494 ( .A(n1604), .B(n1855), .ZN(n824) );
  AOI221_X1 U1495 ( .B1(n1584), .B2(b[2]), .C1(n1585), .C2(b[1]), .A(n1856), 
        .ZN(n1855) );
  OAI22_X1 U1496 ( .A1(n1653), .A2(n1583), .B1(n1565), .B2(n1586), .ZN(n1856)
         );
  XNOR2_X1 U1497 ( .A(n1604), .B(n1858), .ZN(n823) );
  AOI221_X1 U1498 ( .B1(n1584), .B2(b[3]), .C1(n1585), .C2(b[2]), .A(n1859), 
        .ZN(n1858) );
  OAI22_X1 U1499 ( .A1(n1657), .A2(n1583), .B1(n1649), .B2(n1587), .ZN(n1859)
         );
  XNOR2_X1 U1500 ( .A(n1604), .B(n1860), .ZN(n822) );
  AOI221_X1 U1501 ( .B1(n1584), .B2(b[4]), .C1(n1585), .C2(b[3]), .A(n1861), 
        .ZN(n1860) );
  OAI22_X1 U1502 ( .A1(n1660), .A2(n1583), .B1(n1661), .B2(n1587), .ZN(n1861)
         );
  XNOR2_X1 U1503 ( .A(n1604), .B(n1862), .ZN(n821) );
  AOI221_X1 U1504 ( .B1(n1584), .B2(b[5]), .C1(n1585), .C2(b[4]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1505 ( .A1(n1664), .A2(n1583), .B1(n1665), .B2(n1587), .ZN(n1863)
         );
  XNOR2_X1 U1506 ( .A(n1604), .B(n1864), .ZN(n820) );
  AOI221_X1 U1507 ( .B1(n1584), .B2(b[6]), .C1(n1585), .C2(b[5]), .A(n1865), 
        .ZN(n1864) );
  OAI22_X1 U1508 ( .A1(n1668), .A2(n1583), .B1(n1669), .B2(n1587), .ZN(n1865)
         );
  XNOR2_X1 U1509 ( .A(n1604), .B(n1866), .ZN(n819) );
  AOI221_X1 U1510 ( .B1(n1584), .B2(b[7]), .C1(n1585), .C2(b[6]), .A(n1867), 
        .ZN(n1866) );
  OAI22_X1 U1511 ( .A1(n1672), .A2(n1583), .B1(n1673), .B2(n1587), .ZN(n1867)
         );
  XNOR2_X1 U1512 ( .A(n1604), .B(n1868), .ZN(n818) );
  AOI221_X1 U1513 ( .B1(n1584), .B2(b[8]), .C1(n1585), .C2(b[7]), .A(n1869), 
        .ZN(n1868) );
  OAI22_X1 U1514 ( .A1(n1676), .A2(n1583), .B1(n1677), .B2(n1587), .ZN(n1869)
         );
  XNOR2_X1 U1515 ( .A(n1604), .B(n1870), .ZN(n817) );
  AOI221_X1 U1516 ( .B1(n1584), .B2(b[9]), .C1(n1585), .C2(b[8]), .A(n1871), 
        .ZN(n1870) );
  OAI22_X1 U1517 ( .A1(n1680), .A2(n1583), .B1(n1681), .B2(n1587), .ZN(n1871)
         );
  XNOR2_X1 U1518 ( .A(n1604), .B(n1872), .ZN(n816) );
  AOI221_X1 U1519 ( .B1(n1584), .B2(b[10]), .C1(n1585), .C2(b[9]), .A(n1873), 
        .ZN(n1872) );
  OAI22_X1 U1520 ( .A1(n1684), .A2(n1583), .B1(n1685), .B2(n1587), .ZN(n1873)
         );
  XNOR2_X1 U1521 ( .A(n1604), .B(n1874), .ZN(n815) );
  AOI221_X1 U1522 ( .B1(n1584), .B2(b[11]), .C1(n1585), .C2(b[10]), .A(n1875), 
        .ZN(n1874) );
  OAI22_X1 U1523 ( .A1(n1688), .A2(n1583), .B1(n1689), .B2(n1587), .ZN(n1875)
         );
  XNOR2_X1 U1524 ( .A(n1604), .B(n1876), .ZN(n814) );
  AOI221_X1 U1525 ( .B1(n1584), .B2(b[12]), .C1(n1585), .C2(b[11]), .A(n1877), 
        .ZN(n1876) );
  OAI22_X1 U1526 ( .A1(n1692), .A2(n1583), .B1(n1693), .B2(n1587), .ZN(n1877)
         );
  XNOR2_X1 U1527 ( .A(n1604), .B(n1878), .ZN(n813) );
  AOI221_X1 U1528 ( .B1(n1584), .B2(b[13]), .C1(n1585), .C2(b[12]), .A(n1879), 
        .ZN(n1878) );
  OAI22_X1 U1529 ( .A1(n1696), .A2(n1583), .B1(n1697), .B2(n1586), .ZN(n1879)
         );
  XNOR2_X1 U1530 ( .A(n1604), .B(n1880), .ZN(n812) );
  AOI221_X1 U1531 ( .B1(n1584), .B2(b[14]), .C1(n1585), .C2(b[13]), .A(n1881), 
        .ZN(n1880) );
  OAI22_X1 U1532 ( .A1(n1700), .A2(n1583), .B1(n1701), .B2(n1586), .ZN(n1881)
         );
  XNOR2_X1 U1533 ( .A(n1604), .B(n1882), .ZN(n811) );
  AOI221_X1 U1534 ( .B1(n1584), .B2(b[15]), .C1(n1585), .C2(b[14]), .A(n1883), 
        .ZN(n1882) );
  OAI22_X1 U1535 ( .A1(n1704), .A2(n1583), .B1(n1705), .B2(n1586), .ZN(n1883)
         );
  XNOR2_X1 U1536 ( .A(n1604), .B(n1884), .ZN(n810) );
  AOI221_X1 U1537 ( .B1(n1584), .B2(b[16]), .C1(n1585), .C2(b[15]), .A(n1885), 
        .ZN(n1884) );
  OAI22_X1 U1538 ( .A1(n1708), .A2(n1583), .B1(n1709), .B2(n1586), .ZN(n1885)
         );
  XNOR2_X1 U1539 ( .A(n1604), .B(n1886), .ZN(n809) );
  AOI221_X1 U1540 ( .B1(n1584), .B2(b[17]), .C1(n1585), .C2(b[16]), .A(n1887), 
        .ZN(n1886) );
  OAI22_X1 U1541 ( .A1(n1712), .A2(n1583), .B1(n1713), .B2(n1586), .ZN(n1887)
         );
  XNOR2_X1 U1542 ( .A(n1604), .B(n1888), .ZN(n808) );
  AOI221_X1 U1543 ( .B1(n1584), .B2(b[18]), .C1(n1585), .C2(b[17]), .A(n1889), 
        .ZN(n1888) );
  OAI22_X1 U1544 ( .A1(n1716), .A2(n1583), .B1(n1717), .B2(n1586), .ZN(n1889)
         );
  XNOR2_X1 U1545 ( .A(n1604), .B(n1890), .ZN(n807) );
  AOI221_X1 U1546 ( .B1(n1584), .B2(b[19]), .C1(n1585), .C2(b[18]), .A(n1891), 
        .ZN(n1890) );
  OAI22_X1 U1547 ( .A1(n1720), .A2(n1583), .B1(n1721), .B2(n1586), .ZN(n1891)
         );
  XNOR2_X1 U1548 ( .A(n1604), .B(n1892), .ZN(n806) );
  AOI221_X1 U1549 ( .B1(n1584), .B2(b[20]), .C1(n1585), .C2(b[19]), .A(n1893), 
        .ZN(n1892) );
  OAI22_X1 U1550 ( .A1(n1724), .A2(n1583), .B1(n1725), .B2(n1586), .ZN(n1893)
         );
  XNOR2_X1 U1551 ( .A(a[14]), .B(n1894), .ZN(n805) );
  AOI221_X1 U1552 ( .B1(n1584), .B2(b[21]), .C1(n1585), .C2(b[20]), .A(n1895), 
        .ZN(n1894) );
  OAI22_X1 U1553 ( .A1(n1728), .A2(n1583), .B1(n1729), .B2(n1586), .ZN(n1895)
         );
  XNOR2_X1 U1554 ( .A(a[14]), .B(n1896), .ZN(n804) );
  AOI221_X1 U1555 ( .B1(n1584), .B2(b[22]), .C1(n1553), .C2(n1376), .A(n1897), 
        .ZN(n1896) );
  OAI22_X1 U1556 ( .A1(n1640), .A2(n1587), .B1(n1643), .B2(n1550), .ZN(n1897)
         );
  XNOR2_X1 U1557 ( .A(a[14]), .B(n1898), .ZN(n803) );
  AOI221_X1 U1558 ( .B1(n1585), .B2(b[22]), .C1(n1553), .C2(n1375), .A(n1899), 
        .ZN(n1898) );
  OAI22_X1 U1559 ( .A1(n1617), .A2(n1541), .B1(n1643), .B2(n1586), .ZN(n1899)
         );
  XNOR2_X1 U1560 ( .A(a[14]), .B(n1900), .ZN(n802) );
  AOI221_X1 U1561 ( .B1(n1584), .B2(n1614), .C1(n1585), .C2(n1614), .A(n1901), 
        .ZN(n1900) );
  OAI22_X1 U1562 ( .A1(n1633), .A2(n1583), .B1(n1634), .B2(n1586), .ZN(n1901)
         );
  XNOR2_X1 U1563 ( .A(a[14]), .B(n1902), .ZN(n801) );
  OAI221_X1 U1564 ( .B1(n1617), .B2(n1587), .C1(n1619), .C2(n1583), .A(n1903), 
        .ZN(n1902) );
  OAI21_X1 U1565 ( .B1(n1584), .B2(n1585), .A(n1614), .ZN(n1903) );
  INV_X1 U1566 ( .A(n1907), .ZN(n1904) );
  NAND3_X1 U1567 ( .A1(n1907), .A2(n1906), .A3(n1905), .ZN(n1857) );
  XNOR2_X1 U1568 ( .A(a[12]), .B(a[13]), .ZN(n1905) );
  XNOR2_X1 U1569 ( .A(a[13]), .B(n1605), .ZN(n1906) );
  XOR2_X1 U1570 ( .A(a[12]), .B(n1607), .Z(n1907) );
  XNOR2_X1 U1571 ( .A(n1908), .B(n1603), .ZN(n800) );
  OAI22_X1 U1572 ( .A1(n1565), .A2(n1540), .B1(n1566), .B2(n1588), .ZN(n1908)
         );
  XNOR2_X1 U1573 ( .A(n1909), .B(n1603), .ZN(n799) );
  OAI222_X1 U1574 ( .A1(n1649), .A2(n1540), .B1(n1566), .B2(n1549), .C1(n1650), 
        .C2(n1588), .ZN(n1909) );
  XNOR2_X1 U1575 ( .A(n1602), .B(n1910), .ZN(n798) );
  AOI221_X1 U1576 ( .B1(n1589), .B2(b[2]), .C1(n1590), .C2(b[1]), .A(n1911), 
        .ZN(n1910) );
  OAI22_X1 U1577 ( .A1(n1653), .A2(n1588), .B1(n1566), .B2(n1591), .ZN(n1911)
         );
  XNOR2_X1 U1578 ( .A(n1602), .B(n1913), .ZN(n797) );
  AOI221_X1 U1579 ( .B1(n1589), .B2(b[3]), .C1(n1590), .C2(b[2]), .A(n1914), 
        .ZN(n1913) );
  OAI22_X1 U1580 ( .A1(n1657), .A2(n1588), .B1(n1649), .B2(n1592), .ZN(n1914)
         );
  XNOR2_X1 U1581 ( .A(n1602), .B(n1915), .ZN(n796) );
  AOI221_X1 U1582 ( .B1(n1589), .B2(b[4]), .C1(n1590), .C2(b[3]), .A(n1916), 
        .ZN(n1915) );
  OAI22_X1 U1583 ( .A1(n1660), .A2(n1588), .B1(n1661), .B2(n1592), .ZN(n1916)
         );
  XNOR2_X1 U1584 ( .A(n1602), .B(n1917), .ZN(n795) );
  AOI221_X1 U1585 ( .B1(n1589), .B2(b[5]), .C1(n1590), .C2(b[4]), .A(n1918), 
        .ZN(n1917) );
  OAI22_X1 U1586 ( .A1(n1664), .A2(n1588), .B1(n1665), .B2(n1592), .ZN(n1918)
         );
  XNOR2_X1 U1587 ( .A(n1602), .B(n1919), .ZN(n794) );
  AOI221_X1 U1588 ( .B1(n1589), .B2(b[6]), .C1(n1590), .C2(b[5]), .A(n1920), 
        .ZN(n1919) );
  OAI22_X1 U1589 ( .A1(n1668), .A2(n1588), .B1(n1669), .B2(n1592), .ZN(n1920)
         );
  XNOR2_X1 U1590 ( .A(n1602), .B(n1921), .ZN(n793) );
  AOI221_X1 U1591 ( .B1(n1589), .B2(b[7]), .C1(n1590), .C2(b[6]), .A(n1922), 
        .ZN(n1921) );
  OAI22_X1 U1592 ( .A1(n1672), .A2(n1588), .B1(n1673), .B2(n1592), .ZN(n1922)
         );
  XNOR2_X1 U1593 ( .A(n1602), .B(n1923), .ZN(n792) );
  AOI221_X1 U1594 ( .B1(n1589), .B2(b[8]), .C1(n1590), .C2(b[7]), .A(n1924), 
        .ZN(n1923) );
  OAI22_X1 U1595 ( .A1(n1676), .A2(n1588), .B1(n1677), .B2(n1592), .ZN(n1924)
         );
  XNOR2_X1 U1596 ( .A(n1602), .B(n1925), .ZN(n791) );
  AOI221_X1 U1597 ( .B1(n1589), .B2(b[9]), .C1(n1590), .C2(b[8]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1598 ( .A1(n1680), .A2(n1588), .B1(n1681), .B2(n1592), .ZN(n1926)
         );
  XNOR2_X1 U1599 ( .A(n1602), .B(n1927), .ZN(n790) );
  AOI221_X1 U1600 ( .B1(n1589), .B2(b[10]), .C1(n1590), .C2(b[9]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1601 ( .A1(n1684), .A2(n1588), .B1(n1685), .B2(n1592), .ZN(n1928)
         );
  XNOR2_X1 U1602 ( .A(n1602), .B(n1929), .ZN(n789) );
  AOI221_X1 U1603 ( .B1(n1589), .B2(b[11]), .C1(n1590), .C2(b[10]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1604 ( .A1(n1688), .A2(n1588), .B1(n1689), .B2(n1592), .ZN(n1930)
         );
  XNOR2_X1 U1605 ( .A(n1602), .B(n1931), .ZN(n788) );
  AOI221_X1 U1606 ( .B1(n1589), .B2(b[12]), .C1(n1590), .C2(b[11]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1607 ( .A1(n1692), .A2(n1588), .B1(n1693), .B2(n1592), .ZN(n1932)
         );
  XNOR2_X1 U1608 ( .A(n1602), .B(n1933), .ZN(n787) );
  AOI221_X1 U1609 ( .B1(n1589), .B2(b[13]), .C1(n1590), .C2(b[12]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1610 ( .A1(n1696), .A2(n1588), .B1(n1697), .B2(n1591), .ZN(n1934)
         );
  XNOR2_X1 U1611 ( .A(n1602), .B(n1935), .ZN(n786) );
  AOI221_X1 U1612 ( .B1(n1589), .B2(b[14]), .C1(n1590), .C2(b[13]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1613 ( .A1(n1700), .A2(n1588), .B1(n1701), .B2(n1591), .ZN(n1936)
         );
  XNOR2_X1 U1614 ( .A(n1602), .B(n1937), .ZN(n785) );
  AOI221_X1 U1615 ( .B1(n1589), .B2(b[15]), .C1(n1590), .C2(b[14]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1616 ( .A1(n1704), .A2(n1588), .B1(n1705), .B2(n1591), .ZN(n1938)
         );
  XNOR2_X1 U1617 ( .A(n1602), .B(n1939), .ZN(n784) );
  AOI221_X1 U1618 ( .B1(n1589), .B2(b[16]), .C1(n1590), .C2(b[15]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1619 ( .A1(n1708), .A2(n1588), .B1(n1709), .B2(n1591), .ZN(n1940)
         );
  XNOR2_X1 U1620 ( .A(n1602), .B(n1941), .ZN(n783) );
  AOI221_X1 U1621 ( .B1(n1589), .B2(b[17]), .C1(n1590), .C2(b[16]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1622 ( .A1(n1712), .A2(n1588), .B1(n1713), .B2(n1591), .ZN(n1942)
         );
  XNOR2_X1 U1623 ( .A(n1602), .B(n1943), .ZN(n782) );
  AOI221_X1 U1624 ( .B1(n1589), .B2(b[18]), .C1(n1590), .C2(b[17]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1625 ( .A1(n1716), .A2(n1588), .B1(n1717), .B2(n1591), .ZN(n1944)
         );
  XNOR2_X1 U1626 ( .A(n1602), .B(n1945), .ZN(n781) );
  AOI221_X1 U1627 ( .B1(n1589), .B2(b[19]), .C1(n1590), .C2(b[18]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1628 ( .A1(n1720), .A2(n1588), .B1(n1721), .B2(n1591), .ZN(n1946)
         );
  XNOR2_X1 U1629 ( .A(n1602), .B(n1947), .ZN(n780) );
  AOI221_X1 U1630 ( .B1(n1589), .B2(b[20]), .C1(n1590), .C2(b[19]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1631 ( .A1(n1724), .A2(n1588), .B1(n1725), .B2(n1591), .ZN(n1948)
         );
  XNOR2_X1 U1632 ( .A(a[17]), .B(n1949), .ZN(n779) );
  AOI221_X1 U1633 ( .B1(n1589), .B2(b[21]), .C1(n1590), .C2(b[20]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1634 ( .A1(n1728), .A2(n1588), .B1(n1729), .B2(n1591), .ZN(n1950)
         );
  XNOR2_X1 U1635 ( .A(a[17]), .B(n1951), .ZN(n778) );
  AOI221_X1 U1636 ( .B1(n1589), .B2(b[22]), .C1(n1552), .C2(n1376), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1637 ( .A1(n1640), .A2(n1592), .B1(n1643), .B2(n1549), .ZN(n1952)
         );
  XNOR2_X1 U1638 ( .A(a[17]), .B(n1953), .ZN(n777) );
  AOI221_X1 U1639 ( .B1(n1590), .B2(b[22]), .C1(n1552), .C2(n1375), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1640 ( .A1(n1617), .A2(n1540), .B1(n1643), .B2(n1591), .ZN(n1954)
         );
  XNOR2_X1 U1641 ( .A(a[17]), .B(n1955), .ZN(n776) );
  AOI221_X1 U1642 ( .B1(n1589), .B2(n1613), .C1(n1590), .C2(n1614), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1643 ( .A1(n1633), .A2(n1588), .B1(n1634), .B2(n1591), .ZN(n1956)
         );
  XNOR2_X1 U1644 ( .A(a[17]), .B(n1957), .ZN(n775) );
  OAI221_X1 U1645 ( .B1(n1618), .B2(n1592), .C1(n1617), .C2(n1588), .A(n1958), 
        .ZN(n1957) );
  OAI21_X1 U1646 ( .B1(n1589), .B2(n1590), .A(n1614), .ZN(n1958) );
  INV_X1 U1647 ( .A(n1962), .ZN(n1959) );
  NAND3_X1 U1648 ( .A1(n1962), .A2(n1961), .A3(n1960), .ZN(n1912) );
  XNOR2_X1 U1649 ( .A(a[15]), .B(a[16]), .ZN(n1960) );
  XNOR2_X1 U1650 ( .A(a[16]), .B(n1603), .ZN(n1961) );
  XOR2_X1 U1651 ( .A(a[15]), .B(n1605), .Z(n1962) );
  XOR2_X1 U1652 ( .A(n1963), .B(n1600), .Z(n774) );
  OAI22_X1 U1653 ( .A1(n1565), .A2(n1539), .B1(n1566), .B2(n1593), .ZN(n1963)
         );
  XOR2_X1 U1654 ( .A(n1964), .B(n1600), .Z(n773) );
  OAI222_X1 U1655 ( .A1(n1649), .A2(n1539), .B1(n1566), .B2(n1548), .C1(n1650), 
        .C2(n1593), .ZN(n1964) );
  XNOR2_X1 U1656 ( .A(n1600), .B(n1965), .ZN(n772) );
  AOI221_X1 U1657 ( .B1(n1594), .B2(b[2]), .C1(n1595), .C2(b[1]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1658 ( .A1(n1653), .A2(n1593), .B1(n1566), .B2(n1596), .ZN(n1966)
         );
  XNOR2_X1 U1659 ( .A(n1600), .B(n1968), .ZN(n771) );
  AOI221_X1 U1660 ( .B1(n1594), .B2(b[3]), .C1(n1595), .C2(b[2]), .A(n1969), 
        .ZN(n1968) );
  OAI22_X1 U1661 ( .A1(n1657), .A2(n1593), .B1(n1649), .B2(n1597), .ZN(n1969)
         );
  XNOR2_X1 U1662 ( .A(n1600), .B(n1970), .ZN(n770) );
  AOI221_X1 U1663 ( .B1(n1594), .B2(b[4]), .C1(n1595), .C2(b[3]), .A(n1971), 
        .ZN(n1970) );
  OAI22_X1 U1664 ( .A1(n1660), .A2(n1593), .B1(n1661), .B2(n1597), .ZN(n1971)
         );
  XNOR2_X1 U1665 ( .A(n1600), .B(n1972), .ZN(n769) );
  AOI221_X1 U1666 ( .B1(n1594), .B2(b[5]), .C1(n1595), .C2(b[4]), .A(n1973), 
        .ZN(n1972) );
  OAI22_X1 U1667 ( .A1(n1664), .A2(n1593), .B1(n1665), .B2(n1597), .ZN(n1973)
         );
  XNOR2_X1 U1668 ( .A(n1600), .B(n1974), .ZN(n768) );
  AOI221_X1 U1669 ( .B1(n1594), .B2(b[6]), .C1(n1595), .C2(b[5]), .A(n1975), 
        .ZN(n1974) );
  OAI22_X1 U1670 ( .A1(n1668), .A2(n1593), .B1(n1669), .B2(n1597), .ZN(n1975)
         );
  XNOR2_X1 U1671 ( .A(n1600), .B(n1976), .ZN(n767) );
  AOI221_X1 U1672 ( .B1(n1594), .B2(b[7]), .C1(n1595), .C2(b[6]), .A(n1977), 
        .ZN(n1976) );
  OAI22_X1 U1673 ( .A1(n1672), .A2(n1593), .B1(n1673), .B2(n1597), .ZN(n1977)
         );
  XNOR2_X1 U1674 ( .A(n1600), .B(n1978), .ZN(n766) );
  AOI221_X1 U1675 ( .B1(n1594), .B2(b[8]), .C1(n1595), .C2(b[7]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1676 ( .A1(n1676), .A2(n1593), .B1(n1677), .B2(n1597), .ZN(n1979)
         );
  XNOR2_X1 U1677 ( .A(n1600), .B(n1980), .ZN(n765) );
  AOI221_X1 U1678 ( .B1(n1594), .B2(b[9]), .C1(n1595), .C2(b[8]), .A(n1981), 
        .ZN(n1980) );
  OAI22_X1 U1679 ( .A1(n1680), .A2(n1593), .B1(n1681), .B2(n1597), .ZN(n1981)
         );
  XNOR2_X1 U1680 ( .A(n1600), .B(n1982), .ZN(n764) );
  AOI221_X1 U1681 ( .B1(n1594), .B2(b[10]), .C1(n1595), .C2(b[9]), .A(n1983), 
        .ZN(n1982) );
  OAI22_X1 U1682 ( .A1(n1684), .A2(n1593), .B1(n1685), .B2(n1597), .ZN(n1983)
         );
  XNOR2_X1 U1683 ( .A(n1600), .B(n1984), .ZN(n763) );
  AOI221_X1 U1684 ( .B1(n1594), .B2(b[11]), .C1(n1595), .C2(b[10]), .A(n1985), 
        .ZN(n1984) );
  OAI22_X1 U1685 ( .A1(n1688), .A2(n1593), .B1(n1689), .B2(n1597), .ZN(n1985)
         );
  XNOR2_X1 U1686 ( .A(n1601), .B(n1986), .ZN(n762) );
  AOI221_X1 U1687 ( .B1(n1594), .B2(b[12]), .C1(n1595), .C2(b[11]), .A(n1987), 
        .ZN(n1986) );
  OAI22_X1 U1688 ( .A1(n1692), .A2(n1593), .B1(n1693), .B2(n1597), .ZN(n1987)
         );
  XNOR2_X1 U1689 ( .A(n1601), .B(n1988), .ZN(n761) );
  AOI221_X1 U1690 ( .B1(n1594), .B2(b[13]), .C1(n1595), .C2(b[12]), .A(n1989), 
        .ZN(n1988) );
  OAI22_X1 U1691 ( .A1(n1696), .A2(n1593), .B1(n1697), .B2(n1596), .ZN(n1989)
         );
  XNOR2_X1 U1692 ( .A(n1601), .B(n1990), .ZN(n760) );
  AOI221_X1 U1693 ( .B1(n1594), .B2(b[14]), .C1(n1595), .C2(b[13]), .A(n1991), 
        .ZN(n1990) );
  OAI22_X1 U1694 ( .A1(n1700), .A2(n1593), .B1(n1701), .B2(n1596), .ZN(n1991)
         );
  XNOR2_X1 U1695 ( .A(n1601), .B(n1992), .ZN(n759) );
  AOI221_X1 U1696 ( .B1(n1594), .B2(b[15]), .C1(n1595), .C2(b[14]), .A(n1993), 
        .ZN(n1992) );
  OAI22_X1 U1697 ( .A1(n1704), .A2(n1593), .B1(n1705), .B2(n1596), .ZN(n1993)
         );
  XNOR2_X1 U1698 ( .A(n1601), .B(n1994), .ZN(n758) );
  AOI221_X1 U1699 ( .B1(n1594), .B2(b[16]), .C1(n1595), .C2(b[15]), .A(n1995), 
        .ZN(n1994) );
  OAI22_X1 U1700 ( .A1(n1708), .A2(n1593), .B1(n1709), .B2(n1596), .ZN(n1995)
         );
  XNOR2_X1 U1701 ( .A(n1601), .B(n1996), .ZN(n757) );
  AOI221_X1 U1702 ( .B1(n1594), .B2(b[17]), .C1(n1595), .C2(b[16]), .A(n1997), 
        .ZN(n1996) );
  OAI22_X1 U1703 ( .A1(n1712), .A2(n1593), .B1(n1713), .B2(n1596), .ZN(n1997)
         );
  XNOR2_X1 U1704 ( .A(n1601), .B(n1998), .ZN(n756) );
  AOI221_X1 U1705 ( .B1(n1594), .B2(b[18]), .C1(n1595), .C2(b[17]), .A(n1999), 
        .ZN(n1998) );
  OAI22_X1 U1706 ( .A1(n1716), .A2(n1593), .B1(n1717), .B2(n1596), .ZN(n1999)
         );
  XNOR2_X1 U1707 ( .A(n1601), .B(n2000), .ZN(n755) );
  AOI221_X1 U1708 ( .B1(n1594), .B2(b[19]), .C1(n1595), .C2(b[18]), .A(n2001), 
        .ZN(n2000) );
  OAI22_X1 U1709 ( .A1(n1720), .A2(n1593), .B1(n1721), .B2(n1596), .ZN(n2001)
         );
  XNOR2_X1 U1710 ( .A(n1601), .B(n2002), .ZN(n754) );
  AOI221_X1 U1711 ( .B1(n1594), .B2(b[20]), .C1(n1595), .C2(b[19]), .A(n2003), 
        .ZN(n2002) );
  OAI22_X1 U1712 ( .A1(n1724), .A2(n1593), .B1(n1725), .B2(n1596), .ZN(n2003)
         );
  XNOR2_X1 U1713 ( .A(n1601), .B(n2004), .ZN(n753) );
  AOI221_X1 U1714 ( .B1(n1594), .B2(b[21]), .C1(n1595), .C2(b[20]), .A(n2005), 
        .ZN(n2004) );
  OAI22_X1 U1715 ( .A1(n1728), .A2(n1593), .B1(n1729), .B2(n1596), .ZN(n2005)
         );
  XNOR2_X1 U1716 ( .A(n1601), .B(n2006), .ZN(n752) );
  AOI221_X1 U1717 ( .B1(n1594), .B2(b[22]), .C1(n1545), .C2(n1376), .A(n2007), 
        .ZN(n2006) );
  OAI22_X1 U1718 ( .A1(n1640), .A2(n1597), .B1(n1643), .B2(n1548), .ZN(n2007)
         );
  XNOR2_X1 U1719 ( .A(n1601), .B(n2008), .ZN(n751) );
  AOI221_X1 U1720 ( .B1(n1595), .B2(b[22]), .C1(n1545), .C2(n1375), .A(n2009), 
        .ZN(n2008) );
  OAI22_X1 U1721 ( .A1(n1617), .A2(n1539), .B1(n1643), .B2(n1596), .ZN(n2009)
         );
  XNOR2_X1 U1722 ( .A(n1601), .B(n2010), .ZN(n750) );
  AOI221_X1 U1723 ( .B1(n1594), .B2(n1612), .C1(n1595), .C2(n1614), .A(n2011), 
        .ZN(n2010) );
  OAI22_X1 U1724 ( .A1(n1633), .A2(n1593), .B1(n1634), .B2(n1596), .ZN(n2011)
         );
  INV_X1 U1725 ( .A(b[22]), .ZN(n1634) );
  INV_X1 U1726 ( .A(n1374), .ZN(n1633) );
  XNOR2_X1 U1727 ( .A(n1600), .B(n2012), .ZN(n749) );
  OAI221_X1 U1728 ( .B1(n1617), .B2(n1597), .C1(n1619), .C2(n1593), .A(n2013), 
        .ZN(n2012) );
  OAI21_X1 U1729 ( .B1(n1594), .B2(n1595), .A(n1614), .ZN(n2013) );
  INV_X1 U1730 ( .A(n2017), .ZN(n2014) );
  NAND3_X1 U1731 ( .A1(n2017), .A2(n2016), .A3(n2015), .ZN(n1967) );
  XNOR2_X1 U1732 ( .A(a[18]), .B(a[19]), .ZN(n2015) );
  XOR2_X1 U1733 ( .A(a[19]), .B(n1600), .Z(n2016) );
  XOR2_X1 U1734 ( .A(a[18]), .B(n1603), .Z(n2017) );
  XNOR2_X1 U1735 ( .A(n2018), .B(n1599), .ZN(n748) );
  OAI22_X1 U1736 ( .A1(n1538), .A2(n1567), .B1(n1558), .B2(n1567), .ZN(n2018)
         );
  XNOR2_X1 U1737 ( .A(n2019), .B(n1599), .ZN(n747) );
  OAI222_X1 U1738 ( .A1(n1538), .A2(n1649), .B1(n1547), .B2(n1566), .C1(n1558), 
        .C2(n1650), .ZN(n2019) );
  XNOR2_X1 U1739 ( .A(n1598), .B(n2020), .ZN(n746) );
  AOI221_X1 U1740 ( .B1(b[2]), .B2(n1559), .C1(b[1]), .C2(n1560), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1741 ( .A1(n1558), .A2(n1653), .B1(n1557), .B2(n1567), .ZN(n2021)
         );
  INV_X1 U1742 ( .A(b[0]), .ZN(n1647) );
  INV_X1 U1743 ( .A(n1396), .ZN(n1653) );
  XNOR2_X1 U1744 ( .A(n1598), .B(n2022), .ZN(n745) );
  AOI221_X1 U1745 ( .B1(b[3]), .B2(n1559), .C1(b[2]), .C2(n1560), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1746 ( .A1(n1558), .A2(n1657), .B1(n1557), .B2(n1649), .ZN(n2023)
         );
  XNOR2_X1 U1747 ( .A(n1598), .B(n2024), .ZN(n744) );
  AOI221_X1 U1748 ( .B1(b[4]), .B2(n1559), .C1(b[3]), .C2(n1560), .A(n2025), 
        .ZN(n2024) );
  OAI22_X1 U1749 ( .A1(n1558), .A2(n1660), .B1(n1557), .B2(n1661), .ZN(n2025)
         );
  XNOR2_X1 U1750 ( .A(n1598), .B(n2026), .ZN(n743) );
  AOI221_X1 U1751 ( .B1(b[5]), .B2(n1559), .C1(b[4]), .C2(n1560), .A(n2027), 
        .ZN(n2026) );
  OAI22_X1 U1752 ( .A1(n1558), .A2(n1664), .B1(n1557), .B2(n1665), .ZN(n2027)
         );
  XNOR2_X1 U1753 ( .A(n1598), .B(n2028), .ZN(n742) );
  AOI221_X1 U1754 ( .B1(b[6]), .B2(n1559), .C1(b[5]), .C2(n1560), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1755 ( .A1(n1558), .A2(n1668), .B1(n1557), .B2(n1669), .ZN(n2029)
         );
  XNOR2_X1 U1756 ( .A(n1598), .B(n2030), .ZN(n741) );
  AOI221_X1 U1757 ( .B1(b[7]), .B2(n1559), .C1(b[6]), .C2(n1560), .A(n2031), 
        .ZN(n2030) );
  OAI22_X1 U1758 ( .A1(n1558), .A2(n1672), .B1(n1557), .B2(n1673), .ZN(n2031)
         );
  XNOR2_X1 U1759 ( .A(n1598), .B(n2032), .ZN(n740) );
  AOI221_X1 U1760 ( .B1(b[9]), .B2(n1559), .C1(b[8]), .C2(n1560), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1761 ( .A1(n1558), .A2(n1680), .B1(n1557), .B2(n1681), .ZN(n2033)
         );
  XNOR2_X1 U1762 ( .A(n1598), .B(n2034), .ZN(n739) );
  AOI221_X1 U1763 ( .B1(b[10]), .B2(n1559), .C1(b[9]), .C2(n1560), .A(n2035), 
        .ZN(n2034) );
  OAI22_X1 U1764 ( .A1(n1558), .A2(n1684), .B1(n1557), .B2(n1685), .ZN(n2035)
         );
  XNOR2_X1 U1765 ( .A(n1598), .B(n2036), .ZN(n738) );
  AOI221_X1 U1766 ( .B1(b[12]), .B2(n1559), .C1(b[11]), .C2(n1560), .A(n2037), 
        .ZN(n2036) );
  OAI22_X1 U1767 ( .A1(n1558), .A2(n1692), .B1(n1557), .B2(n1693), .ZN(n2037)
         );
  XNOR2_X1 U1768 ( .A(n1598), .B(n2038), .ZN(n737) );
  AOI221_X1 U1769 ( .B1(b[13]), .B2(n1559), .C1(b[12]), .C2(n1560), .A(n2039), 
        .ZN(n2038) );
  OAI22_X1 U1770 ( .A1(n1558), .A2(n1696), .B1(n1557), .B2(n1697), .ZN(n2039)
         );
  XNOR2_X1 U1771 ( .A(n1598), .B(n2040), .ZN(n736) );
  AOI221_X1 U1772 ( .B1(b[14]), .B2(n1559), .C1(b[13]), .C2(n1560), .A(n2041), 
        .ZN(n2040) );
  OAI22_X1 U1773 ( .A1(n1558), .A2(n1700), .B1(n1556), .B2(n1701), .ZN(n2041)
         );
  XNOR2_X1 U1774 ( .A(n1598), .B(n2042), .ZN(n735) );
  AOI221_X1 U1775 ( .B1(b[15]), .B2(n1559), .C1(b[14]), .C2(n1560), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1776 ( .A1(n1558), .A2(n1704), .B1(n1556), .B2(n1705), .ZN(n2043)
         );
  XNOR2_X1 U1777 ( .A(n1598), .B(n2044), .ZN(n734) );
  AOI221_X1 U1778 ( .B1(b[16]), .B2(n1559), .C1(b[15]), .C2(n1560), .A(n2045), 
        .ZN(n2044) );
  OAI22_X1 U1779 ( .A1(n1558), .A2(n1708), .B1(n1556), .B2(n1709), .ZN(n2045)
         );
  XNOR2_X1 U1780 ( .A(n1598), .B(n2046), .ZN(n733) );
  AOI221_X1 U1781 ( .B1(b[18]), .B2(n1559), .C1(b[17]), .C2(n1560), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1782 ( .A1(n1558), .A2(n1716), .B1(n1556), .B2(n1717), .ZN(n2047)
         );
  XNOR2_X1 U1783 ( .A(n1598), .B(n2048), .ZN(n732) );
  AOI221_X1 U1784 ( .B1(b[19]), .B2(n1559), .C1(b[18]), .C2(n1560), .A(n2049), 
        .ZN(n2048) );
  OAI22_X1 U1785 ( .A1(n1558), .A2(n1720), .B1(n1556), .B2(n1721), .ZN(n2049)
         );
  XNOR2_X1 U1786 ( .A(n1598), .B(n2050), .ZN(n731) );
  AOI221_X1 U1787 ( .B1(b[20]), .B2(n1559), .C1(b[19]), .C2(n1560), .A(n2051), 
        .ZN(n2050) );
  OAI22_X1 U1788 ( .A1(n1558), .A2(n1724), .B1(n1556), .B2(n1725), .ZN(n2051)
         );
  XNOR2_X1 U1789 ( .A(a[23]), .B(n2052), .ZN(n730) );
  AOI221_X1 U1790 ( .B1(b[21]), .B2(n1559), .C1(b[20]), .C2(n1560), .A(n2053), 
        .ZN(n2052) );
  OAI22_X1 U1791 ( .A1(n1558), .A2(n1728), .B1(n1556), .B2(n1729), .ZN(n2053)
         );
  XNOR2_X1 U1792 ( .A(a[23]), .B(n2054), .ZN(n729) );
  AOI221_X1 U1793 ( .B1(b[22]), .B2(n1559), .C1(n1376), .C2(n1544), .A(n2055), 
        .ZN(n2054) );
  OAI22_X1 U1794 ( .A1(n1556), .A2(n1640), .B1(n1547), .B2(n1643), .ZN(n2055)
         );
  INV_X1 U1795 ( .A(b[20]), .ZN(n1640) );
  XNOR2_X1 U1796 ( .A(n519), .B(n2056), .ZN(n506) );
  INV_X1 U1797 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1798 ( .A1(n2056), .A2(n519), .ZN(n493) );
  XOR2_X1 U1799 ( .A(n2057), .B(n1742), .Z(n2056) );
  OAI221_X1 U1800 ( .B1(n1618), .B2(n1639), .C1(n1619), .C2(n1564), .A(n2058), 
        .ZN(n2057) );
  OAI21_X1 U1801 ( .B1(n1561), .B2(n1563), .A(n1614), .ZN(n2058) );
  INV_X1 U1802 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1803 ( .A(n1598), .B(n2059), .Z(n454) );
  AOI221_X1 U1804 ( .B1(b[8]), .B2(n1559), .C1(b[7]), .C2(n1560), .A(n2060), 
        .ZN(n2059) );
  OAI22_X1 U1805 ( .A1(n1558), .A2(n1676), .B1(n1556), .B2(n1677), .ZN(n2060)
         );
  INV_X1 U1806 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1807 ( .A(n1598), .B(n2061), .Z(n421) );
  AOI221_X1 U1808 ( .B1(b[11]), .B2(n1559), .C1(b[10]), .C2(n1560), .A(n2062), 
        .ZN(n2061) );
  OAI22_X1 U1809 ( .A1(n1558), .A2(n1688), .B1(n1556), .B2(n1689), .ZN(n2062)
         );
  INV_X1 U1810 ( .A(n387), .ZN(n395) );
  INV_X1 U1811 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1812 ( .A(n1598), .B(n2063), .Z(n374) );
  AOI221_X1 U1813 ( .B1(b[17]), .B2(n1559), .C1(b[16]), .C2(n1560), .A(n2064), 
        .ZN(n2063) );
  OAI22_X1 U1814 ( .A1(n1558), .A2(n1712), .B1(n1556), .B2(n1713), .ZN(n2064)
         );
  INV_X1 U1815 ( .A(n356), .ZN(n360) );
  INV_X1 U1816 ( .A(n1627), .ZN(n351) );
  XOR2_X1 U1817 ( .A(n1599), .B(n2065), .Z(n1627) );
  AOI221_X1 U1818 ( .B1(b[22]), .B2(n1560), .C1(n1375), .C2(n1544), .A(n2066), 
        .ZN(n2065) );
  OAI22_X1 U1819 ( .A1(n1538), .A2(n1618), .B1(n1556), .B2(n1643), .ZN(n2066)
         );
  INV_X1 U1820 ( .A(b[21]), .ZN(n1643) );
  NAND3_X1 U1821 ( .A1(n2067), .A2(n2068), .A3(n2069), .ZN(n1629) );
  XNOR2_X1 U1822 ( .A(a[22]), .B(n1599), .ZN(n2068) );
  XNOR2_X1 U1823 ( .A(a[21]), .B(a[22]), .ZN(n2069) );
  INV_X1 U1824 ( .A(n2067), .ZN(n2070) );
  XNOR2_X1 U1825 ( .A(a[21]), .B(n1600), .ZN(n2067) );
  OAI222_X1 U1826 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n2073), .C1(n2073), 
        .C2(n2072), .ZN(n326) );
  INV_X1 U1827 ( .A(n550), .ZN(n2073) );
  XNOR2_X1 U1828 ( .A(n1742), .B(n2074), .ZN(n2072) );
  AOI221_X1 U1829 ( .B1(n1561), .B2(b[21]), .C1(b[20]), .C2(n1562), .A(n2075), 
        .ZN(n2074) );
  OAI22_X1 U1830 ( .A1(n1564), .A2(n1728), .B1(n1639), .B2(n1729), .ZN(n2075)
         );
  INV_X1 U1831 ( .A(b[19]), .ZN(n1729) );
  INV_X1 U1832 ( .A(n1377), .ZN(n1728) );
  AOI222_X1 U1833 ( .A1(n2076), .A2(n2077), .B1(n2076), .B2(n564), .C1(n564), 
        .C2(n2077), .ZN(n2071) );
  XNOR2_X1 U1834 ( .A(a[2]), .B(n2078), .ZN(n2077) );
  AOI221_X1 U1835 ( .B1(b[20]), .B2(n1561), .C1(b[19]), .C2(n1562), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1836 ( .A1(n1564), .A2(n1724), .B1(n1639), .B2(n1725), .ZN(n2079)
         );
  INV_X1 U1837 ( .A(b[18]), .ZN(n1725) );
  INV_X1 U1838 ( .A(n1378), .ZN(n1724) );
  INV_X1 U1839 ( .A(n2080), .ZN(n2076) );
  AOI222_X1 U1840 ( .A1(n2081), .A2(n2082), .B1(n2081), .B2(n576), .C1(n576), 
        .C2(n2082), .ZN(n2080) );
  XNOR2_X1 U1841 ( .A(a[2]), .B(n2083), .ZN(n2082) );
  AOI221_X1 U1842 ( .B1(b[19]), .B2(n1561), .C1(b[18]), .C2(n1562), .A(n2084), 
        .ZN(n2083) );
  OAI22_X1 U1843 ( .A1(n1564), .A2(n1720), .B1(n1639), .B2(n1721), .ZN(n2084)
         );
  INV_X1 U1844 ( .A(b[17]), .ZN(n1721) );
  INV_X1 U1845 ( .A(n1379), .ZN(n1720) );
  OAI222_X1 U1846 ( .A1(n2085), .A2(n2086), .B1(n2085), .B2(n2087), .C1(n2087), 
        .C2(n2086), .ZN(n2081) );
  INV_X1 U1847 ( .A(n588), .ZN(n2087) );
  XNOR2_X1 U1848 ( .A(n1742), .B(n2088), .ZN(n2086) );
  AOI221_X1 U1849 ( .B1(b[18]), .B2(n1561), .C1(b[17]), .C2(n1562), .A(n2089), 
        .ZN(n2088) );
  OAI22_X1 U1850 ( .A1(n1564), .A2(n1716), .B1(n1639), .B2(n1717), .ZN(n2089)
         );
  INV_X1 U1851 ( .A(b[16]), .ZN(n1717) );
  INV_X1 U1852 ( .A(n1380), .ZN(n1716) );
  AOI222_X1 U1853 ( .A1(n2090), .A2(n2091), .B1(n2090), .B2(n600), .C1(n600), 
        .C2(n2091), .ZN(n2085) );
  XNOR2_X1 U1854 ( .A(a[2]), .B(n2092), .ZN(n2091) );
  AOI221_X1 U1855 ( .B1(b[17]), .B2(n1561), .C1(b[16]), .C2(n1562), .A(n2093), 
        .ZN(n2092) );
  OAI22_X1 U1856 ( .A1(n1564), .A2(n1712), .B1(n1639), .B2(n1713), .ZN(n2093)
         );
  INV_X1 U1857 ( .A(b[15]), .ZN(n1713) );
  INV_X1 U1858 ( .A(n1381), .ZN(n1712) );
  OAI222_X1 U1859 ( .A1(n2094), .A2(n2095), .B1(n2094), .B2(n2096), .C1(n2096), 
        .C2(n2095), .ZN(n2090) );
  INV_X1 U1860 ( .A(n610), .ZN(n2096) );
  XNOR2_X1 U1861 ( .A(n1742), .B(n2097), .ZN(n2095) );
  AOI221_X1 U1862 ( .B1(b[16]), .B2(n1561), .C1(b[15]), .C2(n1562), .A(n2098), 
        .ZN(n2097) );
  OAI22_X1 U1863 ( .A1(n1564), .A2(n1708), .B1(n1639), .B2(n1709), .ZN(n2098)
         );
  INV_X1 U1864 ( .A(b[14]), .ZN(n1709) );
  INV_X1 U1865 ( .A(n1382), .ZN(n1708) );
  AOI222_X1 U1866 ( .A1(n2099), .A2(n2100), .B1(n2099), .B2(n620), .C1(n620), 
        .C2(n2100), .ZN(n2094) );
  XNOR2_X1 U1867 ( .A(a[2]), .B(n2101), .ZN(n2100) );
  AOI221_X1 U1868 ( .B1(b[15]), .B2(n1561), .C1(b[14]), .C2(n1562), .A(n2102), 
        .ZN(n2101) );
  OAI22_X1 U1869 ( .A1(n1564), .A2(n1704), .B1(n1639), .B2(n1705), .ZN(n2102)
         );
  INV_X1 U1870 ( .A(b[13]), .ZN(n1705) );
  INV_X1 U1871 ( .A(n1383), .ZN(n1704) );
  OAI222_X1 U1872 ( .A1(n2103), .A2(n2104), .B1(n2103), .B2(n2105), .C1(n2105), 
        .C2(n2104), .ZN(n2099) );
  INV_X1 U1873 ( .A(n630), .ZN(n2105) );
  XNOR2_X1 U1874 ( .A(n1742), .B(n2106), .ZN(n2104) );
  AOI221_X1 U1875 ( .B1(b[14]), .B2(n1561), .C1(b[13]), .C2(n1562), .A(n2107), 
        .ZN(n2106) );
  OAI22_X1 U1876 ( .A1(n1564), .A2(n1700), .B1(n1639), .B2(n1701), .ZN(n2107)
         );
  INV_X1 U1877 ( .A(b[12]), .ZN(n1701) );
  INV_X1 U1878 ( .A(n1384), .ZN(n1700) );
  AOI222_X1 U1879 ( .A1(n2108), .A2(n2109), .B1(n2108), .B2(n638), .C1(n638), 
        .C2(n2109), .ZN(n2103) );
  XNOR2_X1 U1880 ( .A(a[2]), .B(n2110), .ZN(n2109) );
  AOI221_X1 U1881 ( .B1(b[13]), .B2(n1561), .C1(b[12]), .C2(n1562), .A(n2111), 
        .ZN(n2110) );
  OAI22_X1 U1882 ( .A1(n1564), .A2(n1696), .B1(n1639), .B2(n1697), .ZN(n2111)
         );
  INV_X1 U1883 ( .A(b[11]), .ZN(n1697) );
  INV_X1 U1884 ( .A(n1385), .ZN(n1696) );
  OAI222_X1 U1885 ( .A1(n2112), .A2(n2113), .B1(n2112), .B2(n2114), .C1(n2114), 
        .C2(n2113), .ZN(n2108) );
  INV_X1 U1886 ( .A(n646), .ZN(n2114) );
  XNOR2_X1 U1887 ( .A(n1742), .B(n2115), .ZN(n2113) );
  AOI221_X1 U1888 ( .B1(b[12]), .B2(n1561), .C1(b[11]), .C2(n1562), .A(n2116), 
        .ZN(n2115) );
  OAI22_X1 U1889 ( .A1(n1564), .A2(n1692), .B1(n1639), .B2(n1693), .ZN(n2116)
         );
  INV_X1 U1890 ( .A(b[10]), .ZN(n1693) );
  INV_X1 U1891 ( .A(n1386), .ZN(n1692) );
  AOI222_X1 U1892 ( .A1(n2117), .A2(n2118), .B1(n2117), .B2(n654), .C1(n654), 
        .C2(n2118), .ZN(n2112) );
  XNOR2_X1 U1893 ( .A(a[2]), .B(n2119), .ZN(n2118) );
  AOI221_X1 U1894 ( .B1(b[11]), .B2(n1561), .C1(b[10]), .C2(n1562), .A(n2120), 
        .ZN(n2119) );
  OAI22_X1 U1895 ( .A1(n1564), .A2(n1688), .B1(n1639), .B2(n1689), .ZN(n2120)
         );
  INV_X1 U1896 ( .A(b[9]), .ZN(n1689) );
  INV_X1 U1897 ( .A(n1387), .ZN(n1688) );
  OAI222_X1 U1898 ( .A1(n2121), .A2(n2122), .B1(n2121), .B2(n2123), .C1(n2123), 
        .C2(n2122), .ZN(n2117) );
  INV_X1 U1899 ( .A(n660), .ZN(n2123) );
  XNOR2_X1 U1900 ( .A(n1742), .B(n2124), .ZN(n2122) );
  AOI221_X1 U1901 ( .B1(b[10]), .B2(n1561), .C1(b[9]), .C2(n1563), .A(n2125), 
        .ZN(n2124) );
  OAI22_X1 U1902 ( .A1(n1564), .A2(n1684), .B1(n1639), .B2(n1685), .ZN(n2125)
         );
  INV_X1 U1903 ( .A(b[8]), .ZN(n1685) );
  INV_X1 U1904 ( .A(n1388), .ZN(n1684) );
  AOI222_X1 U1905 ( .A1(n2126), .A2(n2127), .B1(n2126), .B2(n666), .C1(n666), 
        .C2(n2127), .ZN(n2121) );
  XNOR2_X1 U1906 ( .A(a[2]), .B(n2128), .ZN(n2127) );
  AOI221_X1 U1907 ( .B1(b[9]), .B2(n1561), .C1(b[8]), .C2(n1563), .A(n2129), 
        .ZN(n2128) );
  OAI22_X1 U1908 ( .A1(n1564), .A2(n1680), .B1(n1639), .B2(n1681), .ZN(n2129)
         );
  INV_X1 U1909 ( .A(b[7]), .ZN(n1681) );
  INV_X1 U1910 ( .A(n1389), .ZN(n1680) );
  OAI222_X1 U1911 ( .A1(n2130), .A2(n2131), .B1(n2130), .B2(n2132), .C1(n2132), 
        .C2(n2131), .ZN(n2126) );
  INV_X1 U1912 ( .A(n672), .ZN(n2132) );
  XNOR2_X1 U1913 ( .A(n1742), .B(n2133), .ZN(n2131) );
  AOI221_X1 U1914 ( .B1(b[8]), .B2(n1561), .C1(b[7]), .C2(n1562), .A(n2134), 
        .ZN(n2133) );
  OAI22_X1 U1915 ( .A1(n1564), .A2(n1676), .B1(n1639), .B2(n1677), .ZN(n2134)
         );
  INV_X1 U1916 ( .A(b[6]), .ZN(n1677) );
  INV_X1 U1917 ( .A(n1390), .ZN(n1676) );
  AOI222_X1 U1918 ( .A1(n2135), .A2(n2136), .B1(n2135), .B2(n676), .C1(n676), 
        .C2(n2136), .ZN(n2130) );
  XNOR2_X1 U1919 ( .A(a[2]), .B(n2137), .ZN(n2136) );
  AOI221_X1 U1920 ( .B1(b[7]), .B2(n1561), .C1(b[6]), .C2(n1563), .A(n2138), 
        .ZN(n2137) );
  OAI22_X1 U1921 ( .A1(n1564), .A2(n1672), .B1(n1639), .B2(n1673), .ZN(n2138)
         );
  INV_X1 U1922 ( .A(b[5]), .ZN(n1673) );
  INV_X1 U1923 ( .A(n1391), .ZN(n1672) );
  OAI222_X1 U1924 ( .A1(n2139), .A2(n2140), .B1(n2139), .B2(n2141), .C1(n2141), 
        .C2(n2140), .ZN(n2135) );
  INV_X1 U1925 ( .A(n680), .ZN(n2141) );
  XNOR2_X1 U1926 ( .A(n1742), .B(n2142), .ZN(n2140) );
  AOI221_X1 U1927 ( .B1(b[6]), .B2(n1561), .C1(b[5]), .C2(n1563), .A(n2143), 
        .ZN(n2142) );
  OAI22_X1 U1928 ( .A1(n1564), .A2(n1668), .B1(n1639), .B2(n1669), .ZN(n2143)
         );
  INV_X1 U1929 ( .A(b[4]), .ZN(n1669) );
  INV_X1 U1930 ( .A(n1392), .ZN(n1668) );
  AOI222_X1 U1931 ( .A1(n2144), .A2(n2145), .B1(n2144), .B2(n684), .C1(n684), 
        .C2(n2145), .ZN(n2139) );
  XNOR2_X1 U1932 ( .A(a[2]), .B(n2146), .ZN(n2145) );
  AOI221_X1 U1933 ( .B1(b[5]), .B2(n1561), .C1(b[4]), .C2(n1563), .A(n2147), 
        .ZN(n2146) );
  OAI22_X1 U1934 ( .A1(n1564), .A2(n1664), .B1(n1639), .B2(n1665), .ZN(n2147)
         );
  INV_X1 U1935 ( .A(b[3]), .ZN(n1665) );
  INV_X1 U1936 ( .A(n1393), .ZN(n1664) );
  OAI222_X1 U1937 ( .A1(n2148), .A2(n2149), .B1(n2148), .B2(n2150), .C1(n2150), 
        .C2(n2149), .ZN(n2144) );
  INV_X1 U1938 ( .A(n686), .ZN(n2150) );
  XNOR2_X1 U1939 ( .A(n1742), .B(n2151), .ZN(n2149) );
  AOI221_X1 U1940 ( .B1(b[4]), .B2(n1561), .C1(b[3]), .C2(n1563), .A(n2152), 
        .ZN(n2151) );
  OAI22_X1 U1941 ( .A1(n1564), .A2(n1660), .B1(n1639), .B2(n1661), .ZN(n2152)
         );
  INV_X1 U1942 ( .A(n1394), .ZN(n1660) );
  AOI222_X1 U1943 ( .A1(n2153), .A2(n2154), .B1(n2153), .B2(n688), .C1(n688), 
        .C2(n2154), .ZN(n2148) );
  XNOR2_X1 U1944 ( .A(a[2]), .B(n2155), .ZN(n2154) );
  AOI221_X1 U1945 ( .B1(b[3]), .B2(n1561), .C1(b[2]), .C2(n1563), .A(n2156), 
        .ZN(n2155) );
  OAI22_X1 U1946 ( .A1(n1564), .A2(n1657), .B1(n1639), .B2(n1649), .ZN(n2156)
         );
  INV_X1 U1947 ( .A(b[1]), .ZN(n1649) );
  INV_X1 U1948 ( .A(n1395), .ZN(n1657) );
  AND2_X1 U1949 ( .A1(n2160), .A2(n2161), .ZN(n2153) );
  AOI211_X1 U1950 ( .C1(b[1]), .C2(n1561), .A(n2162), .B(b[0]), .ZN(n2161) );
  OAI22_X1 U1951 ( .A1(n1535), .A2(n1661), .B1(n1564), .B2(n1650), .ZN(n2162)
         );
  INV_X1 U1952 ( .A(n1397), .ZN(n1650) );
  INV_X1 U1953 ( .A(b[2]), .ZN(n1661) );
  INV_X1 U1954 ( .A(a[0]), .ZN(n2158) );
  AOI221_X1 U1955 ( .B1(b[1]), .B2(n1563), .C1(n1396), .C2(n1555), .A(n1742), 
        .ZN(n2160) );
  XNOR2_X1 U1956 ( .A(a[1]), .B(n1742), .ZN(n2157) );
  INV_X1 U1957 ( .A(a[2]), .ZN(n1742) );
  NOR2_X1 U1958 ( .A1(n2159), .A2(a[0]), .ZN(n1636) );
  INV_X1 U1959 ( .A(a[1]), .ZN(n2159) );
endmodule


module iir_filter_DW_mult_tc_2 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(product[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(product[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(product[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(product[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(product[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(product[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(product[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(product[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(product[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(product[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(product[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(product[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(product[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(product[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(product[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(product[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(product[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(product[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(product[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(product[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(product[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(product[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(product[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1598), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1600), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1602), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1604), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1606), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1608), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1610), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(b[22]), .B(n1614), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(b[21]), .B(b[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(b[20]), .B(b[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(b[19]), .B(b[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(b[18]), .B(b[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(b[17]), .B(b[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(b[16]), .B(b[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(b[15]), .B(b[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(b[14]), .B(b[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(b[13]), .B(b[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(b[12]), .B(b[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(b[11]), .B(b[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(b[10]), .B(b[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(b[9]), .B(b[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(b[8]), .B(b[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(b[7]), .B(b[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(b[6]), .B(b[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(b[5]), .B(b[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(b[4]), .B(b[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(b[3]), .B(b[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(b[2]), .B(b[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(b[1]), .B(b[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(b[0]), .B(b[1]), .CO(n727), .S(n1397) );
  INV_X1 U1137 ( .A(n1533), .ZN(n1570) );
  INV_X1 U1138 ( .A(n1536), .ZN(n1568) );
  INV_X1 U1139 ( .A(n1535), .ZN(n1561) );
  INV_X1 U1140 ( .A(n1534), .ZN(n1569) );
  BUF_X1 U1141 ( .A(n1654), .Z(n1572) );
  INV_X1 U1142 ( .A(n1547), .ZN(n1560) );
  INV_X1 U1143 ( .A(n1544), .ZN(n1558) );
  INV_X1 U1144 ( .A(n1537), .ZN(n1580) );
  INV_X1 U1145 ( .A(n1551), .ZN(n1575) );
  INV_X1 U1146 ( .A(n1550), .ZN(n1585) );
  INV_X1 U1147 ( .A(n1548), .ZN(n1595) );
  INV_X1 U1148 ( .A(n1549), .ZN(n1590) );
  INV_X1 U1149 ( .A(n1538), .ZN(n1559) );
  INV_X1 U1150 ( .A(n1545), .ZN(n1593) );
  INV_X1 U1151 ( .A(n1553), .ZN(n1583) );
  INV_X1 U1152 ( .A(n1552), .ZN(n1588) );
  INV_X1 U1153 ( .A(n1546), .ZN(n1578) );
  INV_X1 U1154 ( .A(n1554), .ZN(n1573) );
  BUF_X1 U1155 ( .A(n1654), .Z(n1571) );
  BUF_X1 U1156 ( .A(n1629), .Z(n1557) );
  BUF_X1 U1157 ( .A(n1967), .Z(n1596) );
  BUF_X1 U1158 ( .A(n1912), .Z(n1591) );
  BUF_X1 U1159 ( .A(n1857), .Z(n1586) );
  BUF_X1 U1160 ( .A(n1802), .Z(n1581) );
  BUF_X1 U1161 ( .A(n1747), .Z(n1576) );
  BUF_X1 U1162 ( .A(n1912), .Z(n1592) );
  BUF_X1 U1163 ( .A(n1857), .Z(n1587) );
  BUF_X1 U1164 ( .A(n1802), .Z(n1582) );
  BUF_X1 U1165 ( .A(n1747), .Z(n1577) );
  BUF_X1 U1166 ( .A(n1967), .Z(n1597) );
  INV_X1 U1167 ( .A(n1615), .ZN(n1614) );
  INV_X1 U1168 ( .A(n1540), .ZN(n1589) );
  INV_X1 U1169 ( .A(n1541), .ZN(n1584) );
  INV_X1 U1170 ( .A(n1542), .ZN(n1579) );
  INV_X1 U1171 ( .A(n1543), .ZN(n1574) );
  BUF_X1 U1172 ( .A(n1629), .Z(n1556) );
  INV_X1 U1173 ( .A(n1539), .ZN(n1594) );
  NAND3_X1 U1174 ( .A1(n2157), .A2(n2158), .A3(n2159), .ZN(n1639) );
  INV_X1 U1175 ( .A(n1555), .ZN(n1564) );
  OR2_X1 U1176 ( .A1(n1738), .A2(n1739), .ZN(n1533) );
  OR2_X1 U1177 ( .A1(n1740), .A2(n1741), .ZN(n1534) );
  OR2_X1 U1178 ( .A1(n2158), .A2(n2157), .ZN(n1535) );
  AND2_X1 U1179 ( .A1(n1738), .A2(n1740), .ZN(n1536) );
  INV_X1 U1180 ( .A(n1611), .ZN(n1610) );
  INV_X1 U1181 ( .A(n1607), .ZN(n1606) );
  INV_X1 U1182 ( .A(n1609), .ZN(n1608) );
  INV_X1 U1183 ( .A(n1603), .ZN(n1602) );
  INV_X1 U1184 ( .A(n1605), .ZN(n1604) );
  OR2_X1 U1185 ( .A1(n1849), .A2(n1850), .ZN(n1537) );
  BUF_X1 U1186 ( .A(n1636), .Z(n1562) );
  BUF_X1 U1187 ( .A(n1636), .Z(n1563) );
  BUF_X1 U1188 ( .A(n1647), .Z(n1565) );
  BUF_X1 U1189 ( .A(n1647), .Z(n1566) );
  OR2_X1 U1190 ( .A1(n2068), .A2(n2067), .ZN(n1538) );
  OR2_X1 U1191 ( .A1(n2016), .A2(n2017), .ZN(n1539) );
  OR2_X1 U1192 ( .A1(n1961), .A2(n1962), .ZN(n1540) );
  OR2_X1 U1193 ( .A1(n1906), .A2(n1907), .ZN(n1541) );
  OR2_X1 U1194 ( .A1(n1851), .A2(n1852), .ZN(n1542) );
  OR2_X1 U1195 ( .A1(n1796), .A2(n1797), .ZN(n1543) );
  AND2_X1 U1196 ( .A1(n2070), .A2(n2068), .ZN(n1544) );
  AND2_X1 U1197 ( .A1(n2014), .A2(n2016), .ZN(n1545) );
  AND2_X1 U1198 ( .A1(n1849), .A2(n1851), .ZN(n1546) );
  OR2_X1 U1199 ( .A1(n2070), .A2(n2069), .ZN(n1547) );
  OR2_X1 U1200 ( .A1(n2014), .A2(n2015), .ZN(n1548) );
  OR2_X1 U1201 ( .A1(n1959), .A2(n1960), .ZN(n1549) );
  OR2_X1 U1202 ( .A1(n1904), .A2(n1905), .ZN(n1550) );
  OR2_X1 U1203 ( .A1(n1794), .A2(n1795), .ZN(n1551) );
  AND2_X1 U1204 ( .A1(n1959), .A2(n1961), .ZN(n1552) );
  AND2_X1 U1205 ( .A1(n1904), .A2(n1906), .ZN(n1553) );
  AND2_X1 U1206 ( .A1(n1794), .A2(n1796), .ZN(n1554) );
  BUF_X1 U1207 ( .A(n1647), .Z(n1567) );
  INV_X1 U1208 ( .A(n1599), .ZN(n1598) );
  AND2_X1 U1209 ( .A1(a[0]), .A2(n2157), .ZN(n1555) );
  BUF_X1 U1210 ( .A(a[20]), .Z(n1600) );
  INV_X1 U1211 ( .A(a[23]), .ZN(n1599) );
  INV_X1 U1212 ( .A(a[5]), .ZN(n1611) );
  INV_X1 U1213 ( .A(a[11]), .ZN(n1607) );
  INV_X1 U1214 ( .A(a[8]), .ZN(n1609) );
  INV_X1 U1215 ( .A(a[17]), .ZN(n1603) );
  INV_X1 U1216 ( .A(a[14]), .ZN(n1605) );
  BUF_X1 U1217 ( .A(a[20]), .Z(n1601) );
  CLKBUF_X1 U1218 ( .A(b[23]), .Z(n1612) );
  CLKBUF_X1 U1219 ( .A(b[23]), .Z(n1613) );
  INV_X1 U1220 ( .A(b[23]), .ZN(n1615) );
  INV_X1 U1221 ( .A(n1612), .ZN(n1616) );
  INV_X1 U1222 ( .A(n1612), .ZN(n1617) );
  INV_X1 U1223 ( .A(n1612), .ZN(n1618) );
  INV_X1 U1224 ( .A(n1613), .ZN(n1619) );
  INV_X1 U1225 ( .A(n1613), .ZN(n1620) );
  AOI21_X1 U1226 ( .B1(n1621), .B2(n1622), .A(n1623), .ZN(product[47]) );
  OAI22_X1 U1227 ( .A1(n1624), .A2(n1625), .B1(n1624), .B2(n1626), .ZN(n1623)
         );
  INV_X1 U1228 ( .A(n1622), .ZN(n1626) );
  AOI222_X1 U1229 ( .A1(n1627), .A2(n303), .B1(n1625), .B2(n303), .C1(n1627), 
        .C2(n1625), .ZN(n1624) );
  XOR2_X1 U1230 ( .A(n1628), .B(n1599), .Z(n1622) );
  OAI221_X1 U1231 ( .B1(n1617), .B2(n1557), .C1(n1620), .C2(n1558), .A(n1630), 
        .ZN(n1628) );
  OAI21_X1 U1232 ( .B1(n1559), .B2(n1560), .A(n1614), .ZN(n1630) );
  INV_X1 U1233 ( .A(n1625), .ZN(n1621) );
  XOR2_X1 U1234 ( .A(a[23]), .B(n1631), .Z(n1625) );
  AOI221_X1 U1235 ( .B1(n1613), .B2(n1559), .C1(n1560), .C2(n1614), .A(n1632), 
        .ZN(n1631) );
  OAI22_X1 U1236 ( .A1(n1558), .A2(n1633), .B1(n1557), .B2(n1634), .ZN(n1632)
         );
  XNOR2_X1 U1237 ( .A(a[2]), .B(n1635), .ZN(n908) );
  AOI221_X1 U1238 ( .B1(n1561), .B2(b[22]), .C1(n1563), .C2(b[21]), .A(n1637), 
        .ZN(n1635) );
  OAI22_X1 U1239 ( .A1(n1564), .A2(n1638), .B1(n1639), .B2(n1640), .ZN(n1637)
         );
  INV_X1 U1240 ( .A(n1376), .ZN(n1638) );
  XNOR2_X1 U1241 ( .A(a[2]), .B(n1641), .ZN(n907) );
  AOI221_X1 U1242 ( .B1(n1563), .B2(b[22]), .C1(n1555), .C2(n1375), .A(n1642), 
        .ZN(n1641) );
  OAI22_X1 U1243 ( .A1(n1643), .A2(n1639), .B1(n1617), .B2(n1535), .ZN(n1642)
         );
  XNOR2_X1 U1244 ( .A(a[2]), .B(n1644), .ZN(n906) );
  AOI221_X1 U1245 ( .B1(n1561), .B2(n1613), .C1(n1563), .C2(n1614), .A(n1645), 
        .ZN(n1644) );
  OAI22_X1 U1246 ( .A1(n1633), .A2(n1564), .B1(n1634), .B2(n1639), .ZN(n1645)
         );
  XNOR2_X1 U1247 ( .A(n1646), .B(n1611), .ZN(n904) );
  OAI22_X1 U1248 ( .A1(n1565), .A2(n1534), .B1(n1568), .B2(n1567), .ZN(n1646)
         );
  XNOR2_X1 U1249 ( .A(n1648), .B(n1611), .ZN(n903) );
  OAI222_X1 U1250 ( .A1(n1534), .A2(n1649), .B1(n1566), .B2(n1533), .C1(n1568), 
        .C2(n1650), .ZN(n1648) );
  XNOR2_X1 U1251 ( .A(n1610), .B(n1651), .ZN(n902) );
  AOI221_X1 U1252 ( .B1(b[2]), .B2(n1569), .C1(b[1]), .C2(n1570), .A(n1652), 
        .ZN(n1651) );
  OAI22_X1 U1253 ( .A1(n1568), .A2(n1653), .B1(n1565), .B2(n1572), .ZN(n1652)
         );
  XNOR2_X1 U1254 ( .A(n1610), .B(n1655), .ZN(n901) );
  AOI221_X1 U1255 ( .B1(b[3]), .B2(n1569), .C1(b[2]), .C2(n1570), .A(n1656), 
        .ZN(n1655) );
  OAI22_X1 U1256 ( .A1(n1568), .A2(n1657), .B1(n1649), .B2(n1572), .ZN(n1656)
         );
  XNOR2_X1 U1257 ( .A(n1610), .B(n1658), .ZN(n900) );
  AOI221_X1 U1258 ( .B1(b[4]), .B2(n1569), .C1(b[3]), .C2(n1570), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1259 ( .A1(n1568), .A2(n1660), .B1(n1661), .B2(n1572), .ZN(n1659)
         );
  XNOR2_X1 U1260 ( .A(n1610), .B(n1662), .ZN(n899) );
  AOI221_X1 U1261 ( .B1(b[5]), .B2(n1569), .C1(b[4]), .C2(n1570), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1262 ( .A1(n1568), .A2(n1664), .B1(n1572), .B2(n1665), .ZN(n1663)
         );
  XNOR2_X1 U1263 ( .A(n1610), .B(n1666), .ZN(n898) );
  AOI221_X1 U1264 ( .B1(b[6]), .B2(n1569), .C1(b[5]), .C2(n1570), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1265 ( .A1(n1568), .A2(n1668), .B1(n1572), .B2(n1669), .ZN(n1667)
         );
  XNOR2_X1 U1266 ( .A(n1610), .B(n1670), .ZN(n897) );
  AOI221_X1 U1267 ( .B1(b[7]), .B2(n1569), .C1(b[6]), .C2(n1570), .A(n1671), 
        .ZN(n1670) );
  OAI22_X1 U1268 ( .A1(n1568), .A2(n1672), .B1(n1572), .B2(n1673), .ZN(n1671)
         );
  XNOR2_X1 U1269 ( .A(n1610), .B(n1674), .ZN(n896) );
  AOI221_X1 U1270 ( .B1(b[8]), .B2(n1569), .C1(b[7]), .C2(n1570), .A(n1675), 
        .ZN(n1674) );
  OAI22_X1 U1271 ( .A1(n1568), .A2(n1676), .B1(n1571), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1272 ( .A(n1610), .B(n1678), .ZN(n895) );
  AOI221_X1 U1273 ( .B1(b[9]), .B2(n1569), .C1(b[8]), .C2(n1570), .A(n1679), 
        .ZN(n1678) );
  OAI22_X1 U1274 ( .A1(n1568), .A2(n1680), .B1(n1572), .B2(n1681), .ZN(n1679)
         );
  XNOR2_X1 U1275 ( .A(n1610), .B(n1682), .ZN(n894) );
  AOI221_X1 U1276 ( .B1(b[10]), .B2(n1569), .C1(b[9]), .C2(n1570), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1277 ( .A1(n1568), .A2(n1684), .B1(n1572), .B2(n1685), .ZN(n1683)
         );
  XNOR2_X1 U1278 ( .A(n1610), .B(n1686), .ZN(n893) );
  AOI221_X1 U1279 ( .B1(b[11]), .B2(n1569), .C1(b[10]), .C2(n1570), .A(n1687), 
        .ZN(n1686) );
  OAI22_X1 U1280 ( .A1(n1568), .A2(n1688), .B1(n1571), .B2(n1689), .ZN(n1687)
         );
  XNOR2_X1 U1281 ( .A(n1610), .B(n1690), .ZN(n892) );
  AOI221_X1 U1282 ( .B1(b[12]), .B2(n1569), .C1(b[11]), .C2(n1570), .A(n1691), 
        .ZN(n1690) );
  OAI22_X1 U1283 ( .A1(n1568), .A2(n1692), .B1(n1571), .B2(n1693), .ZN(n1691)
         );
  XNOR2_X1 U1284 ( .A(n1610), .B(n1694), .ZN(n891) );
  AOI221_X1 U1285 ( .B1(b[13]), .B2(n1569), .C1(b[12]), .C2(n1570), .A(n1695), 
        .ZN(n1694) );
  OAI22_X1 U1286 ( .A1(n1568), .A2(n1696), .B1(n1571), .B2(n1697), .ZN(n1695)
         );
  XNOR2_X1 U1287 ( .A(n1610), .B(n1698), .ZN(n890) );
  AOI221_X1 U1288 ( .B1(b[14]), .B2(n1569), .C1(b[13]), .C2(n1570), .A(n1699), 
        .ZN(n1698) );
  OAI22_X1 U1289 ( .A1(n1568), .A2(n1700), .B1(n1571), .B2(n1701), .ZN(n1699)
         );
  XNOR2_X1 U1290 ( .A(n1610), .B(n1702), .ZN(n889) );
  AOI221_X1 U1291 ( .B1(b[15]), .B2(n1569), .C1(b[14]), .C2(n1570), .A(n1703), 
        .ZN(n1702) );
  OAI22_X1 U1292 ( .A1(n1568), .A2(n1704), .B1(n1571), .B2(n1705), .ZN(n1703)
         );
  XNOR2_X1 U1293 ( .A(n1610), .B(n1706), .ZN(n888) );
  AOI221_X1 U1294 ( .B1(b[16]), .B2(n1569), .C1(b[15]), .C2(n1570), .A(n1707), 
        .ZN(n1706) );
  OAI22_X1 U1295 ( .A1(n1568), .A2(n1708), .B1(n1571), .B2(n1709), .ZN(n1707)
         );
  XNOR2_X1 U1296 ( .A(n1610), .B(n1710), .ZN(n887) );
  AOI221_X1 U1297 ( .B1(b[17]), .B2(n1569), .C1(b[16]), .C2(n1570), .A(n1711), 
        .ZN(n1710) );
  OAI22_X1 U1298 ( .A1(n1568), .A2(n1712), .B1(n1571), .B2(n1713), .ZN(n1711)
         );
  XNOR2_X1 U1299 ( .A(n1610), .B(n1714), .ZN(n886) );
  AOI221_X1 U1300 ( .B1(b[18]), .B2(n1569), .C1(b[17]), .C2(n1570), .A(n1715), 
        .ZN(n1714) );
  OAI22_X1 U1301 ( .A1(n1568), .A2(n1716), .B1(n1571), .B2(n1717), .ZN(n1715)
         );
  XNOR2_X1 U1302 ( .A(n1610), .B(n1718), .ZN(n885) );
  AOI221_X1 U1303 ( .B1(b[19]), .B2(n1569), .C1(b[18]), .C2(n1570), .A(n1719), 
        .ZN(n1718) );
  OAI22_X1 U1304 ( .A1(n1568), .A2(n1720), .B1(n1571), .B2(n1721), .ZN(n1719)
         );
  XNOR2_X1 U1305 ( .A(a[5]), .B(n1722), .ZN(n884) );
  AOI221_X1 U1306 ( .B1(n1569), .B2(b[20]), .C1(b[19]), .C2(n1570), .A(n1723), 
        .ZN(n1722) );
  OAI22_X1 U1307 ( .A1(n1568), .A2(n1724), .B1(n1571), .B2(n1725), .ZN(n1723)
         );
  XNOR2_X1 U1308 ( .A(a[5]), .B(n1726), .ZN(n883) );
  AOI221_X1 U1309 ( .B1(n1569), .B2(b[21]), .C1(n1570), .C2(b[20]), .A(n1727), 
        .ZN(n1726) );
  OAI22_X1 U1310 ( .A1(n1568), .A2(n1728), .B1(n1571), .B2(n1729), .ZN(n1727)
         );
  XNOR2_X1 U1311 ( .A(a[5]), .B(n1730), .ZN(n882) );
  AOI221_X1 U1312 ( .B1(n1569), .B2(b[22]), .C1(n1536), .C2(n1376), .A(n1731), 
        .ZN(n1730) );
  OAI22_X1 U1313 ( .A1(n1640), .A2(n1572), .B1(n1643), .B2(n1533), .ZN(n1731)
         );
  XNOR2_X1 U1314 ( .A(a[5]), .B(n1732), .ZN(n881) );
  AOI221_X1 U1315 ( .B1(n1570), .B2(b[22]), .C1(n1536), .C2(n1375), .A(n1733), 
        .ZN(n1732) );
  OAI22_X1 U1316 ( .A1(n1615), .A2(n1534), .B1(n1643), .B2(n1572), .ZN(n1733)
         );
  XNOR2_X1 U1317 ( .A(a[5]), .B(n1734), .ZN(n880) );
  AOI221_X1 U1318 ( .B1(n1569), .B2(n1613), .C1(n1570), .C2(n1614), .A(n1735), 
        .ZN(n1734) );
  OAI22_X1 U1319 ( .A1(n1633), .A2(n1568), .B1(n1634), .B2(n1572), .ZN(n1735)
         );
  XNOR2_X1 U1320 ( .A(n1610), .B(n1736), .ZN(n879) );
  OAI221_X1 U1321 ( .B1(n1616), .B2(n1572), .C1(n1620), .C2(n1568), .A(n1737), 
        .ZN(n1736) );
  OAI21_X1 U1322 ( .B1(n1569), .B2(n1570), .A(n1614), .ZN(n1737) );
  INV_X1 U1323 ( .A(n1741), .ZN(n1738) );
  NAND3_X1 U1324 ( .A1(n1741), .A2(n1740), .A3(n1739), .ZN(n1654) );
  XNOR2_X1 U1325 ( .A(a[3]), .B(a[4]), .ZN(n1739) );
  XNOR2_X1 U1326 ( .A(a[4]), .B(n1611), .ZN(n1740) );
  XOR2_X1 U1327 ( .A(a[3]), .B(n1742), .Z(n1741) );
  XNOR2_X1 U1328 ( .A(n1743), .B(n1609), .ZN(n878) );
  OAI22_X1 U1329 ( .A1(n1565), .A2(n1543), .B1(n1565), .B2(n1573), .ZN(n1743)
         );
  XNOR2_X1 U1330 ( .A(n1744), .B(n1609), .ZN(n877) );
  OAI222_X1 U1331 ( .A1(n1649), .A2(n1543), .B1(n1566), .B2(n1551), .C1(n1650), 
        .C2(n1573), .ZN(n1744) );
  XNOR2_X1 U1332 ( .A(n1608), .B(n1745), .ZN(n876) );
  AOI221_X1 U1333 ( .B1(n1574), .B2(b[2]), .C1(n1575), .C2(b[1]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1334 ( .A1(n1653), .A2(n1573), .B1(n1565), .B2(n1576), .ZN(n1746)
         );
  XNOR2_X1 U1335 ( .A(n1608), .B(n1748), .ZN(n875) );
  AOI221_X1 U1336 ( .B1(n1574), .B2(b[3]), .C1(n1575), .C2(b[2]), .A(n1749), 
        .ZN(n1748) );
  OAI22_X1 U1337 ( .A1(n1657), .A2(n1573), .B1(n1649), .B2(n1577), .ZN(n1749)
         );
  XNOR2_X1 U1338 ( .A(n1608), .B(n1750), .ZN(n874) );
  AOI221_X1 U1339 ( .B1(n1574), .B2(b[4]), .C1(n1575), .C2(b[3]), .A(n1751), 
        .ZN(n1750) );
  OAI22_X1 U1340 ( .A1(n1660), .A2(n1573), .B1(n1661), .B2(n1577), .ZN(n1751)
         );
  XNOR2_X1 U1341 ( .A(n1608), .B(n1752), .ZN(n873) );
  AOI221_X1 U1342 ( .B1(n1574), .B2(b[5]), .C1(n1575), .C2(b[4]), .A(n1753), 
        .ZN(n1752) );
  OAI22_X1 U1343 ( .A1(n1664), .A2(n1573), .B1(n1665), .B2(n1577), .ZN(n1753)
         );
  XNOR2_X1 U1344 ( .A(n1608), .B(n1754), .ZN(n872) );
  AOI221_X1 U1345 ( .B1(n1574), .B2(b[6]), .C1(n1575), .C2(b[5]), .A(n1755), 
        .ZN(n1754) );
  OAI22_X1 U1346 ( .A1(n1668), .A2(n1573), .B1(n1669), .B2(n1577), .ZN(n1755)
         );
  XNOR2_X1 U1347 ( .A(n1608), .B(n1756), .ZN(n871) );
  AOI221_X1 U1348 ( .B1(n1574), .B2(b[7]), .C1(n1575), .C2(b[6]), .A(n1757), 
        .ZN(n1756) );
  OAI22_X1 U1349 ( .A1(n1672), .A2(n1573), .B1(n1673), .B2(n1577), .ZN(n1757)
         );
  XNOR2_X1 U1350 ( .A(n1608), .B(n1758), .ZN(n870) );
  AOI221_X1 U1351 ( .B1(n1574), .B2(b[8]), .C1(n1575), .C2(b[7]), .A(n1759), 
        .ZN(n1758) );
  OAI22_X1 U1352 ( .A1(n1676), .A2(n1573), .B1(n1677), .B2(n1577), .ZN(n1759)
         );
  XNOR2_X1 U1353 ( .A(n1608), .B(n1760), .ZN(n869) );
  AOI221_X1 U1354 ( .B1(n1574), .B2(b[9]), .C1(n1575), .C2(b[8]), .A(n1761), 
        .ZN(n1760) );
  OAI22_X1 U1355 ( .A1(n1680), .A2(n1573), .B1(n1681), .B2(n1577), .ZN(n1761)
         );
  XNOR2_X1 U1356 ( .A(n1608), .B(n1762), .ZN(n868) );
  AOI221_X1 U1357 ( .B1(n1574), .B2(b[10]), .C1(n1575), .C2(b[9]), .A(n1763), 
        .ZN(n1762) );
  OAI22_X1 U1358 ( .A1(n1684), .A2(n1573), .B1(n1685), .B2(n1577), .ZN(n1763)
         );
  XNOR2_X1 U1359 ( .A(n1608), .B(n1764), .ZN(n867) );
  AOI221_X1 U1360 ( .B1(n1574), .B2(b[11]), .C1(n1575), .C2(b[10]), .A(n1765), 
        .ZN(n1764) );
  OAI22_X1 U1361 ( .A1(n1688), .A2(n1573), .B1(n1689), .B2(n1577), .ZN(n1765)
         );
  XNOR2_X1 U1362 ( .A(n1608), .B(n1766), .ZN(n866) );
  AOI221_X1 U1363 ( .B1(n1574), .B2(b[12]), .C1(n1575), .C2(b[11]), .A(n1767), 
        .ZN(n1766) );
  OAI22_X1 U1364 ( .A1(n1692), .A2(n1573), .B1(n1693), .B2(n1577), .ZN(n1767)
         );
  XNOR2_X1 U1365 ( .A(n1608), .B(n1768), .ZN(n865) );
  AOI221_X1 U1366 ( .B1(n1574), .B2(b[13]), .C1(n1575), .C2(b[12]), .A(n1769), 
        .ZN(n1768) );
  OAI22_X1 U1367 ( .A1(n1696), .A2(n1573), .B1(n1697), .B2(n1576), .ZN(n1769)
         );
  XNOR2_X1 U1368 ( .A(n1608), .B(n1770), .ZN(n864) );
  AOI221_X1 U1369 ( .B1(n1574), .B2(b[14]), .C1(n1575), .C2(b[13]), .A(n1771), 
        .ZN(n1770) );
  OAI22_X1 U1370 ( .A1(n1700), .A2(n1573), .B1(n1701), .B2(n1576), .ZN(n1771)
         );
  XNOR2_X1 U1371 ( .A(n1608), .B(n1772), .ZN(n863) );
  AOI221_X1 U1372 ( .B1(n1574), .B2(b[15]), .C1(n1575), .C2(b[14]), .A(n1773), 
        .ZN(n1772) );
  OAI22_X1 U1373 ( .A1(n1704), .A2(n1573), .B1(n1705), .B2(n1576), .ZN(n1773)
         );
  XNOR2_X1 U1374 ( .A(n1608), .B(n1774), .ZN(n862) );
  AOI221_X1 U1375 ( .B1(n1574), .B2(b[16]), .C1(n1575), .C2(b[15]), .A(n1775), 
        .ZN(n1774) );
  OAI22_X1 U1376 ( .A1(n1708), .A2(n1573), .B1(n1709), .B2(n1576), .ZN(n1775)
         );
  XNOR2_X1 U1377 ( .A(n1608), .B(n1776), .ZN(n861) );
  AOI221_X1 U1378 ( .B1(n1574), .B2(b[17]), .C1(n1575), .C2(b[16]), .A(n1777), 
        .ZN(n1776) );
  OAI22_X1 U1379 ( .A1(n1712), .A2(n1573), .B1(n1713), .B2(n1576), .ZN(n1777)
         );
  XNOR2_X1 U1380 ( .A(n1608), .B(n1778), .ZN(n860) );
  AOI221_X1 U1381 ( .B1(n1574), .B2(b[18]), .C1(n1575), .C2(b[17]), .A(n1779), 
        .ZN(n1778) );
  OAI22_X1 U1382 ( .A1(n1716), .A2(n1573), .B1(n1717), .B2(n1576), .ZN(n1779)
         );
  XNOR2_X1 U1383 ( .A(n1608), .B(n1780), .ZN(n859) );
  AOI221_X1 U1384 ( .B1(n1574), .B2(b[19]), .C1(n1575), .C2(b[18]), .A(n1781), 
        .ZN(n1780) );
  OAI22_X1 U1385 ( .A1(n1720), .A2(n1573), .B1(n1721), .B2(n1576), .ZN(n1781)
         );
  XNOR2_X1 U1386 ( .A(a[8]), .B(n1782), .ZN(n858) );
  AOI221_X1 U1387 ( .B1(n1574), .B2(b[20]), .C1(n1575), .C2(b[19]), .A(n1783), 
        .ZN(n1782) );
  OAI22_X1 U1388 ( .A1(n1724), .A2(n1573), .B1(n1725), .B2(n1576), .ZN(n1783)
         );
  XNOR2_X1 U1389 ( .A(a[8]), .B(n1784), .ZN(n857) );
  AOI221_X1 U1390 ( .B1(n1574), .B2(b[21]), .C1(n1575), .C2(b[20]), .A(n1785), 
        .ZN(n1784) );
  OAI22_X1 U1391 ( .A1(n1728), .A2(n1573), .B1(n1729), .B2(n1576), .ZN(n1785)
         );
  XNOR2_X1 U1392 ( .A(a[8]), .B(n1786), .ZN(n856) );
  AOI221_X1 U1393 ( .B1(n1574), .B2(b[22]), .C1(n1554), .C2(n1376), .A(n1787), 
        .ZN(n1786) );
  OAI22_X1 U1394 ( .A1(n1640), .A2(n1577), .B1(n1643), .B2(n1551), .ZN(n1787)
         );
  XNOR2_X1 U1395 ( .A(a[8]), .B(n1788), .ZN(n855) );
  AOI221_X1 U1396 ( .B1(n1575), .B2(b[22]), .C1(n1554), .C2(n1375), .A(n1789), 
        .ZN(n1788) );
  OAI22_X1 U1397 ( .A1(n1617), .A2(n1543), .B1(n1643), .B2(n1576), .ZN(n1789)
         );
  XNOR2_X1 U1398 ( .A(a[8]), .B(n1790), .ZN(n854) );
  AOI221_X1 U1399 ( .B1(n1574), .B2(n1613), .C1(n1575), .C2(n1614), .A(n1791), 
        .ZN(n1790) );
  OAI22_X1 U1400 ( .A1(n1633), .A2(n1573), .B1(n1634), .B2(n1576), .ZN(n1791)
         );
  XNOR2_X1 U1401 ( .A(n1608), .B(n1792), .ZN(n853) );
  OAI221_X1 U1402 ( .B1(n1616), .B2(n1577), .C1(n1617), .C2(n1573), .A(n1793), 
        .ZN(n1792) );
  OAI21_X1 U1403 ( .B1(n1574), .B2(n1575), .A(n1614), .ZN(n1793) );
  INV_X1 U1404 ( .A(n1797), .ZN(n1794) );
  NAND3_X1 U1405 ( .A1(n1797), .A2(n1796), .A3(n1795), .ZN(n1747) );
  XNOR2_X1 U1406 ( .A(a[6]), .B(a[7]), .ZN(n1795) );
  XNOR2_X1 U1407 ( .A(a[7]), .B(n1609), .ZN(n1796) );
  XOR2_X1 U1408 ( .A(a[6]), .B(n1611), .Z(n1797) );
  XNOR2_X1 U1409 ( .A(n1798), .B(n1607), .ZN(n852) );
  OAI22_X1 U1410 ( .A1(n1565), .A2(n1542), .B1(n1565), .B2(n1578), .ZN(n1798)
         );
  XNOR2_X1 U1411 ( .A(n1799), .B(n1607), .ZN(n851) );
  OAI222_X1 U1412 ( .A1(n1649), .A2(n1542), .B1(n1566), .B2(n1537), .C1(n1650), 
        .C2(n1578), .ZN(n1799) );
  XNOR2_X1 U1413 ( .A(n1606), .B(n1800), .ZN(n850) );
  AOI221_X1 U1414 ( .B1(n1579), .B2(b[2]), .C1(n1580), .C2(b[1]), .A(n1801), 
        .ZN(n1800) );
  OAI22_X1 U1415 ( .A1(n1653), .A2(n1578), .B1(n1566), .B2(n1581), .ZN(n1801)
         );
  XNOR2_X1 U1416 ( .A(n1606), .B(n1803), .ZN(n849) );
  AOI221_X1 U1417 ( .B1(n1579), .B2(b[3]), .C1(n1580), .C2(b[2]), .A(n1804), 
        .ZN(n1803) );
  OAI22_X1 U1418 ( .A1(n1657), .A2(n1578), .B1(n1649), .B2(n1582), .ZN(n1804)
         );
  XNOR2_X1 U1419 ( .A(n1606), .B(n1805), .ZN(n848) );
  AOI221_X1 U1420 ( .B1(n1579), .B2(b[4]), .C1(n1580), .C2(b[3]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1421 ( .A1(n1660), .A2(n1578), .B1(n1661), .B2(n1582), .ZN(n1806)
         );
  XNOR2_X1 U1422 ( .A(n1606), .B(n1807), .ZN(n847) );
  AOI221_X1 U1423 ( .B1(n1579), .B2(b[5]), .C1(n1580), .C2(b[4]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1424 ( .A1(n1664), .A2(n1578), .B1(n1665), .B2(n1582), .ZN(n1808)
         );
  XNOR2_X1 U1425 ( .A(n1606), .B(n1809), .ZN(n846) );
  AOI221_X1 U1426 ( .B1(n1579), .B2(b[6]), .C1(n1580), .C2(b[5]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1427 ( .A1(n1668), .A2(n1578), .B1(n1669), .B2(n1582), .ZN(n1810)
         );
  XNOR2_X1 U1428 ( .A(n1606), .B(n1811), .ZN(n845) );
  AOI221_X1 U1429 ( .B1(n1579), .B2(b[7]), .C1(n1580), .C2(b[6]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1430 ( .A1(n1672), .A2(n1578), .B1(n1673), .B2(n1582), .ZN(n1812)
         );
  XNOR2_X1 U1431 ( .A(n1606), .B(n1813), .ZN(n844) );
  AOI221_X1 U1432 ( .B1(n1579), .B2(b[8]), .C1(n1580), .C2(b[7]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1433 ( .A1(n1676), .A2(n1578), .B1(n1677), .B2(n1582), .ZN(n1814)
         );
  XNOR2_X1 U1434 ( .A(n1606), .B(n1815), .ZN(n843) );
  AOI221_X1 U1435 ( .B1(n1579), .B2(b[9]), .C1(n1580), .C2(b[8]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1436 ( .A1(n1680), .A2(n1578), .B1(n1681), .B2(n1582), .ZN(n1816)
         );
  XNOR2_X1 U1437 ( .A(n1606), .B(n1817), .ZN(n842) );
  AOI221_X1 U1438 ( .B1(n1579), .B2(b[10]), .C1(n1580), .C2(b[9]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1439 ( .A1(n1684), .A2(n1578), .B1(n1685), .B2(n1582), .ZN(n1818)
         );
  XNOR2_X1 U1440 ( .A(n1606), .B(n1819), .ZN(n841) );
  AOI221_X1 U1441 ( .B1(n1579), .B2(b[11]), .C1(n1580), .C2(b[10]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1442 ( .A1(n1688), .A2(n1578), .B1(n1689), .B2(n1582), .ZN(n1820)
         );
  XNOR2_X1 U1443 ( .A(n1606), .B(n1821), .ZN(n840) );
  AOI221_X1 U1444 ( .B1(n1579), .B2(b[12]), .C1(n1580), .C2(b[11]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1445 ( .A1(n1692), .A2(n1578), .B1(n1693), .B2(n1582), .ZN(n1822)
         );
  XNOR2_X1 U1446 ( .A(n1606), .B(n1823), .ZN(n839) );
  AOI221_X1 U1447 ( .B1(n1579), .B2(b[13]), .C1(n1580), .C2(b[12]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1448 ( .A1(n1696), .A2(n1578), .B1(n1697), .B2(n1581), .ZN(n1824)
         );
  XNOR2_X1 U1449 ( .A(n1606), .B(n1825), .ZN(n838) );
  AOI221_X1 U1450 ( .B1(n1579), .B2(b[14]), .C1(n1580), .C2(b[13]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1451 ( .A1(n1700), .A2(n1578), .B1(n1701), .B2(n1581), .ZN(n1826)
         );
  XNOR2_X1 U1452 ( .A(n1606), .B(n1827), .ZN(n837) );
  AOI221_X1 U1453 ( .B1(n1579), .B2(b[15]), .C1(n1580), .C2(b[14]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1454 ( .A1(n1704), .A2(n1578), .B1(n1705), .B2(n1581), .ZN(n1828)
         );
  XNOR2_X1 U1455 ( .A(n1606), .B(n1829), .ZN(n836) );
  AOI221_X1 U1456 ( .B1(n1579), .B2(b[16]), .C1(n1580), .C2(b[15]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1457 ( .A1(n1708), .A2(n1578), .B1(n1709), .B2(n1581), .ZN(n1830)
         );
  XNOR2_X1 U1458 ( .A(n1606), .B(n1831), .ZN(n835) );
  AOI221_X1 U1459 ( .B1(n1579), .B2(b[17]), .C1(n1580), .C2(b[16]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1460 ( .A1(n1712), .A2(n1578), .B1(n1713), .B2(n1581), .ZN(n1832)
         );
  XNOR2_X1 U1461 ( .A(n1606), .B(n1833), .ZN(n834) );
  AOI221_X1 U1462 ( .B1(n1579), .B2(b[18]), .C1(n1580), .C2(b[17]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1463 ( .A1(n1716), .A2(n1578), .B1(n1717), .B2(n1581), .ZN(n1834)
         );
  XNOR2_X1 U1464 ( .A(n1606), .B(n1835), .ZN(n833) );
  AOI221_X1 U1465 ( .B1(n1579), .B2(b[19]), .C1(n1580), .C2(b[18]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1466 ( .A1(n1720), .A2(n1578), .B1(n1721), .B2(n1581), .ZN(n1836)
         );
  XNOR2_X1 U1467 ( .A(n1606), .B(n1837), .ZN(n832) );
  AOI221_X1 U1468 ( .B1(n1579), .B2(b[20]), .C1(n1580), .C2(b[19]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1469 ( .A1(n1724), .A2(n1578), .B1(n1725), .B2(n1581), .ZN(n1838)
         );
  XNOR2_X1 U1470 ( .A(a[11]), .B(n1839), .ZN(n831) );
  AOI221_X1 U1471 ( .B1(n1579), .B2(b[21]), .C1(n1580), .C2(b[20]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1472 ( .A1(n1728), .A2(n1578), .B1(n1729), .B2(n1581), .ZN(n1840)
         );
  XNOR2_X1 U1473 ( .A(a[11]), .B(n1841), .ZN(n830) );
  AOI221_X1 U1474 ( .B1(n1579), .B2(b[22]), .C1(n1546), .C2(n1376), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1475 ( .A1(n1640), .A2(n1582), .B1(n1643), .B2(n1537), .ZN(n1842)
         );
  XNOR2_X1 U1476 ( .A(a[11]), .B(n1843), .ZN(n829) );
  AOI221_X1 U1477 ( .B1(n1580), .B2(b[22]), .C1(n1546), .C2(n1375), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1478 ( .A1(n1617), .A2(n1542), .B1(n1643), .B2(n1581), .ZN(n1844)
         );
  XNOR2_X1 U1479 ( .A(a[11]), .B(n1845), .ZN(n828) );
  AOI221_X1 U1480 ( .B1(n1579), .B2(n1614), .C1(n1580), .C2(n1614), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1481 ( .A1(n1633), .A2(n1578), .B1(n1634), .B2(n1581), .ZN(n1846)
         );
  XNOR2_X1 U1482 ( .A(a[11]), .B(n1847), .ZN(n827) );
  OAI221_X1 U1483 ( .B1(n1616), .B2(n1582), .C1(n1617), .C2(n1578), .A(n1848), 
        .ZN(n1847) );
  OAI21_X1 U1484 ( .B1(n1579), .B2(n1580), .A(n1614), .ZN(n1848) );
  INV_X1 U1485 ( .A(n1852), .ZN(n1849) );
  NAND3_X1 U1486 ( .A1(n1852), .A2(n1851), .A3(n1850), .ZN(n1802) );
  XNOR2_X1 U1487 ( .A(a[10]), .B(a[9]), .ZN(n1850) );
  XNOR2_X1 U1488 ( .A(a[10]), .B(n1607), .ZN(n1851) );
  XOR2_X1 U1489 ( .A(a[9]), .B(n1609), .Z(n1852) );
  XNOR2_X1 U1490 ( .A(n1853), .B(n1605), .ZN(n826) );
  OAI22_X1 U1491 ( .A1(n1565), .A2(n1541), .B1(n1565), .B2(n1583), .ZN(n1853)
         );
  XNOR2_X1 U1492 ( .A(n1854), .B(n1605), .ZN(n825) );
  OAI222_X1 U1493 ( .A1(n1649), .A2(n1541), .B1(n1566), .B2(n1550), .C1(n1650), 
        .C2(n1583), .ZN(n1854) );
  XNOR2_X1 U1494 ( .A(n1604), .B(n1855), .ZN(n824) );
  AOI221_X1 U1495 ( .B1(n1584), .B2(b[2]), .C1(n1585), .C2(b[1]), .A(n1856), 
        .ZN(n1855) );
  OAI22_X1 U1496 ( .A1(n1653), .A2(n1583), .B1(n1565), .B2(n1586), .ZN(n1856)
         );
  XNOR2_X1 U1497 ( .A(n1604), .B(n1858), .ZN(n823) );
  AOI221_X1 U1498 ( .B1(n1584), .B2(b[3]), .C1(n1585), .C2(b[2]), .A(n1859), 
        .ZN(n1858) );
  OAI22_X1 U1499 ( .A1(n1657), .A2(n1583), .B1(n1649), .B2(n1587), .ZN(n1859)
         );
  XNOR2_X1 U1500 ( .A(n1604), .B(n1860), .ZN(n822) );
  AOI221_X1 U1501 ( .B1(n1584), .B2(b[4]), .C1(n1585), .C2(b[3]), .A(n1861), 
        .ZN(n1860) );
  OAI22_X1 U1502 ( .A1(n1660), .A2(n1583), .B1(n1661), .B2(n1587), .ZN(n1861)
         );
  XNOR2_X1 U1503 ( .A(n1604), .B(n1862), .ZN(n821) );
  AOI221_X1 U1504 ( .B1(n1584), .B2(b[5]), .C1(n1585), .C2(b[4]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1505 ( .A1(n1664), .A2(n1583), .B1(n1665), .B2(n1587), .ZN(n1863)
         );
  XNOR2_X1 U1506 ( .A(n1604), .B(n1864), .ZN(n820) );
  AOI221_X1 U1507 ( .B1(n1584), .B2(b[6]), .C1(n1585), .C2(b[5]), .A(n1865), 
        .ZN(n1864) );
  OAI22_X1 U1508 ( .A1(n1668), .A2(n1583), .B1(n1669), .B2(n1587), .ZN(n1865)
         );
  XNOR2_X1 U1509 ( .A(n1604), .B(n1866), .ZN(n819) );
  AOI221_X1 U1510 ( .B1(n1584), .B2(b[7]), .C1(n1585), .C2(b[6]), .A(n1867), 
        .ZN(n1866) );
  OAI22_X1 U1511 ( .A1(n1672), .A2(n1583), .B1(n1673), .B2(n1587), .ZN(n1867)
         );
  XNOR2_X1 U1512 ( .A(n1604), .B(n1868), .ZN(n818) );
  AOI221_X1 U1513 ( .B1(n1584), .B2(b[8]), .C1(n1585), .C2(b[7]), .A(n1869), 
        .ZN(n1868) );
  OAI22_X1 U1514 ( .A1(n1676), .A2(n1583), .B1(n1677), .B2(n1587), .ZN(n1869)
         );
  XNOR2_X1 U1515 ( .A(n1604), .B(n1870), .ZN(n817) );
  AOI221_X1 U1516 ( .B1(n1584), .B2(b[9]), .C1(n1585), .C2(b[8]), .A(n1871), 
        .ZN(n1870) );
  OAI22_X1 U1517 ( .A1(n1680), .A2(n1583), .B1(n1681), .B2(n1587), .ZN(n1871)
         );
  XNOR2_X1 U1518 ( .A(n1604), .B(n1872), .ZN(n816) );
  AOI221_X1 U1519 ( .B1(n1584), .B2(b[10]), .C1(n1585), .C2(b[9]), .A(n1873), 
        .ZN(n1872) );
  OAI22_X1 U1520 ( .A1(n1684), .A2(n1583), .B1(n1685), .B2(n1587), .ZN(n1873)
         );
  XNOR2_X1 U1521 ( .A(n1604), .B(n1874), .ZN(n815) );
  AOI221_X1 U1522 ( .B1(n1584), .B2(b[11]), .C1(n1585), .C2(b[10]), .A(n1875), 
        .ZN(n1874) );
  OAI22_X1 U1523 ( .A1(n1688), .A2(n1583), .B1(n1689), .B2(n1587), .ZN(n1875)
         );
  XNOR2_X1 U1524 ( .A(n1604), .B(n1876), .ZN(n814) );
  AOI221_X1 U1525 ( .B1(n1584), .B2(b[12]), .C1(n1585), .C2(b[11]), .A(n1877), 
        .ZN(n1876) );
  OAI22_X1 U1526 ( .A1(n1692), .A2(n1583), .B1(n1693), .B2(n1587), .ZN(n1877)
         );
  XNOR2_X1 U1527 ( .A(n1604), .B(n1878), .ZN(n813) );
  AOI221_X1 U1528 ( .B1(n1584), .B2(b[13]), .C1(n1585), .C2(b[12]), .A(n1879), 
        .ZN(n1878) );
  OAI22_X1 U1529 ( .A1(n1696), .A2(n1583), .B1(n1697), .B2(n1586), .ZN(n1879)
         );
  XNOR2_X1 U1530 ( .A(n1604), .B(n1880), .ZN(n812) );
  AOI221_X1 U1531 ( .B1(n1584), .B2(b[14]), .C1(n1585), .C2(b[13]), .A(n1881), 
        .ZN(n1880) );
  OAI22_X1 U1532 ( .A1(n1700), .A2(n1583), .B1(n1701), .B2(n1586), .ZN(n1881)
         );
  XNOR2_X1 U1533 ( .A(n1604), .B(n1882), .ZN(n811) );
  AOI221_X1 U1534 ( .B1(n1584), .B2(b[15]), .C1(n1585), .C2(b[14]), .A(n1883), 
        .ZN(n1882) );
  OAI22_X1 U1535 ( .A1(n1704), .A2(n1583), .B1(n1705), .B2(n1586), .ZN(n1883)
         );
  XNOR2_X1 U1536 ( .A(n1604), .B(n1884), .ZN(n810) );
  AOI221_X1 U1537 ( .B1(n1584), .B2(b[16]), .C1(n1585), .C2(b[15]), .A(n1885), 
        .ZN(n1884) );
  OAI22_X1 U1538 ( .A1(n1708), .A2(n1583), .B1(n1709), .B2(n1586), .ZN(n1885)
         );
  XNOR2_X1 U1539 ( .A(n1604), .B(n1886), .ZN(n809) );
  AOI221_X1 U1540 ( .B1(n1584), .B2(b[17]), .C1(n1585), .C2(b[16]), .A(n1887), 
        .ZN(n1886) );
  OAI22_X1 U1541 ( .A1(n1712), .A2(n1583), .B1(n1713), .B2(n1586), .ZN(n1887)
         );
  XNOR2_X1 U1542 ( .A(n1604), .B(n1888), .ZN(n808) );
  AOI221_X1 U1543 ( .B1(n1584), .B2(b[18]), .C1(n1585), .C2(b[17]), .A(n1889), 
        .ZN(n1888) );
  OAI22_X1 U1544 ( .A1(n1716), .A2(n1583), .B1(n1717), .B2(n1586), .ZN(n1889)
         );
  XNOR2_X1 U1545 ( .A(n1604), .B(n1890), .ZN(n807) );
  AOI221_X1 U1546 ( .B1(n1584), .B2(b[19]), .C1(n1585), .C2(b[18]), .A(n1891), 
        .ZN(n1890) );
  OAI22_X1 U1547 ( .A1(n1720), .A2(n1583), .B1(n1721), .B2(n1586), .ZN(n1891)
         );
  XNOR2_X1 U1548 ( .A(n1604), .B(n1892), .ZN(n806) );
  AOI221_X1 U1549 ( .B1(n1584), .B2(b[20]), .C1(n1585), .C2(b[19]), .A(n1893), 
        .ZN(n1892) );
  OAI22_X1 U1550 ( .A1(n1724), .A2(n1583), .B1(n1725), .B2(n1586), .ZN(n1893)
         );
  XNOR2_X1 U1551 ( .A(a[14]), .B(n1894), .ZN(n805) );
  AOI221_X1 U1552 ( .B1(n1584), .B2(b[21]), .C1(n1585), .C2(b[20]), .A(n1895), 
        .ZN(n1894) );
  OAI22_X1 U1553 ( .A1(n1728), .A2(n1583), .B1(n1729), .B2(n1586), .ZN(n1895)
         );
  XNOR2_X1 U1554 ( .A(a[14]), .B(n1896), .ZN(n804) );
  AOI221_X1 U1555 ( .B1(n1584), .B2(b[22]), .C1(n1553), .C2(n1376), .A(n1897), 
        .ZN(n1896) );
  OAI22_X1 U1556 ( .A1(n1640), .A2(n1587), .B1(n1643), .B2(n1550), .ZN(n1897)
         );
  XNOR2_X1 U1557 ( .A(a[14]), .B(n1898), .ZN(n803) );
  AOI221_X1 U1558 ( .B1(n1585), .B2(b[22]), .C1(n1553), .C2(n1375), .A(n1899), 
        .ZN(n1898) );
  OAI22_X1 U1559 ( .A1(n1617), .A2(n1541), .B1(n1643), .B2(n1586), .ZN(n1899)
         );
  XNOR2_X1 U1560 ( .A(a[14]), .B(n1900), .ZN(n802) );
  AOI221_X1 U1561 ( .B1(n1584), .B2(n1614), .C1(n1585), .C2(n1614), .A(n1901), 
        .ZN(n1900) );
  OAI22_X1 U1562 ( .A1(n1633), .A2(n1583), .B1(n1634), .B2(n1586), .ZN(n1901)
         );
  XNOR2_X1 U1563 ( .A(a[14]), .B(n1902), .ZN(n801) );
  OAI221_X1 U1564 ( .B1(n1617), .B2(n1587), .C1(n1619), .C2(n1583), .A(n1903), 
        .ZN(n1902) );
  OAI21_X1 U1565 ( .B1(n1584), .B2(n1585), .A(n1614), .ZN(n1903) );
  INV_X1 U1566 ( .A(n1907), .ZN(n1904) );
  NAND3_X1 U1567 ( .A1(n1907), .A2(n1906), .A3(n1905), .ZN(n1857) );
  XNOR2_X1 U1568 ( .A(a[12]), .B(a[13]), .ZN(n1905) );
  XNOR2_X1 U1569 ( .A(a[13]), .B(n1605), .ZN(n1906) );
  XOR2_X1 U1570 ( .A(a[12]), .B(n1607), .Z(n1907) );
  XNOR2_X1 U1571 ( .A(n1908), .B(n1603), .ZN(n800) );
  OAI22_X1 U1572 ( .A1(n1565), .A2(n1540), .B1(n1566), .B2(n1588), .ZN(n1908)
         );
  XNOR2_X1 U1573 ( .A(n1909), .B(n1603), .ZN(n799) );
  OAI222_X1 U1574 ( .A1(n1649), .A2(n1540), .B1(n1566), .B2(n1549), .C1(n1650), 
        .C2(n1588), .ZN(n1909) );
  XNOR2_X1 U1575 ( .A(n1602), .B(n1910), .ZN(n798) );
  AOI221_X1 U1576 ( .B1(n1589), .B2(b[2]), .C1(n1590), .C2(b[1]), .A(n1911), 
        .ZN(n1910) );
  OAI22_X1 U1577 ( .A1(n1653), .A2(n1588), .B1(n1566), .B2(n1591), .ZN(n1911)
         );
  XNOR2_X1 U1578 ( .A(n1602), .B(n1913), .ZN(n797) );
  AOI221_X1 U1579 ( .B1(n1589), .B2(b[3]), .C1(n1590), .C2(b[2]), .A(n1914), 
        .ZN(n1913) );
  OAI22_X1 U1580 ( .A1(n1657), .A2(n1588), .B1(n1649), .B2(n1592), .ZN(n1914)
         );
  XNOR2_X1 U1581 ( .A(n1602), .B(n1915), .ZN(n796) );
  AOI221_X1 U1582 ( .B1(n1589), .B2(b[4]), .C1(n1590), .C2(b[3]), .A(n1916), 
        .ZN(n1915) );
  OAI22_X1 U1583 ( .A1(n1660), .A2(n1588), .B1(n1661), .B2(n1592), .ZN(n1916)
         );
  XNOR2_X1 U1584 ( .A(n1602), .B(n1917), .ZN(n795) );
  AOI221_X1 U1585 ( .B1(n1589), .B2(b[5]), .C1(n1590), .C2(b[4]), .A(n1918), 
        .ZN(n1917) );
  OAI22_X1 U1586 ( .A1(n1664), .A2(n1588), .B1(n1665), .B2(n1592), .ZN(n1918)
         );
  XNOR2_X1 U1587 ( .A(n1602), .B(n1919), .ZN(n794) );
  AOI221_X1 U1588 ( .B1(n1589), .B2(b[6]), .C1(n1590), .C2(b[5]), .A(n1920), 
        .ZN(n1919) );
  OAI22_X1 U1589 ( .A1(n1668), .A2(n1588), .B1(n1669), .B2(n1592), .ZN(n1920)
         );
  XNOR2_X1 U1590 ( .A(n1602), .B(n1921), .ZN(n793) );
  AOI221_X1 U1591 ( .B1(n1589), .B2(b[7]), .C1(n1590), .C2(b[6]), .A(n1922), 
        .ZN(n1921) );
  OAI22_X1 U1592 ( .A1(n1672), .A2(n1588), .B1(n1673), .B2(n1592), .ZN(n1922)
         );
  XNOR2_X1 U1593 ( .A(n1602), .B(n1923), .ZN(n792) );
  AOI221_X1 U1594 ( .B1(n1589), .B2(b[8]), .C1(n1590), .C2(b[7]), .A(n1924), 
        .ZN(n1923) );
  OAI22_X1 U1595 ( .A1(n1676), .A2(n1588), .B1(n1677), .B2(n1592), .ZN(n1924)
         );
  XNOR2_X1 U1596 ( .A(n1602), .B(n1925), .ZN(n791) );
  AOI221_X1 U1597 ( .B1(n1589), .B2(b[9]), .C1(n1590), .C2(b[8]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1598 ( .A1(n1680), .A2(n1588), .B1(n1681), .B2(n1592), .ZN(n1926)
         );
  XNOR2_X1 U1599 ( .A(n1602), .B(n1927), .ZN(n790) );
  AOI221_X1 U1600 ( .B1(n1589), .B2(b[10]), .C1(n1590), .C2(b[9]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1601 ( .A1(n1684), .A2(n1588), .B1(n1685), .B2(n1592), .ZN(n1928)
         );
  XNOR2_X1 U1602 ( .A(n1602), .B(n1929), .ZN(n789) );
  AOI221_X1 U1603 ( .B1(n1589), .B2(b[11]), .C1(n1590), .C2(b[10]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1604 ( .A1(n1688), .A2(n1588), .B1(n1689), .B2(n1592), .ZN(n1930)
         );
  XNOR2_X1 U1605 ( .A(n1602), .B(n1931), .ZN(n788) );
  AOI221_X1 U1606 ( .B1(n1589), .B2(b[12]), .C1(n1590), .C2(b[11]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1607 ( .A1(n1692), .A2(n1588), .B1(n1693), .B2(n1592), .ZN(n1932)
         );
  XNOR2_X1 U1608 ( .A(n1602), .B(n1933), .ZN(n787) );
  AOI221_X1 U1609 ( .B1(n1589), .B2(b[13]), .C1(n1590), .C2(b[12]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1610 ( .A1(n1696), .A2(n1588), .B1(n1697), .B2(n1591), .ZN(n1934)
         );
  XNOR2_X1 U1611 ( .A(n1602), .B(n1935), .ZN(n786) );
  AOI221_X1 U1612 ( .B1(n1589), .B2(b[14]), .C1(n1590), .C2(b[13]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1613 ( .A1(n1700), .A2(n1588), .B1(n1701), .B2(n1591), .ZN(n1936)
         );
  XNOR2_X1 U1614 ( .A(n1602), .B(n1937), .ZN(n785) );
  AOI221_X1 U1615 ( .B1(n1589), .B2(b[15]), .C1(n1590), .C2(b[14]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1616 ( .A1(n1704), .A2(n1588), .B1(n1705), .B2(n1591), .ZN(n1938)
         );
  XNOR2_X1 U1617 ( .A(n1602), .B(n1939), .ZN(n784) );
  AOI221_X1 U1618 ( .B1(n1589), .B2(b[16]), .C1(n1590), .C2(b[15]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1619 ( .A1(n1708), .A2(n1588), .B1(n1709), .B2(n1591), .ZN(n1940)
         );
  XNOR2_X1 U1620 ( .A(n1602), .B(n1941), .ZN(n783) );
  AOI221_X1 U1621 ( .B1(n1589), .B2(b[17]), .C1(n1590), .C2(b[16]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1622 ( .A1(n1712), .A2(n1588), .B1(n1713), .B2(n1591), .ZN(n1942)
         );
  XNOR2_X1 U1623 ( .A(n1602), .B(n1943), .ZN(n782) );
  AOI221_X1 U1624 ( .B1(n1589), .B2(b[18]), .C1(n1590), .C2(b[17]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1625 ( .A1(n1716), .A2(n1588), .B1(n1717), .B2(n1591), .ZN(n1944)
         );
  XNOR2_X1 U1626 ( .A(n1602), .B(n1945), .ZN(n781) );
  AOI221_X1 U1627 ( .B1(n1589), .B2(b[19]), .C1(n1590), .C2(b[18]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1628 ( .A1(n1720), .A2(n1588), .B1(n1721), .B2(n1591), .ZN(n1946)
         );
  XNOR2_X1 U1629 ( .A(n1602), .B(n1947), .ZN(n780) );
  AOI221_X1 U1630 ( .B1(n1589), .B2(b[20]), .C1(n1590), .C2(b[19]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1631 ( .A1(n1724), .A2(n1588), .B1(n1725), .B2(n1591), .ZN(n1948)
         );
  XNOR2_X1 U1632 ( .A(a[17]), .B(n1949), .ZN(n779) );
  AOI221_X1 U1633 ( .B1(n1589), .B2(b[21]), .C1(n1590), .C2(b[20]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1634 ( .A1(n1728), .A2(n1588), .B1(n1729), .B2(n1591), .ZN(n1950)
         );
  XNOR2_X1 U1635 ( .A(a[17]), .B(n1951), .ZN(n778) );
  AOI221_X1 U1636 ( .B1(n1589), .B2(b[22]), .C1(n1552), .C2(n1376), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1637 ( .A1(n1640), .A2(n1592), .B1(n1643), .B2(n1549), .ZN(n1952)
         );
  XNOR2_X1 U1638 ( .A(a[17]), .B(n1953), .ZN(n777) );
  AOI221_X1 U1639 ( .B1(n1590), .B2(b[22]), .C1(n1552), .C2(n1375), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1640 ( .A1(n1617), .A2(n1540), .B1(n1643), .B2(n1591), .ZN(n1954)
         );
  XNOR2_X1 U1641 ( .A(a[17]), .B(n1955), .ZN(n776) );
  AOI221_X1 U1642 ( .B1(n1589), .B2(n1613), .C1(n1590), .C2(n1614), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1643 ( .A1(n1633), .A2(n1588), .B1(n1634), .B2(n1591), .ZN(n1956)
         );
  XNOR2_X1 U1644 ( .A(a[17]), .B(n1957), .ZN(n775) );
  OAI221_X1 U1645 ( .B1(n1618), .B2(n1592), .C1(n1617), .C2(n1588), .A(n1958), 
        .ZN(n1957) );
  OAI21_X1 U1646 ( .B1(n1589), .B2(n1590), .A(n1614), .ZN(n1958) );
  INV_X1 U1647 ( .A(n1962), .ZN(n1959) );
  NAND3_X1 U1648 ( .A1(n1962), .A2(n1961), .A3(n1960), .ZN(n1912) );
  XNOR2_X1 U1649 ( .A(a[15]), .B(a[16]), .ZN(n1960) );
  XNOR2_X1 U1650 ( .A(a[16]), .B(n1603), .ZN(n1961) );
  XOR2_X1 U1651 ( .A(a[15]), .B(n1605), .Z(n1962) );
  XOR2_X1 U1652 ( .A(n1963), .B(n1600), .Z(n774) );
  OAI22_X1 U1653 ( .A1(n1565), .A2(n1539), .B1(n1566), .B2(n1593), .ZN(n1963)
         );
  XOR2_X1 U1654 ( .A(n1964), .B(n1600), .Z(n773) );
  OAI222_X1 U1655 ( .A1(n1649), .A2(n1539), .B1(n1566), .B2(n1548), .C1(n1650), 
        .C2(n1593), .ZN(n1964) );
  XNOR2_X1 U1656 ( .A(n1600), .B(n1965), .ZN(n772) );
  AOI221_X1 U1657 ( .B1(n1594), .B2(b[2]), .C1(n1595), .C2(b[1]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1658 ( .A1(n1653), .A2(n1593), .B1(n1566), .B2(n1596), .ZN(n1966)
         );
  XNOR2_X1 U1659 ( .A(n1600), .B(n1968), .ZN(n771) );
  AOI221_X1 U1660 ( .B1(n1594), .B2(b[3]), .C1(n1595), .C2(b[2]), .A(n1969), 
        .ZN(n1968) );
  OAI22_X1 U1661 ( .A1(n1657), .A2(n1593), .B1(n1649), .B2(n1597), .ZN(n1969)
         );
  XNOR2_X1 U1662 ( .A(n1600), .B(n1970), .ZN(n770) );
  AOI221_X1 U1663 ( .B1(n1594), .B2(b[4]), .C1(n1595), .C2(b[3]), .A(n1971), 
        .ZN(n1970) );
  OAI22_X1 U1664 ( .A1(n1660), .A2(n1593), .B1(n1661), .B2(n1597), .ZN(n1971)
         );
  XNOR2_X1 U1665 ( .A(n1600), .B(n1972), .ZN(n769) );
  AOI221_X1 U1666 ( .B1(n1594), .B2(b[5]), .C1(n1595), .C2(b[4]), .A(n1973), 
        .ZN(n1972) );
  OAI22_X1 U1667 ( .A1(n1664), .A2(n1593), .B1(n1665), .B2(n1597), .ZN(n1973)
         );
  XNOR2_X1 U1668 ( .A(n1600), .B(n1974), .ZN(n768) );
  AOI221_X1 U1669 ( .B1(n1594), .B2(b[6]), .C1(n1595), .C2(b[5]), .A(n1975), 
        .ZN(n1974) );
  OAI22_X1 U1670 ( .A1(n1668), .A2(n1593), .B1(n1669), .B2(n1597), .ZN(n1975)
         );
  XNOR2_X1 U1671 ( .A(n1600), .B(n1976), .ZN(n767) );
  AOI221_X1 U1672 ( .B1(n1594), .B2(b[7]), .C1(n1595), .C2(b[6]), .A(n1977), 
        .ZN(n1976) );
  OAI22_X1 U1673 ( .A1(n1672), .A2(n1593), .B1(n1673), .B2(n1597), .ZN(n1977)
         );
  XNOR2_X1 U1674 ( .A(n1600), .B(n1978), .ZN(n766) );
  AOI221_X1 U1675 ( .B1(n1594), .B2(b[8]), .C1(n1595), .C2(b[7]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1676 ( .A1(n1676), .A2(n1593), .B1(n1677), .B2(n1597), .ZN(n1979)
         );
  XNOR2_X1 U1677 ( .A(n1600), .B(n1980), .ZN(n765) );
  AOI221_X1 U1678 ( .B1(n1594), .B2(b[9]), .C1(n1595), .C2(b[8]), .A(n1981), 
        .ZN(n1980) );
  OAI22_X1 U1679 ( .A1(n1680), .A2(n1593), .B1(n1681), .B2(n1597), .ZN(n1981)
         );
  XNOR2_X1 U1680 ( .A(n1600), .B(n1982), .ZN(n764) );
  AOI221_X1 U1681 ( .B1(n1594), .B2(b[10]), .C1(n1595), .C2(b[9]), .A(n1983), 
        .ZN(n1982) );
  OAI22_X1 U1682 ( .A1(n1684), .A2(n1593), .B1(n1685), .B2(n1597), .ZN(n1983)
         );
  XNOR2_X1 U1683 ( .A(n1600), .B(n1984), .ZN(n763) );
  AOI221_X1 U1684 ( .B1(n1594), .B2(b[11]), .C1(n1595), .C2(b[10]), .A(n1985), 
        .ZN(n1984) );
  OAI22_X1 U1685 ( .A1(n1688), .A2(n1593), .B1(n1689), .B2(n1597), .ZN(n1985)
         );
  XNOR2_X1 U1686 ( .A(n1601), .B(n1986), .ZN(n762) );
  AOI221_X1 U1687 ( .B1(n1594), .B2(b[12]), .C1(n1595), .C2(b[11]), .A(n1987), 
        .ZN(n1986) );
  OAI22_X1 U1688 ( .A1(n1692), .A2(n1593), .B1(n1693), .B2(n1597), .ZN(n1987)
         );
  XNOR2_X1 U1689 ( .A(n1601), .B(n1988), .ZN(n761) );
  AOI221_X1 U1690 ( .B1(n1594), .B2(b[13]), .C1(n1595), .C2(b[12]), .A(n1989), 
        .ZN(n1988) );
  OAI22_X1 U1691 ( .A1(n1696), .A2(n1593), .B1(n1697), .B2(n1596), .ZN(n1989)
         );
  XNOR2_X1 U1692 ( .A(n1601), .B(n1990), .ZN(n760) );
  AOI221_X1 U1693 ( .B1(n1594), .B2(b[14]), .C1(n1595), .C2(b[13]), .A(n1991), 
        .ZN(n1990) );
  OAI22_X1 U1694 ( .A1(n1700), .A2(n1593), .B1(n1701), .B2(n1596), .ZN(n1991)
         );
  XNOR2_X1 U1695 ( .A(n1601), .B(n1992), .ZN(n759) );
  AOI221_X1 U1696 ( .B1(n1594), .B2(b[15]), .C1(n1595), .C2(b[14]), .A(n1993), 
        .ZN(n1992) );
  OAI22_X1 U1697 ( .A1(n1704), .A2(n1593), .B1(n1705), .B2(n1596), .ZN(n1993)
         );
  XNOR2_X1 U1698 ( .A(n1601), .B(n1994), .ZN(n758) );
  AOI221_X1 U1699 ( .B1(n1594), .B2(b[16]), .C1(n1595), .C2(b[15]), .A(n1995), 
        .ZN(n1994) );
  OAI22_X1 U1700 ( .A1(n1708), .A2(n1593), .B1(n1709), .B2(n1596), .ZN(n1995)
         );
  XNOR2_X1 U1701 ( .A(n1601), .B(n1996), .ZN(n757) );
  AOI221_X1 U1702 ( .B1(n1594), .B2(b[17]), .C1(n1595), .C2(b[16]), .A(n1997), 
        .ZN(n1996) );
  OAI22_X1 U1703 ( .A1(n1712), .A2(n1593), .B1(n1713), .B2(n1596), .ZN(n1997)
         );
  XNOR2_X1 U1704 ( .A(n1601), .B(n1998), .ZN(n756) );
  AOI221_X1 U1705 ( .B1(n1594), .B2(b[18]), .C1(n1595), .C2(b[17]), .A(n1999), 
        .ZN(n1998) );
  OAI22_X1 U1706 ( .A1(n1716), .A2(n1593), .B1(n1717), .B2(n1596), .ZN(n1999)
         );
  XNOR2_X1 U1707 ( .A(n1601), .B(n2000), .ZN(n755) );
  AOI221_X1 U1708 ( .B1(n1594), .B2(b[19]), .C1(n1595), .C2(b[18]), .A(n2001), 
        .ZN(n2000) );
  OAI22_X1 U1709 ( .A1(n1720), .A2(n1593), .B1(n1721), .B2(n1596), .ZN(n2001)
         );
  XNOR2_X1 U1710 ( .A(n1601), .B(n2002), .ZN(n754) );
  AOI221_X1 U1711 ( .B1(n1594), .B2(b[20]), .C1(n1595), .C2(b[19]), .A(n2003), 
        .ZN(n2002) );
  OAI22_X1 U1712 ( .A1(n1724), .A2(n1593), .B1(n1725), .B2(n1596), .ZN(n2003)
         );
  XNOR2_X1 U1713 ( .A(n1601), .B(n2004), .ZN(n753) );
  AOI221_X1 U1714 ( .B1(n1594), .B2(b[21]), .C1(n1595), .C2(b[20]), .A(n2005), 
        .ZN(n2004) );
  OAI22_X1 U1715 ( .A1(n1728), .A2(n1593), .B1(n1729), .B2(n1596), .ZN(n2005)
         );
  XNOR2_X1 U1716 ( .A(n1601), .B(n2006), .ZN(n752) );
  AOI221_X1 U1717 ( .B1(n1594), .B2(b[22]), .C1(n1545), .C2(n1376), .A(n2007), 
        .ZN(n2006) );
  OAI22_X1 U1718 ( .A1(n1640), .A2(n1597), .B1(n1643), .B2(n1548), .ZN(n2007)
         );
  XNOR2_X1 U1719 ( .A(n1601), .B(n2008), .ZN(n751) );
  AOI221_X1 U1720 ( .B1(n1595), .B2(b[22]), .C1(n1545), .C2(n1375), .A(n2009), 
        .ZN(n2008) );
  OAI22_X1 U1721 ( .A1(n1617), .A2(n1539), .B1(n1643), .B2(n1596), .ZN(n2009)
         );
  XNOR2_X1 U1722 ( .A(n1601), .B(n2010), .ZN(n750) );
  AOI221_X1 U1723 ( .B1(n1594), .B2(n1612), .C1(n1595), .C2(n1614), .A(n2011), 
        .ZN(n2010) );
  OAI22_X1 U1724 ( .A1(n1633), .A2(n1593), .B1(n1634), .B2(n1596), .ZN(n2011)
         );
  INV_X1 U1725 ( .A(b[22]), .ZN(n1634) );
  INV_X1 U1726 ( .A(n1374), .ZN(n1633) );
  XNOR2_X1 U1727 ( .A(n1600), .B(n2012), .ZN(n749) );
  OAI221_X1 U1728 ( .B1(n1617), .B2(n1597), .C1(n1619), .C2(n1593), .A(n2013), 
        .ZN(n2012) );
  OAI21_X1 U1729 ( .B1(n1594), .B2(n1595), .A(n1614), .ZN(n2013) );
  INV_X1 U1730 ( .A(n2017), .ZN(n2014) );
  NAND3_X1 U1731 ( .A1(n2017), .A2(n2016), .A3(n2015), .ZN(n1967) );
  XNOR2_X1 U1732 ( .A(a[18]), .B(a[19]), .ZN(n2015) );
  XOR2_X1 U1733 ( .A(a[19]), .B(n1600), .Z(n2016) );
  XOR2_X1 U1734 ( .A(a[18]), .B(n1603), .Z(n2017) );
  XNOR2_X1 U1735 ( .A(n2018), .B(n1599), .ZN(n748) );
  OAI22_X1 U1736 ( .A1(n1538), .A2(n1567), .B1(n1558), .B2(n1567), .ZN(n2018)
         );
  XNOR2_X1 U1737 ( .A(n2019), .B(n1599), .ZN(n747) );
  OAI222_X1 U1738 ( .A1(n1538), .A2(n1649), .B1(n1547), .B2(n1566), .C1(n1558), 
        .C2(n1650), .ZN(n2019) );
  XNOR2_X1 U1739 ( .A(n1598), .B(n2020), .ZN(n746) );
  AOI221_X1 U1740 ( .B1(b[2]), .B2(n1559), .C1(b[1]), .C2(n1560), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1741 ( .A1(n1558), .A2(n1653), .B1(n1557), .B2(n1567), .ZN(n2021)
         );
  INV_X1 U1742 ( .A(b[0]), .ZN(n1647) );
  INV_X1 U1743 ( .A(n1396), .ZN(n1653) );
  XNOR2_X1 U1744 ( .A(n1598), .B(n2022), .ZN(n745) );
  AOI221_X1 U1745 ( .B1(b[3]), .B2(n1559), .C1(b[2]), .C2(n1560), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1746 ( .A1(n1558), .A2(n1657), .B1(n1557), .B2(n1649), .ZN(n2023)
         );
  XNOR2_X1 U1747 ( .A(n1598), .B(n2024), .ZN(n744) );
  AOI221_X1 U1748 ( .B1(b[4]), .B2(n1559), .C1(b[3]), .C2(n1560), .A(n2025), 
        .ZN(n2024) );
  OAI22_X1 U1749 ( .A1(n1558), .A2(n1660), .B1(n1557), .B2(n1661), .ZN(n2025)
         );
  XNOR2_X1 U1750 ( .A(n1598), .B(n2026), .ZN(n743) );
  AOI221_X1 U1751 ( .B1(b[5]), .B2(n1559), .C1(b[4]), .C2(n1560), .A(n2027), 
        .ZN(n2026) );
  OAI22_X1 U1752 ( .A1(n1558), .A2(n1664), .B1(n1557), .B2(n1665), .ZN(n2027)
         );
  XNOR2_X1 U1753 ( .A(n1598), .B(n2028), .ZN(n742) );
  AOI221_X1 U1754 ( .B1(b[6]), .B2(n1559), .C1(b[5]), .C2(n1560), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1755 ( .A1(n1558), .A2(n1668), .B1(n1557), .B2(n1669), .ZN(n2029)
         );
  XNOR2_X1 U1756 ( .A(n1598), .B(n2030), .ZN(n741) );
  AOI221_X1 U1757 ( .B1(b[7]), .B2(n1559), .C1(b[6]), .C2(n1560), .A(n2031), 
        .ZN(n2030) );
  OAI22_X1 U1758 ( .A1(n1558), .A2(n1672), .B1(n1557), .B2(n1673), .ZN(n2031)
         );
  XNOR2_X1 U1759 ( .A(n1598), .B(n2032), .ZN(n740) );
  AOI221_X1 U1760 ( .B1(b[9]), .B2(n1559), .C1(b[8]), .C2(n1560), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1761 ( .A1(n1558), .A2(n1680), .B1(n1557), .B2(n1681), .ZN(n2033)
         );
  XNOR2_X1 U1762 ( .A(n1598), .B(n2034), .ZN(n739) );
  AOI221_X1 U1763 ( .B1(b[10]), .B2(n1559), .C1(b[9]), .C2(n1560), .A(n2035), 
        .ZN(n2034) );
  OAI22_X1 U1764 ( .A1(n1558), .A2(n1684), .B1(n1557), .B2(n1685), .ZN(n2035)
         );
  XNOR2_X1 U1765 ( .A(n1598), .B(n2036), .ZN(n738) );
  AOI221_X1 U1766 ( .B1(b[12]), .B2(n1559), .C1(b[11]), .C2(n1560), .A(n2037), 
        .ZN(n2036) );
  OAI22_X1 U1767 ( .A1(n1558), .A2(n1692), .B1(n1557), .B2(n1693), .ZN(n2037)
         );
  XNOR2_X1 U1768 ( .A(n1598), .B(n2038), .ZN(n737) );
  AOI221_X1 U1769 ( .B1(b[13]), .B2(n1559), .C1(b[12]), .C2(n1560), .A(n2039), 
        .ZN(n2038) );
  OAI22_X1 U1770 ( .A1(n1558), .A2(n1696), .B1(n1557), .B2(n1697), .ZN(n2039)
         );
  XNOR2_X1 U1771 ( .A(n1598), .B(n2040), .ZN(n736) );
  AOI221_X1 U1772 ( .B1(b[14]), .B2(n1559), .C1(b[13]), .C2(n1560), .A(n2041), 
        .ZN(n2040) );
  OAI22_X1 U1773 ( .A1(n1558), .A2(n1700), .B1(n1556), .B2(n1701), .ZN(n2041)
         );
  XNOR2_X1 U1774 ( .A(n1598), .B(n2042), .ZN(n735) );
  AOI221_X1 U1775 ( .B1(b[15]), .B2(n1559), .C1(b[14]), .C2(n1560), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1776 ( .A1(n1558), .A2(n1704), .B1(n1556), .B2(n1705), .ZN(n2043)
         );
  XNOR2_X1 U1777 ( .A(n1598), .B(n2044), .ZN(n734) );
  AOI221_X1 U1778 ( .B1(b[16]), .B2(n1559), .C1(b[15]), .C2(n1560), .A(n2045), 
        .ZN(n2044) );
  OAI22_X1 U1779 ( .A1(n1558), .A2(n1708), .B1(n1556), .B2(n1709), .ZN(n2045)
         );
  XNOR2_X1 U1780 ( .A(n1598), .B(n2046), .ZN(n733) );
  AOI221_X1 U1781 ( .B1(b[18]), .B2(n1559), .C1(b[17]), .C2(n1560), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1782 ( .A1(n1558), .A2(n1716), .B1(n1556), .B2(n1717), .ZN(n2047)
         );
  XNOR2_X1 U1783 ( .A(n1598), .B(n2048), .ZN(n732) );
  AOI221_X1 U1784 ( .B1(b[19]), .B2(n1559), .C1(b[18]), .C2(n1560), .A(n2049), 
        .ZN(n2048) );
  OAI22_X1 U1785 ( .A1(n1558), .A2(n1720), .B1(n1556), .B2(n1721), .ZN(n2049)
         );
  XNOR2_X1 U1786 ( .A(n1598), .B(n2050), .ZN(n731) );
  AOI221_X1 U1787 ( .B1(b[20]), .B2(n1559), .C1(b[19]), .C2(n1560), .A(n2051), 
        .ZN(n2050) );
  OAI22_X1 U1788 ( .A1(n1558), .A2(n1724), .B1(n1556), .B2(n1725), .ZN(n2051)
         );
  XNOR2_X1 U1789 ( .A(a[23]), .B(n2052), .ZN(n730) );
  AOI221_X1 U1790 ( .B1(b[21]), .B2(n1559), .C1(b[20]), .C2(n1560), .A(n2053), 
        .ZN(n2052) );
  OAI22_X1 U1791 ( .A1(n1558), .A2(n1728), .B1(n1556), .B2(n1729), .ZN(n2053)
         );
  XNOR2_X1 U1792 ( .A(a[23]), .B(n2054), .ZN(n729) );
  AOI221_X1 U1793 ( .B1(b[22]), .B2(n1559), .C1(n1376), .C2(n1544), .A(n2055), 
        .ZN(n2054) );
  OAI22_X1 U1794 ( .A1(n1556), .A2(n1640), .B1(n1547), .B2(n1643), .ZN(n2055)
         );
  INV_X1 U1795 ( .A(b[20]), .ZN(n1640) );
  XNOR2_X1 U1796 ( .A(n519), .B(n2056), .ZN(n506) );
  INV_X1 U1797 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1798 ( .A1(n2056), .A2(n519), .ZN(n493) );
  XOR2_X1 U1799 ( .A(n2057), .B(n1742), .Z(n2056) );
  OAI221_X1 U1800 ( .B1(n1618), .B2(n1639), .C1(n1619), .C2(n1564), .A(n2058), 
        .ZN(n2057) );
  OAI21_X1 U1801 ( .B1(n1561), .B2(n1563), .A(n1614), .ZN(n2058) );
  INV_X1 U1802 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1803 ( .A(n1598), .B(n2059), .Z(n454) );
  AOI221_X1 U1804 ( .B1(b[8]), .B2(n1559), .C1(b[7]), .C2(n1560), .A(n2060), 
        .ZN(n2059) );
  OAI22_X1 U1805 ( .A1(n1558), .A2(n1676), .B1(n1556), .B2(n1677), .ZN(n2060)
         );
  INV_X1 U1806 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1807 ( .A(n1598), .B(n2061), .Z(n421) );
  AOI221_X1 U1808 ( .B1(b[11]), .B2(n1559), .C1(b[10]), .C2(n1560), .A(n2062), 
        .ZN(n2061) );
  OAI22_X1 U1809 ( .A1(n1558), .A2(n1688), .B1(n1556), .B2(n1689), .ZN(n2062)
         );
  INV_X1 U1810 ( .A(n387), .ZN(n395) );
  INV_X1 U1811 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1812 ( .A(n1598), .B(n2063), .Z(n374) );
  AOI221_X1 U1813 ( .B1(b[17]), .B2(n1559), .C1(b[16]), .C2(n1560), .A(n2064), 
        .ZN(n2063) );
  OAI22_X1 U1814 ( .A1(n1558), .A2(n1712), .B1(n1556), .B2(n1713), .ZN(n2064)
         );
  INV_X1 U1815 ( .A(n356), .ZN(n360) );
  INV_X1 U1816 ( .A(n1627), .ZN(n351) );
  XOR2_X1 U1817 ( .A(n1599), .B(n2065), .Z(n1627) );
  AOI221_X1 U1818 ( .B1(b[22]), .B2(n1560), .C1(n1375), .C2(n1544), .A(n2066), 
        .ZN(n2065) );
  OAI22_X1 U1819 ( .A1(n1538), .A2(n1618), .B1(n1556), .B2(n1643), .ZN(n2066)
         );
  INV_X1 U1820 ( .A(b[21]), .ZN(n1643) );
  NAND3_X1 U1821 ( .A1(n2067), .A2(n2068), .A3(n2069), .ZN(n1629) );
  XNOR2_X1 U1822 ( .A(a[22]), .B(n1599), .ZN(n2068) );
  XNOR2_X1 U1823 ( .A(a[21]), .B(a[22]), .ZN(n2069) );
  INV_X1 U1824 ( .A(n2067), .ZN(n2070) );
  XNOR2_X1 U1825 ( .A(a[21]), .B(n1600), .ZN(n2067) );
  OAI222_X1 U1826 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n2073), .C1(n2073), 
        .C2(n2072), .ZN(n326) );
  INV_X1 U1827 ( .A(n550), .ZN(n2073) );
  XNOR2_X1 U1828 ( .A(n1742), .B(n2074), .ZN(n2072) );
  AOI221_X1 U1829 ( .B1(n1561), .B2(b[21]), .C1(b[20]), .C2(n1562), .A(n2075), 
        .ZN(n2074) );
  OAI22_X1 U1830 ( .A1(n1564), .A2(n1728), .B1(n1639), .B2(n1729), .ZN(n2075)
         );
  INV_X1 U1831 ( .A(b[19]), .ZN(n1729) );
  INV_X1 U1832 ( .A(n1377), .ZN(n1728) );
  AOI222_X1 U1833 ( .A1(n2076), .A2(n2077), .B1(n2076), .B2(n564), .C1(n564), 
        .C2(n2077), .ZN(n2071) );
  XNOR2_X1 U1834 ( .A(a[2]), .B(n2078), .ZN(n2077) );
  AOI221_X1 U1835 ( .B1(b[20]), .B2(n1561), .C1(b[19]), .C2(n1562), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1836 ( .A1(n1564), .A2(n1724), .B1(n1639), .B2(n1725), .ZN(n2079)
         );
  INV_X1 U1837 ( .A(b[18]), .ZN(n1725) );
  INV_X1 U1838 ( .A(n1378), .ZN(n1724) );
  INV_X1 U1839 ( .A(n2080), .ZN(n2076) );
  AOI222_X1 U1840 ( .A1(n2081), .A2(n2082), .B1(n2081), .B2(n576), .C1(n576), 
        .C2(n2082), .ZN(n2080) );
  XNOR2_X1 U1841 ( .A(a[2]), .B(n2083), .ZN(n2082) );
  AOI221_X1 U1842 ( .B1(b[19]), .B2(n1561), .C1(b[18]), .C2(n1562), .A(n2084), 
        .ZN(n2083) );
  OAI22_X1 U1843 ( .A1(n1564), .A2(n1720), .B1(n1639), .B2(n1721), .ZN(n2084)
         );
  INV_X1 U1844 ( .A(b[17]), .ZN(n1721) );
  INV_X1 U1845 ( .A(n1379), .ZN(n1720) );
  OAI222_X1 U1846 ( .A1(n2085), .A2(n2086), .B1(n2085), .B2(n2087), .C1(n2087), 
        .C2(n2086), .ZN(n2081) );
  INV_X1 U1847 ( .A(n588), .ZN(n2087) );
  XNOR2_X1 U1848 ( .A(n1742), .B(n2088), .ZN(n2086) );
  AOI221_X1 U1849 ( .B1(b[18]), .B2(n1561), .C1(b[17]), .C2(n1562), .A(n2089), 
        .ZN(n2088) );
  OAI22_X1 U1850 ( .A1(n1564), .A2(n1716), .B1(n1639), .B2(n1717), .ZN(n2089)
         );
  INV_X1 U1851 ( .A(b[16]), .ZN(n1717) );
  INV_X1 U1852 ( .A(n1380), .ZN(n1716) );
  AOI222_X1 U1853 ( .A1(n2090), .A2(n2091), .B1(n2090), .B2(n600), .C1(n600), 
        .C2(n2091), .ZN(n2085) );
  XNOR2_X1 U1854 ( .A(a[2]), .B(n2092), .ZN(n2091) );
  AOI221_X1 U1855 ( .B1(b[17]), .B2(n1561), .C1(b[16]), .C2(n1562), .A(n2093), 
        .ZN(n2092) );
  OAI22_X1 U1856 ( .A1(n1564), .A2(n1712), .B1(n1639), .B2(n1713), .ZN(n2093)
         );
  INV_X1 U1857 ( .A(b[15]), .ZN(n1713) );
  INV_X1 U1858 ( .A(n1381), .ZN(n1712) );
  OAI222_X1 U1859 ( .A1(n2094), .A2(n2095), .B1(n2094), .B2(n2096), .C1(n2096), 
        .C2(n2095), .ZN(n2090) );
  INV_X1 U1860 ( .A(n610), .ZN(n2096) );
  XNOR2_X1 U1861 ( .A(n1742), .B(n2097), .ZN(n2095) );
  AOI221_X1 U1862 ( .B1(b[16]), .B2(n1561), .C1(b[15]), .C2(n1562), .A(n2098), 
        .ZN(n2097) );
  OAI22_X1 U1863 ( .A1(n1564), .A2(n1708), .B1(n1639), .B2(n1709), .ZN(n2098)
         );
  INV_X1 U1864 ( .A(b[14]), .ZN(n1709) );
  INV_X1 U1865 ( .A(n1382), .ZN(n1708) );
  AOI222_X1 U1866 ( .A1(n2099), .A2(n2100), .B1(n2099), .B2(n620), .C1(n620), 
        .C2(n2100), .ZN(n2094) );
  XNOR2_X1 U1867 ( .A(a[2]), .B(n2101), .ZN(n2100) );
  AOI221_X1 U1868 ( .B1(b[15]), .B2(n1561), .C1(b[14]), .C2(n1562), .A(n2102), 
        .ZN(n2101) );
  OAI22_X1 U1869 ( .A1(n1564), .A2(n1704), .B1(n1639), .B2(n1705), .ZN(n2102)
         );
  INV_X1 U1870 ( .A(b[13]), .ZN(n1705) );
  INV_X1 U1871 ( .A(n1383), .ZN(n1704) );
  OAI222_X1 U1872 ( .A1(n2103), .A2(n2104), .B1(n2103), .B2(n2105), .C1(n2105), 
        .C2(n2104), .ZN(n2099) );
  INV_X1 U1873 ( .A(n630), .ZN(n2105) );
  XNOR2_X1 U1874 ( .A(n1742), .B(n2106), .ZN(n2104) );
  AOI221_X1 U1875 ( .B1(b[14]), .B2(n1561), .C1(b[13]), .C2(n1562), .A(n2107), 
        .ZN(n2106) );
  OAI22_X1 U1876 ( .A1(n1564), .A2(n1700), .B1(n1639), .B2(n1701), .ZN(n2107)
         );
  INV_X1 U1877 ( .A(b[12]), .ZN(n1701) );
  INV_X1 U1878 ( .A(n1384), .ZN(n1700) );
  AOI222_X1 U1879 ( .A1(n2108), .A2(n2109), .B1(n2108), .B2(n638), .C1(n638), 
        .C2(n2109), .ZN(n2103) );
  XNOR2_X1 U1880 ( .A(a[2]), .B(n2110), .ZN(n2109) );
  AOI221_X1 U1881 ( .B1(b[13]), .B2(n1561), .C1(b[12]), .C2(n1562), .A(n2111), 
        .ZN(n2110) );
  OAI22_X1 U1882 ( .A1(n1564), .A2(n1696), .B1(n1639), .B2(n1697), .ZN(n2111)
         );
  INV_X1 U1883 ( .A(b[11]), .ZN(n1697) );
  INV_X1 U1884 ( .A(n1385), .ZN(n1696) );
  OAI222_X1 U1885 ( .A1(n2112), .A2(n2113), .B1(n2112), .B2(n2114), .C1(n2114), 
        .C2(n2113), .ZN(n2108) );
  INV_X1 U1886 ( .A(n646), .ZN(n2114) );
  XNOR2_X1 U1887 ( .A(n1742), .B(n2115), .ZN(n2113) );
  AOI221_X1 U1888 ( .B1(b[12]), .B2(n1561), .C1(b[11]), .C2(n1562), .A(n2116), 
        .ZN(n2115) );
  OAI22_X1 U1889 ( .A1(n1564), .A2(n1692), .B1(n1639), .B2(n1693), .ZN(n2116)
         );
  INV_X1 U1890 ( .A(b[10]), .ZN(n1693) );
  INV_X1 U1891 ( .A(n1386), .ZN(n1692) );
  AOI222_X1 U1892 ( .A1(n2117), .A2(n2118), .B1(n2117), .B2(n654), .C1(n654), 
        .C2(n2118), .ZN(n2112) );
  XNOR2_X1 U1893 ( .A(a[2]), .B(n2119), .ZN(n2118) );
  AOI221_X1 U1894 ( .B1(b[11]), .B2(n1561), .C1(b[10]), .C2(n1562), .A(n2120), 
        .ZN(n2119) );
  OAI22_X1 U1895 ( .A1(n1564), .A2(n1688), .B1(n1639), .B2(n1689), .ZN(n2120)
         );
  INV_X1 U1896 ( .A(b[9]), .ZN(n1689) );
  INV_X1 U1897 ( .A(n1387), .ZN(n1688) );
  OAI222_X1 U1898 ( .A1(n2121), .A2(n2122), .B1(n2121), .B2(n2123), .C1(n2123), 
        .C2(n2122), .ZN(n2117) );
  INV_X1 U1899 ( .A(n660), .ZN(n2123) );
  XNOR2_X1 U1900 ( .A(n1742), .B(n2124), .ZN(n2122) );
  AOI221_X1 U1901 ( .B1(b[10]), .B2(n1561), .C1(b[9]), .C2(n1563), .A(n2125), 
        .ZN(n2124) );
  OAI22_X1 U1902 ( .A1(n1564), .A2(n1684), .B1(n1639), .B2(n1685), .ZN(n2125)
         );
  INV_X1 U1903 ( .A(b[8]), .ZN(n1685) );
  INV_X1 U1904 ( .A(n1388), .ZN(n1684) );
  AOI222_X1 U1905 ( .A1(n2126), .A2(n2127), .B1(n2126), .B2(n666), .C1(n666), 
        .C2(n2127), .ZN(n2121) );
  XNOR2_X1 U1906 ( .A(a[2]), .B(n2128), .ZN(n2127) );
  AOI221_X1 U1907 ( .B1(b[9]), .B2(n1561), .C1(b[8]), .C2(n1563), .A(n2129), 
        .ZN(n2128) );
  OAI22_X1 U1908 ( .A1(n1564), .A2(n1680), .B1(n1639), .B2(n1681), .ZN(n2129)
         );
  INV_X1 U1909 ( .A(b[7]), .ZN(n1681) );
  INV_X1 U1910 ( .A(n1389), .ZN(n1680) );
  OAI222_X1 U1911 ( .A1(n2130), .A2(n2131), .B1(n2130), .B2(n2132), .C1(n2132), 
        .C2(n2131), .ZN(n2126) );
  INV_X1 U1912 ( .A(n672), .ZN(n2132) );
  XNOR2_X1 U1913 ( .A(n1742), .B(n2133), .ZN(n2131) );
  AOI221_X1 U1914 ( .B1(b[8]), .B2(n1561), .C1(b[7]), .C2(n1562), .A(n2134), 
        .ZN(n2133) );
  OAI22_X1 U1915 ( .A1(n1564), .A2(n1676), .B1(n1639), .B2(n1677), .ZN(n2134)
         );
  INV_X1 U1916 ( .A(b[6]), .ZN(n1677) );
  INV_X1 U1917 ( .A(n1390), .ZN(n1676) );
  AOI222_X1 U1918 ( .A1(n2135), .A2(n2136), .B1(n2135), .B2(n676), .C1(n676), 
        .C2(n2136), .ZN(n2130) );
  XNOR2_X1 U1919 ( .A(a[2]), .B(n2137), .ZN(n2136) );
  AOI221_X1 U1920 ( .B1(b[7]), .B2(n1561), .C1(b[6]), .C2(n1563), .A(n2138), 
        .ZN(n2137) );
  OAI22_X1 U1921 ( .A1(n1564), .A2(n1672), .B1(n1639), .B2(n1673), .ZN(n2138)
         );
  INV_X1 U1922 ( .A(b[5]), .ZN(n1673) );
  INV_X1 U1923 ( .A(n1391), .ZN(n1672) );
  OAI222_X1 U1924 ( .A1(n2139), .A2(n2140), .B1(n2139), .B2(n2141), .C1(n2141), 
        .C2(n2140), .ZN(n2135) );
  INV_X1 U1925 ( .A(n680), .ZN(n2141) );
  XNOR2_X1 U1926 ( .A(n1742), .B(n2142), .ZN(n2140) );
  AOI221_X1 U1927 ( .B1(b[6]), .B2(n1561), .C1(b[5]), .C2(n1563), .A(n2143), 
        .ZN(n2142) );
  OAI22_X1 U1928 ( .A1(n1564), .A2(n1668), .B1(n1639), .B2(n1669), .ZN(n2143)
         );
  INV_X1 U1929 ( .A(b[4]), .ZN(n1669) );
  INV_X1 U1930 ( .A(n1392), .ZN(n1668) );
  AOI222_X1 U1931 ( .A1(n2144), .A2(n2145), .B1(n2144), .B2(n684), .C1(n684), 
        .C2(n2145), .ZN(n2139) );
  XNOR2_X1 U1932 ( .A(a[2]), .B(n2146), .ZN(n2145) );
  AOI221_X1 U1933 ( .B1(b[5]), .B2(n1561), .C1(b[4]), .C2(n1563), .A(n2147), 
        .ZN(n2146) );
  OAI22_X1 U1934 ( .A1(n1564), .A2(n1664), .B1(n1639), .B2(n1665), .ZN(n2147)
         );
  INV_X1 U1935 ( .A(b[3]), .ZN(n1665) );
  INV_X1 U1936 ( .A(n1393), .ZN(n1664) );
  OAI222_X1 U1937 ( .A1(n2148), .A2(n2149), .B1(n2148), .B2(n2150), .C1(n2150), 
        .C2(n2149), .ZN(n2144) );
  INV_X1 U1938 ( .A(n686), .ZN(n2150) );
  XNOR2_X1 U1939 ( .A(n1742), .B(n2151), .ZN(n2149) );
  AOI221_X1 U1940 ( .B1(b[4]), .B2(n1561), .C1(b[3]), .C2(n1563), .A(n2152), 
        .ZN(n2151) );
  OAI22_X1 U1941 ( .A1(n1564), .A2(n1660), .B1(n1639), .B2(n1661), .ZN(n2152)
         );
  INV_X1 U1942 ( .A(n1394), .ZN(n1660) );
  AOI222_X1 U1943 ( .A1(n2153), .A2(n2154), .B1(n2153), .B2(n688), .C1(n688), 
        .C2(n2154), .ZN(n2148) );
  XNOR2_X1 U1944 ( .A(a[2]), .B(n2155), .ZN(n2154) );
  AOI221_X1 U1945 ( .B1(b[3]), .B2(n1561), .C1(b[2]), .C2(n1563), .A(n2156), 
        .ZN(n2155) );
  OAI22_X1 U1946 ( .A1(n1564), .A2(n1657), .B1(n1639), .B2(n1649), .ZN(n2156)
         );
  INV_X1 U1947 ( .A(b[1]), .ZN(n1649) );
  INV_X1 U1948 ( .A(n1395), .ZN(n1657) );
  AND2_X1 U1949 ( .A1(n2160), .A2(n2161), .ZN(n2153) );
  AOI211_X1 U1950 ( .C1(b[1]), .C2(n1561), .A(n2162), .B(b[0]), .ZN(n2161) );
  OAI22_X1 U1951 ( .A1(n1535), .A2(n1661), .B1(n1564), .B2(n1650), .ZN(n2162)
         );
  INV_X1 U1952 ( .A(n1397), .ZN(n1650) );
  INV_X1 U1953 ( .A(b[2]), .ZN(n1661) );
  INV_X1 U1954 ( .A(a[0]), .ZN(n2158) );
  AOI221_X1 U1955 ( .B1(b[1]), .B2(n1563), .C1(n1396), .C2(n1555), .A(n1742), 
        .ZN(n2160) );
  XNOR2_X1 U1956 ( .A(a[1]), .B(n1742), .ZN(n2157) );
  INV_X1 U1957 ( .A(a[2]), .ZN(n1742) );
  NOR2_X1 U1958 ( .A1(n2159), .A2(a[0]), .ZN(n1636) );
  INV_X1 U1959 ( .A(a[1]), .ZN(n2159) );
endmodule


module iir_filter_DW_mult_tc_1 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(product[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(product[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(product[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(product[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(product[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(product[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(product[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(product[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(product[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(product[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(product[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(product[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(product[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(product[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(product[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(product[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(product[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(product[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(product[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(product[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(product[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(product[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(product[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1598), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1600), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1602), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1604), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1606), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1608), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1610), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(b[22]), .B(n1614), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(b[21]), .B(b[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(b[20]), .B(b[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(b[19]), .B(b[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(b[18]), .B(b[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(b[17]), .B(b[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(b[16]), .B(b[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(b[15]), .B(b[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(b[14]), .B(b[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(b[13]), .B(b[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(b[12]), .B(b[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(b[11]), .B(b[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(b[10]), .B(b[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(b[9]), .B(b[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(b[8]), .B(b[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(b[7]), .B(b[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(b[6]), .B(b[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(b[5]), .B(b[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(b[4]), .B(b[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(b[3]), .B(b[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(b[2]), .B(b[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(b[1]), .B(b[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(b[0]), .B(b[1]), .CO(n727), .S(n1397) );
  INV_X1 U1137 ( .A(n1533), .ZN(n1570) );
  INV_X1 U1138 ( .A(n1536), .ZN(n1568) );
  INV_X1 U1139 ( .A(n1535), .ZN(n1561) );
  INV_X1 U1140 ( .A(n1534), .ZN(n1569) );
  BUF_X1 U1141 ( .A(n1654), .Z(n1572) );
  INV_X1 U1142 ( .A(n1547), .ZN(n1560) );
  INV_X1 U1143 ( .A(n1544), .ZN(n1558) );
  INV_X1 U1144 ( .A(n1537), .ZN(n1580) );
  INV_X1 U1145 ( .A(n1551), .ZN(n1575) );
  INV_X1 U1146 ( .A(n1550), .ZN(n1585) );
  INV_X1 U1147 ( .A(n1548), .ZN(n1595) );
  INV_X1 U1148 ( .A(n1549), .ZN(n1590) );
  INV_X1 U1149 ( .A(n1538), .ZN(n1559) );
  INV_X1 U1150 ( .A(n1545), .ZN(n1593) );
  INV_X1 U1151 ( .A(n1553), .ZN(n1583) );
  INV_X1 U1152 ( .A(n1552), .ZN(n1588) );
  INV_X1 U1153 ( .A(n1546), .ZN(n1578) );
  INV_X1 U1154 ( .A(n1554), .ZN(n1573) );
  BUF_X1 U1155 ( .A(n1654), .Z(n1571) );
  BUF_X1 U1156 ( .A(n1629), .Z(n1557) );
  BUF_X1 U1157 ( .A(n1967), .Z(n1596) );
  BUF_X1 U1158 ( .A(n1912), .Z(n1591) );
  BUF_X1 U1159 ( .A(n1857), .Z(n1586) );
  BUF_X1 U1160 ( .A(n1802), .Z(n1581) );
  BUF_X1 U1161 ( .A(n1747), .Z(n1576) );
  BUF_X1 U1162 ( .A(n1912), .Z(n1592) );
  BUF_X1 U1163 ( .A(n1857), .Z(n1587) );
  BUF_X1 U1164 ( .A(n1802), .Z(n1582) );
  BUF_X1 U1165 ( .A(n1747), .Z(n1577) );
  BUF_X1 U1166 ( .A(n1967), .Z(n1597) );
  INV_X1 U1167 ( .A(n1615), .ZN(n1614) );
  INV_X1 U1168 ( .A(n1540), .ZN(n1589) );
  INV_X1 U1169 ( .A(n1541), .ZN(n1584) );
  INV_X1 U1170 ( .A(n1542), .ZN(n1579) );
  INV_X1 U1171 ( .A(n1543), .ZN(n1574) );
  BUF_X1 U1172 ( .A(n1629), .Z(n1556) );
  INV_X1 U1173 ( .A(n1539), .ZN(n1594) );
  NAND3_X1 U1174 ( .A1(n2157), .A2(n2158), .A3(n2159), .ZN(n1639) );
  INV_X1 U1175 ( .A(n1555), .ZN(n1564) );
  OR2_X1 U1176 ( .A1(n1738), .A2(n1739), .ZN(n1533) );
  OR2_X1 U1177 ( .A1(n1740), .A2(n1741), .ZN(n1534) );
  OR2_X1 U1178 ( .A1(n2158), .A2(n2157), .ZN(n1535) );
  AND2_X1 U1179 ( .A1(n1738), .A2(n1740), .ZN(n1536) );
  INV_X1 U1180 ( .A(n1611), .ZN(n1610) );
  INV_X1 U1181 ( .A(n1607), .ZN(n1606) );
  INV_X1 U1182 ( .A(n1609), .ZN(n1608) );
  INV_X1 U1183 ( .A(n1603), .ZN(n1602) );
  INV_X1 U1184 ( .A(n1605), .ZN(n1604) );
  OR2_X1 U1185 ( .A1(n1849), .A2(n1850), .ZN(n1537) );
  BUF_X1 U1186 ( .A(n1636), .Z(n1562) );
  BUF_X1 U1187 ( .A(n1636), .Z(n1563) );
  BUF_X1 U1188 ( .A(n1647), .Z(n1565) );
  BUF_X1 U1189 ( .A(n1647), .Z(n1566) );
  OR2_X1 U1190 ( .A1(n2068), .A2(n2067), .ZN(n1538) );
  OR2_X1 U1191 ( .A1(n2016), .A2(n2017), .ZN(n1539) );
  OR2_X1 U1192 ( .A1(n1961), .A2(n1962), .ZN(n1540) );
  OR2_X1 U1193 ( .A1(n1906), .A2(n1907), .ZN(n1541) );
  OR2_X1 U1194 ( .A1(n1851), .A2(n1852), .ZN(n1542) );
  OR2_X1 U1195 ( .A1(n1796), .A2(n1797), .ZN(n1543) );
  AND2_X1 U1196 ( .A1(n2070), .A2(n2068), .ZN(n1544) );
  AND2_X1 U1197 ( .A1(n2014), .A2(n2016), .ZN(n1545) );
  AND2_X1 U1198 ( .A1(n1849), .A2(n1851), .ZN(n1546) );
  OR2_X1 U1199 ( .A1(n2070), .A2(n2069), .ZN(n1547) );
  OR2_X1 U1200 ( .A1(n2014), .A2(n2015), .ZN(n1548) );
  OR2_X1 U1201 ( .A1(n1959), .A2(n1960), .ZN(n1549) );
  OR2_X1 U1202 ( .A1(n1904), .A2(n1905), .ZN(n1550) );
  OR2_X1 U1203 ( .A1(n1794), .A2(n1795), .ZN(n1551) );
  AND2_X1 U1204 ( .A1(n1959), .A2(n1961), .ZN(n1552) );
  AND2_X1 U1205 ( .A1(n1904), .A2(n1906), .ZN(n1553) );
  AND2_X1 U1206 ( .A1(n1794), .A2(n1796), .ZN(n1554) );
  BUF_X1 U1207 ( .A(n1647), .Z(n1567) );
  INV_X1 U1208 ( .A(n1599), .ZN(n1598) );
  AND2_X1 U1209 ( .A1(a[0]), .A2(n2157), .ZN(n1555) );
  BUF_X1 U1210 ( .A(a[20]), .Z(n1600) );
  INV_X1 U1211 ( .A(a[23]), .ZN(n1599) );
  INV_X1 U1212 ( .A(a[5]), .ZN(n1611) );
  INV_X1 U1213 ( .A(a[11]), .ZN(n1607) );
  INV_X1 U1214 ( .A(a[8]), .ZN(n1609) );
  INV_X1 U1215 ( .A(a[17]), .ZN(n1603) );
  INV_X1 U1216 ( .A(a[14]), .ZN(n1605) );
  BUF_X1 U1217 ( .A(a[20]), .Z(n1601) );
  CLKBUF_X1 U1218 ( .A(b[23]), .Z(n1612) );
  CLKBUF_X1 U1219 ( .A(b[23]), .Z(n1613) );
  INV_X1 U1220 ( .A(b[23]), .ZN(n1615) );
  INV_X1 U1221 ( .A(n1612), .ZN(n1616) );
  INV_X1 U1222 ( .A(n1612), .ZN(n1617) );
  INV_X1 U1223 ( .A(n1612), .ZN(n1618) );
  INV_X1 U1224 ( .A(n1613), .ZN(n1619) );
  INV_X1 U1225 ( .A(n1613), .ZN(n1620) );
  AOI21_X1 U1226 ( .B1(n1621), .B2(n1622), .A(n1623), .ZN(product[47]) );
  OAI22_X1 U1227 ( .A1(n1624), .A2(n1625), .B1(n1624), .B2(n1626), .ZN(n1623)
         );
  INV_X1 U1228 ( .A(n1622), .ZN(n1626) );
  AOI222_X1 U1229 ( .A1(n1627), .A2(n303), .B1(n1625), .B2(n303), .C1(n1627), 
        .C2(n1625), .ZN(n1624) );
  XOR2_X1 U1230 ( .A(n1628), .B(n1599), .Z(n1622) );
  OAI221_X1 U1231 ( .B1(n1617), .B2(n1557), .C1(n1620), .C2(n1558), .A(n1630), 
        .ZN(n1628) );
  OAI21_X1 U1232 ( .B1(n1559), .B2(n1560), .A(n1614), .ZN(n1630) );
  INV_X1 U1233 ( .A(n1625), .ZN(n1621) );
  XOR2_X1 U1234 ( .A(a[23]), .B(n1631), .Z(n1625) );
  AOI221_X1 U1235 ( .B1(n1613), .B2(n1559), .C1(n1560), .C2(n1614), .A(n1632), 
        .ZN(n1631) );
  OAI22_X1 U1236 ( .A1(n1558), .A2(n1633), .B1(n1557), .B2(n1634), .ZN(n1632)
         );
  XNOR2_X1 U1237 ( .A(a[2]), .B(n1635), .ZN(n908) );
  AOI221_X1 U1238 ( .B1(n1561), .B2(b[22]), .C1(n1563), .C2(b[21]), .A(n1637), 
        .ZN(n1635) );
  OAI22_X1 U1239 ( .A1(n1564), .A2(n1638), .B1(n1639), .B2(n1640), .ZN(n1637)
         );
  INV_X1 U1240 ( .A(n1376), .ZN(n1638) );
  XNOR2_X1 U1241 ( .A(a[2]), .B(n1641), .ZN(n907) );
  AOI221_X1 U1242 ( .B1(n1563), .B2(b[22]), .C1(n1555), .C2(n1375), .A(n1642), 
        .ZN(n1641) );
  OAI22_X1 U1243 ( .A1(n1643), .A2(n1639), .B1(n1617), .B2(n1535), .ZN(n1642)
         );
  XNOR2_X1 U1244 ( .A(a[2]), .B(n1644), .ZN(n906) );
  AOI221_X1 U1245 ( .B1(n1561), .B2(n1613), .C1(n1563), .C2(n1614), .A(n1645), 
        .ZN(n1644) );
  OAI22_X1 U1246 ( .A1(n1633), .A2(n1564), .B1(n1634), .B2(n1639), .ZN(n1645)
         );
  XNOR2_X1 U1247 ( .A(n1646), .B(n1611), .ZN(n904) );
  OAI22_X1 U1248 ( .A1(n1565), .A2(n1534), .B1(n1568), .B2(n1567), .ZN(n1646)
         );
  XNOR2_X1 U1249 ( .A(n1648), .B(n1611), .ZN(n903) );
  OAI222_X1 U1250 ( .A1(n1534), .A2(n1649), .B1(n1566), .B2(n1533), .C1(n1568), 
        .C2(n1650), .ZN(n1648) );
  XNOR2_X1 U1251 ( .A(n1610), .B(n1651), .ZN(n902) );
  AOI221_X1 U1252 ( .B1(b[2]), .B2(n1569), .C1(b[1]), .C2(n1570), .A(n1652), 
        .ZN(n1651) );
  OAI22_X1 U1253 ( .A1(n1568), .A2(n1653), .B1(n1565), .B2(n1572), .ZN(n1652)
         );
  XNOR2_X1 U1254 ( .A(n1610), .B(n1655), .ZN(n901) );
  AOI221_X1 U1255 ( .B1(b[3]), .B2(n1569), .C1(b[2]), .C2(n1570), .A(n1656), 
        .ZN(n1655) );
  OAI22_X1 U1256 ( .A1(n1568), .A2(n1657), .B1(n1649), .B2(n1572), .ZN(n1656)
         );
  XNOR2_X1 U1257 ( .A(n1610), .B(n1658), .ZN(n900) );
  AOI221_X1 U1258 ( .B1(b[4]), .B2(n1569), .C1(b[3]), .C2(n1570), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1259 ( .A1(n1568), .A2(n1660), .B1(n1661), .B2(n1572), .ZN(n1659)
         );
  XNOR2_X1 U1260 ( .A(n1610), .B(n1662), .ZN(n899) );
  AOI221_X1 U1261 ( .B1(b[5]), .B2(n1569), .C1(b[4]), .C2(n1570), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1262 ( .A1(n1568), .A2(n1664), .B1(n1572), .B2(n1665), .ZN(n1663)
         );
  XNOR2_X1 U1263 ( .A(n1610), .B(n1666), .ZN(n898) );
  AOI221_X1 U1264 ( .B1(b[6]), .B2(n1569), .C1(b[5]), .C2(n1570), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1265 ( .A1(n1568), .A2(n1668), .B1(n1572), .B2(n1669), .ZN(n1667)
         );
  XNOR2_X1 U1266 ( .A(n1610), .B(n1670), .ZN(n897) );
  AOI221_X1 U1267 ( .B1(b[7]), .B2(n1569), .C1(b[6]), .C2(n1570), .A(n1671), 
        .ZN(n1670) );
  OAI22_X1 U1268 ( .A1(n1568), .A2(n1672), .B1(n1572), .B2(n1673), .ZN(n1671)
         );
  XNOR2_X1 U1269 ( .A(n1610), .B(n1674), .ZN(n896) );
  AOI221_X1 U1270 ( .B1(b[8]), .B2(n1569), .C1(b[7]), .C2(n1570), .A(n1675), 
        .ZN(n1674) );
  OAI22_X1 U1271 ( .A1(n1568), .A2(n1676), .B1(n1571), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1272 ( .A(n1610), .B(n1678), .ZN(n895) );
  AOI221_X1 U1273 ( .B1(b[9]), .B2(n1569), .C1(b[8]), .C2(n1570), .A(n1679), 
        .ZN(n1678) );
  OAI22_X1 U1274 ( .A1(n1568), .A2(n1680), .B1(n1572), .B2(n1681), .ZN(n1679)
         );
  XNOR2_X1 U1275 ( .A(n1610), .B(n1682), .ZN(n894) );
  AOI221_X1 U1276 ( .B1(b[10]), .B2(n1569), .C1(b[9]), .C2(n1570), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1277 ( .A1(n1568), .A2(n1684), .B1(n1572), .B2(n1685), .ZN(n1683)
         );
  XNOR2_X1 U1278 ( .A(n1610), .B(n1686), .ZN(n893) );
  AOI221_X1 U1279 ( .B1(b[11]), .B2(n1569), .C1(b[10]), .C2(n1570), .A(n1687), 
        .ZN(n1686) );
  OAI22_X1 U1280 ( .A1(n1568), .A2(n1688), .B1(n1571), .B2(n1689), .ZN(n1687)
         );
  XNOR2_X1 U1281 ( .A(n1610), .B(n1690), .ZN(n892) );
  AOI221_X1 U1282 ( .B1(b[12]), .B2(n1569), .C1(b[11]), .C2(n1570), .A(n1691), 
        .ZN(n1690) );
  OAI22_X1 U1283 ( .A1(n1568), .A2(n1692), .B1(n1571), .B2(n1693), .ZN(n1691)
         );
  XNOR2_X1 U1284 ( .A(n1610), .B(n1694), .ZN(n891) );
  AOI221_X1 U1285 ( .B1(b[13]), .B2(n1569), .C1(b[12]), .C2(n1570), .A(n1695), 
        .ZN(n1694) );
  OAI22_X1 U1286 ( .A1(n1568), .A2(n1696), .B1(n1571), .B2(n1697), .ZN(n1695)
         );
  XNOR2_X1 U1287 ( .A(n1610), .B(n1698), .ZN(n890) );
  AOI221_X1 U1288 ( .B1(b[14]), .B2(n1569), .C1(b[13]), .C2(n1570), .A(n1699), 
        .ZN(n1698) );
  OAI22_X1 U1289 ( .A1(n1568), .A2(n1700), .B1(n1571), .B2(n1701), .ZN(n1699)
         );
  XNOR2_X1 U1290 ( .A(n1610), .B(n1702), .ZN(n889) );
  AOI221_X1 U1291 ( .B1(b[15]), .B2(n1569), .C1(b[14]), .C2(n1570), .A(n1703), 
        .ZN(n1702) );
  OAI22_X1 U1292 ( .A1(n1568), .A2(n1704), .B1(n1571), .B2(n1705), .ZN(n1703)
         );
  XNOR2_X1 U1293 ( .A(n1610), .B(n1706), .ZN(n888) );
  AOI221_X1 U1294 ( .B1(b[16]), .B2(n1569), .C1(b[15]), .C2(n1570), .A(n1707), 
        .ZN(n1706) );
  OAI22_X1 U1295 ( .A1(n1568), .A2(n1708), .B1(n1571), .B2(n1709), .ZN(n1707)
         );
  XNOR2_X1 U1296 ( .A(n1610), .B(n1710), .ZN(n887) );
  AOI221_X1 U1297 ( .B1(b[17]), .B2(n1569), .C1(b[16]), .C2(n1570), .A(n1711), 
        .ZN(n1710) );
  OAI22_X1 U1298 ( .A1(n1568), .A2(n1712), .B1(n1571), .B2(n1713), .ZN(n1711)
         );
  XNOR2_X1 U1299 ( .A(n1610), .B(n1714), .ZN(n886) );
  AOI221_X1 U1300 ( .B1(b[18]), .B2(n1569), .C1(b[17]), .C2(n1570), .A(n1715), 
        .ZN(n1714) );
  OAI22_X1 U1301 ( .A1(n1568), .A2(n1716), .B1(n1571), .B2(n1717), .ZN(n1715)
         );
  XNOR2_X1 U1302 ( .A(n1610), .B(n1718), .ZN(n885) );
  AOI221_X1 U1303 ( .B1(b[19]), .B2(n1569), .C1(b[18]), .C2(n1570), .A(n1719), 
        .ZN(n1718) );
  OAI22_X1 U1304 ( .A1(n1568), .A2(n1720), .B1(n1571), .B2(n1721), .ZN(n1719)
         );
  XNOR2_X1 U1305 ( .A(a[5]), .B(n1722), .ZN(n884) );
  AOI221_X1 U1306 ( .B1(n1569), .B2(b[20]), .C1(b[19]), .C2(n1570), .A(n1723), 
        .ZN(n1722) );
  OAI22_X1 U1307 ( .A1(n1568), .A2(n1724), .B1(n1571), .B2(n1725), .ZN(n1723)
         );
  XNOR2_X1 U1308 ( .A(a[5]), .B(n1726), .ZN(n883) );
  AOI221_X1 U1309 ( .B1(n1569), .B2(b[21]), .C1(n1570), .C2(b[20]), .A(n1727), 
        .ZN(n1726) );
  OAI22_X1 U1310 ( .A1(n1568), .A2(n1728), .B1(n1571), .B2(n1729), .ZN(n1727)
         );
  XNOR2_X1 U1311 ( .A(a[5]), .B(n1730), .ZN(n882) );
  AOI221_X1 U1312 ( .B1(n1569), .B2(b[22]), .C1(n1536), .C2(n1376), .A(n1731), 
        .ZN(n1730) );
  OAI22_X1 U1313 ( .A1(n1640), .A2(n1572), .B1(n1643), .B2(n1533), .ZN(n1731)
         );
  XNOR2_X1 U1314 ( .A(a[5]), .B(n1732), .ZN(n881) );
  AOI221_X1 U1315 ( .B1(n1570), .B2(b[22]), .C1(n1536), .C2(n1375), .A(n1733), 
        .ZN(n1732) );
  OAI22_X1 U1316 ( .A1(n1615), .A2(n1534), .B1(n1643), .B2(n1572), .ZN(n1733)
         );
  XNOR2_X1 U1317 ( .A(a[5]), .B(n1734), .ZN(n880) );
  AOI221_X1 U1318 ( .B1(n1569), .B2(n1613), .C1(n1570), .C2(n1614), .A(n1735), 
        .ZN(n1734) );
  OAI22_X1 U1319 ( .A1(n1633), .A2(n1568), .B1(n1634), .B2(n1572), .ZN(n1735)
         );
  XNOR2_X1 U1320 ( .A(n1610), .B(n1736), .ZN(n879) );
  OAI221_X1 U1321 ( .B1(n1616), .B2(n1572), .C1(n1620), .C2(n1568), .A(n1737), 
        .ZN(n1736) );
  OAI21_X1 U1322 ( .B1(n1569), .B2(n1570), .A(n1614), .ZN(n1737) );
  INV_X1 U1323 ( .A(n1741), .ZN(n1738) );
  NAND3_X1 U1324 ( .A1(n1741), .A2(n1740), .A3(n1739), .ZN(n1654) );
  XNOR2_X1 U1325 ( .A(a[3]), .B(a[4]), .ZN(n1739) );
  XNOR2_X1 U1326 ( .A(a[4]), .B(n1611), .ZN(n1740) );
  XOR2_X1 U1327 ( .A(a[3]), .B(n1742), .Z(n1741) );
  XNOR2_X1 U1328 ( .A(n1743), .B(n1609), .ZN(n878) );
  OAI22_X1 U1329 ( .A1(n1565), .A2(n1543), .B1(n1565), .B2(n1573), .ZN(n1743)
         );
  XNOR2_X1 U1330 ( .A(n1744), .B(n1609), .ZN(n877) );
  OAI222_X1 U1331 ( .A1(n1649), .A2(n1543), .B1(n1566), .B2(n1551), .C1(n1650), 
        .C2(n1573), .ZN(n1744) );
  XNOR2_X1 U1332 ( .A(n1608), .B(n1745), .ZN(n876) );
  AOI221_X1 U1333 ( .B1(n1574), .B2(b[2]), .C1(n1575), .C2(b[1]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1334 ( .A1(n1653), .A2(n1573), .B1(n1565), .B2(n1576), .ZN(n1746)
         );
  XNOR2_X1 U1335 ( .A(n1608), .B(n1748), .ZN(n875) );
  AOI221_X1 U1336 ( .B1(n1574), .B2(b[3]), .C1(n1575), .C2(b[2]), .A(n1749), 
        .ZN(n1748) );
  OAI22_X1 U1337 ( .A1(n1657), .A2(n1573), .B1(n1649), .B2(n1577), .ZN(n1749)
         );
  XNOR2_X1 U1338 ( .A(n1608), .B(n1750), .ZN(n874) );
  AOI221_X1 U1339 ( .B1(n1574), .B2(b[4]), .C1(n1575), .C2(b[3]), .A(n1751), 
        .ZN(n1750) );
  OAI22_X1 U1340 ( .A1(n1660), .A2(n1573), .B1(n1661), .B2(n1577), .ZN(n1751)
         );
  XNOR2_X1 U1341 ( .A(n1608), .B(n1752), .ZN(n873) );
  AOI221_X1 U1342 ( .B1(n1574), .B2(b[5]), .C1(n1575), .C2(b[4]), .A(n1753), 
        .ZN(n1752) );
  OAI22_X1 U1343 ( .A1(n1664), .A2(n1573), .B1(n1665), .B2(n1577), .ZN(n1753)
         );
  XNOR2_X1 U1344 ( .A(n1608), .B(n1754), .ZN(n872) );
  AOI221_X1 U1345 ( .B1(n1574), .B2(b[6]), .C1(n1575), .C2(b[5]), .A(n1755), 
        .ZN(n1754) );
  OAI22_X1 U1346 ( .A1(n1668), .A2(n1573), .B1(n1669), .B2(n1577), .ZN(n1755)
         );
  XNOR2_X1 U1347 ( .A(n1608), .B(n1756), .ZN(n871) );
  AOI221_X1 U1348 ( .B1(n1574), .B2(b[7]), .C1(n1575), .C2(b[6]), .A(n1757), 
        .ZN(n1756) );
  OAI22_X1 U1349 ( .A1(n1672), .A2(n1573), .B1(n1673), .B2(n1577), .ZN(n1757)
         );
  XNOR2_X1 U1350 ( .A(n1608), .B(n1758), .ZN(n870) );
  AOI221_X1 U1351 ( .B1(n1574), .B2(b[8]), .C1(n1575), .C2(b[7]), .A(n1759), 
        .ZN(n1758) );
  OAI22_X1 U1352 ( .A1(n1676), .A2(n1573), .B1(n1677), .B2(n1577), .ZN(n1759)
         );
  XNOR2_X1 U1353 ( .A(n1608), .B(n1760), .ZN(n869) );
  AOI221_X1 U1354 ( .B1(n1574), .B2(b[9]), .C1(n1575), .C2(b[8]), .A(n1761), 
        .ZN(n1760) );
  OAI22_X1 U1355 ( .A1(n1680), .A2(n1573), .B1(n1681), .B2(n1577), .ZN(n1761)
         );
  XNOR2_X1 U1356 ( .A(n1608), .B(n1762), .ZN(n868) );
  AOI221_X1 U1357 ( .B1(n1574), .B2(b[10]), .C1(n1575), .C2(b[9]), .A(n1763), 
        .ZN(n1762) );
  OAI22_X1 U1358 ( .A1(n1684), .A2(n1573), .B1(n1685), .B2(n1577), .ZN(n1763)
         );
  XNOR2_X1 U1359 ( .A(n1608), .B(n1764), .ZN(n867) );
  AOI221_X1 U1360 ( .B1(n1574), .B2(b[11]), .C1(n1575), .C2(b[10]), .A(n1765), 
        .ZN(n1764) );
  OAI22_X1 U1361 ( .A1(n1688), .A2(n1573), .B1(n1689), .B2(n1577), .ZN(n1765)
         );
  XNOR2_X1 U1362 ( .A(n1608), .B(n1766), .ZN(n866) );
  AOI221_X1 U1363 ( .B1(n1574), .B2(b[12]), .C1(n1575), .C2(b[11]), .A(n1767), 
        .ZN(n1766) );
  OAI22_X1 U1364 ( .A1(n1692), .A2(n1573), .B1(n1693), .B2(n1577), .ZN(n1767)
         );
  XNOR2_X1 U1365 ( .A(n1608), .B(n1768), .ZN(n865) );
  AOI221_X1 U1366 ( .B1(n1574), .B2(b[13]), .C1(n1575), .C2(b[12]), .A(n1769), 
        .ZN(n1768) );
  OAI22_X1 U1367 ( .A1(n1696), .A2(n1573), .B1(n1697), .B2(n1576), .ZN(n1769)
         );
  XNOR2_X1 U1368 ( .A(n1608), .B(n1770), .ZN(n864) );
  AOI221_X1 U1369 ( .B1(n1574), .B2(b[14]), .C1(n1575), .C2(b[13]), .A(n1771), 
        .ZN(n1770) );
  OAI22_X1 U1370 ( .A1(n1700), .A2(n1573), .B1(n1701), .B2(n1576), .ZN(n1771)
         );
  XNOR2_X1 U1371 ( .A(n1608), .B(n1772), .ZN(n863) );
  AOI221_X1 U1372 ( .B1(n1574), .B2(b[15]), .C1(n1575), .C2(b[14]), .A(n1773), 
        .ZN(n1772) );
  OAI22_X1 U1373 ( .A1(n1704), .A2(n1573), .B1(n1705), .B2(n1576), .ZN(n1773)
         );
  XNOR2_X1 U1374 ( .A(n1608), .B(n1774), .ZN(n862) );
  AOI221_X1 U1375 ( .B1(n1574), .B2(b[16]), .C1(n1575), .C2(b[15]), .A(n1775), 
        .ZN(n1774) );
  OAI22_X1 U1376 ( .A1(n1708), .A2(n1573), .B1(n1709), .B2(n1576), .ZN(n1775)
         );
  XNOR2_X1 U1377 ( .A(n1608), .B(n1776), .ZN(n861) );
  AOI221_X1 U1378 ( .B1(n1574), .B2(b[17]), .C1(n1575), .C2(b[16]), .A(n1777), 
        .ZN(n1776) );
  OAI22_X1 U1379 ( .A1(n1712), .A2(n1573), .B1(n1713), .B2(n1576), .ZN(n1777)
         );
  XNOR2_X1 U1380 ( .A(n1608), .B(n1778), .ZN(n860) );
  AOI221_X1 U1381 ( .B1(n1574), .B2(b[18]), .C1(n1575), .C2(b[17]), .A(n1779), 
        .ZN(n1778) );
  OAI22_X1 U1382 ( .A1(n1716), .A2(n1573), .B1(n1717), .B2(n1576), .ZN(n1779)
         );
  XNOR2_X1 U1383 ( .A(n1608), .B(n1780), .ZN(n859) );
  AOI221_X1 U1384 ( .B1(n1574), .B2(b[19]), .C1(n1575), .C2(b[18]), .A(n1781), 
        .ZN(n1780) );
  OAI22_X1 U1385 ( .A1(n1720), .A2(n1573), .B1(n1721), .B2(n1576), .ZN(n1781)
         );
  XNOR2_X1 U1386 ( .A(a[8]), .B(n1782), .ZN(n858) );
  AOI221_X1 U1387 ( .B1(n1574), .B2(b[20]), .C1(n1575), .C2(b[19]), .A(n1783), 
        .ZN(n1782) );
  OAI22_X1 U1388 ( .A1(n1724), .A2(n1573), .B1(n1725), .B2(n1576), .ZN(n1783)
         );
  XNOR2_X1 U1389 ( .A(a[8]), .B(n1784), .ZN(n857) );
  AOI221_X1 U1390 ( .B1(n1574), .B2(b[21]), .C1(n1575), .C2(b[20]), .A(n1785), 
        .ZN(n1784) );
  OAI22_X1 U1391 ( .A1(n1728), .A2(n1573), .B1(n1729), .B2(n1576), .ZN(n1785)
         );
  XNOR2_X1 U1392 ( .A(a[8]), .B(n1786), .ZN(n856) );
  AOI221_X1 U1393 ( .B1(n1574), .B2(b[22]), .C1(n1554), .C2(n1376), .A(n1787), 
        .ZN(n1786) );
  OAI22_X1 U1394 ( .A1(n1640), .A2(n1577), .B1(n1643), .B2(n1551), .ZN(n1787)
         );
  XNOR2_X1 U1395 ( .A(a[8]), .B(n1788), .ZN(n855) );
  AOI221_X1 U1396 ( .B1(n1575), .B2(b[22]), .C1(n1554), .C2(n1375), .A(n1789), 
        .ZN(n1788) );
  OAI22_X1 U1397 ( .A1(n1617), .A2(n1543), .B1(n1643), .B2(n1576), .ZN(n1789)
         );
  XNOR2_X1 U1398 ( .A(a[8]), .B(n1790), .ZN(n854) );
  AOI221_X1 U1399 ( .B1(n1574), .B2(n1613), .C1(n1575), .C2(n1614), .A(n1791), 
        .ZN(n1790) );
  OAI22_X1 U1400 ( .A1(n1633), .A2(n1573), .B1(n1634), .B2(n1576), .ZN(n1791)
         );
  XNOR2_X1 U1401 ( .A(n1608), .B(n1792), .ZN(n853) );
  OAI221_X1 U1402 ( .B1(n1616), .B2(n1577), .C1(n1617), .C2(n1573), .A(n1793), 
        .ZN(n1792) );
  OAI21_X1 U1403 ( .B1(n1574), .B2(n1575), .A(n1614), .ZN(n1793) );
  INV_X1 U1404 ( .A(n1797), .ZN(n1794) );
  NAND3_X1 U1405 ( .A1(n1797), .A2(n1796), .A3(n1795), .ZN(n1747) );
  XNOR2_X1 U1406 ( .A(a[6]), .B(a[7]), .ZN(n1795) );
  XNOR2_X1 U1407 ( .A(a[7]), .B(n1609), .ZN(n1796) );
  XOR2_X1 U1408 ( .A(a[6]), .B(n1611), .Z(n1797) );
  XNOR2_X1 U1409 ( .A(n1798), .B(n1607), .ZN(n852) );
  OAI22_X1 U1410 ( .A1(n1565), .A2(n1542), .B1(n1565), .B2(n1578), .ZN(n1798)
         );
  XNOR2_X1 U1411 ( .A(n1799), .B(n1607), .ZN(n851) );
  OAI222_X1 U1412 ( .A1(n1649), .A2(n1542), .B1(n1566), .B2(n1537), .C1(n1650), 
        .C2(n1578), .ZN(n1799) );
  XNOR2_X1 U1413 ( .A(n1606), .B(n1800), .ZN(n850) );
  AOI221_X1 U1414 ( .B1(n1579), .B2(b[2]), .C1(n1580), .C2(b[1]), .A(n1801), 
        .ZN(n1800) );
  OAI22_X1 U1415 ( .A1(n1653), .A2(n1578), .B1(n1566), .B2(n1581), .ZN(n1801)
         );
  XNOR2_X1 U1416 ( .A(n1606), .B(n1803), .ZN(n849) );
  AOI221_X1 U1417 ( .B1(n1579), .B2(b[3]), .C1(n1580), .C2(b[2]), .A(n1804), 
        .ZN(n1803) );
  OAI22_X1 U1418 ( .A1(n1657), .A2(n1578), .B1(n1649), .B2(n1582), .ZN(n1804)
         );
  XNOR2_X1 U1419 ( .A(n1606), .B(n1805), .ZN(n848) );
  AOI221_X1 U1420 ( .B1(n1579), .B2(b[4]), .C1(n1580), .C2(b[3]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1421 ( .A1(n1660), .A2(n1578), .B1(n1661), .B2(n1582), .ZN(n1806)
         );
  XNOR2_X1 U1422 ( .A(n1606), .B(n1807), .ZN(n847) );
  AOI221_X1 U1423 ( .B1(n1579), .B2(b[5]), .C1(n1580), .C2(b[4]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1424 ( .A1(n1664), .A2(n1578), .B1(n1665), .B2(n1582), .ZN(n1808)
         );
  XNOR2_X1 U1425 ( .A(n1606), .B(n1809), .ZN(n846) );
  AOI221_X1 U1426 ( .B1(n1579), .B2(b[6]), .C1(n1580), .C2(b[5]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1427 ( .A1(n1668), .A2(n1578), .B1(n1669), .B2(n1582), .ZN(n1810)
         );
  XNOR2_X1 U1428 ( .A(n1606), .B(n1811), .ZN(n845) );
  AOI221_X1 U1429 ( .B1(n1579), .B2(b[7]), .C1(n1580), .C2(b[6]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1430 ( .A1(n1672), .A2(n1578), .B1(n1673), .B2(n1582), .ZN(n1812)
         );
  XNOR2_X1 U1431 ( .A(n1606), .B(n1813), .ZN(n844) );
  AOI221_X1 U1432 ( .B1(n1579), .B2(b[8]), .C1(n1580), .C2(b[7]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1433 ( .A1(n1676), .A2(n1578), .B1(n1677), .B2(n1582), .ZN(n1814)
         );
  XNOR2_X1 U1434 ( .A(n1606), .B(n1815), .ZN(n843) );
  AOI221_X1 U1435 ( .B1(n1579), .B2(b[9]), .C1(n1580), .C2(b[8]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1436 ( .A1(n1680), .A2(n1578), .B1(n1681), .B2(n1582), .ZN(n1816)
         );
  XNOR2_X1 U1437 ( .A(n1606), .B(n1817), .ZN(n842) );
  AOI221_X1 U1438 ( .B1(n1579), .B2(b[10]), .C1(n1580), .C2(b[9]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1439 ( .A1(n1684), .A2(n1578), .B1(n1685), .B2(n1582), .ZN(n1818)
         );
  XNOR2_X1 U1440 ( .A(n1606), .B(n1819), .ZN(n841) );
  AOI221_X1 U1441 ( .B1(n1579), .B2(b[11]), .C1(n1580), .C2(b[10]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1442 ( .A1(n1688), .A2(n1578), .B1(n1689), .B2(n1582), .ZN(n1820)
         );
  XNOR2_X1 U1443 ( .A(n1606), .B(n1821), .ZN(n840) );
  AOI221_X1 U1444 ( .B1(n1579), .B2(b[12]), .C1(n1580), .C2(b[11]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1445 ( .A1(n1692), .A2(n1578), .B1(n1693), .B2(n1582), .ZN(n1822)
         );
  XNOR2_X1 U1446 ( .A(n1606), .B(n1823), .ZN(n839) );
  AOI221_X1 U1447 ( .B1(n1579), .B2(b[13]), .C1(n1580), .C2(b[12]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1448 ( .A1(n1696), .A2(n1578), .B1(n1697), .B2(n1581), .ZN(n1824)
         );
  XNOR2_X1 U1449 ( .A(n1606), .B(n1825), .ZN(n838) );
  AOI221_X1 U1450 ( .B1(n1579), .B2(b[14]), .C1(n1580), .C2(b[13]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1451 ( .A1(n1700), .A2(n1578), .B1(n1701), .B2(n1581), .ZN(n1826)
         );
  XNOR2_X1 U1452 ( .A(n1606), .B(n1827), .ZN(n837) );
  AOI221_X1 U1453 ( .B1(n1579), .B2(b[15]), .C1(n1580), .C2(b[14]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1454 ( .A1(n1704), .A2(n1578), .B1(n1705), .B2(n1581), .ZN(n1828)
         );
  XNOR2_X1 U1455 ( .A(n1606), .B(n1829), .ZN(n836) );
  AOI221_X1 U1456 ( .B1(n1579), .B2(b[16]), .C1(n1580), .C2(b[15]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1457 ( .A1(n1708), .A2(n1578), .B1(n1709), .B2(n1581), .ZN(n1830)
         );
  XNOR2_X1 U1458 ( .A(n1606), .B(n1831), .ZN(n835) );
  AOI221_X1 U1459 ( .B1(n1579), .B2(b[17]), .C1(n1580), .C2(b[16]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1460 ( .A1(n1712), .A2(n1578), .B1(n1713), .B2(n1581), .ZN(n1832)
         );
  XNOR2_X1 U1461 ( .A(n1606), .B(n1833), .ZN(n834) );
  AOI221_X1 U1462 ( .B1(n1579), .B2(b[18]), .C1(n1580), .C2(b[17]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1463 ( .A1(n1716), .A2(n1578), .B1(n1717), .B2(n1581), .ZN(n1834)
         );
  XNOR2_X1 U1464 ( .A(n1606), .B(n1835), .ZN(n833) );
  AOI221_X1 U1465 ( .B1(n1579), .B2(b[19]), .C1(n1580), .C2(b[18]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1466 ( .A1(n1720), .A2(n1578), .B1(n1721), .B2(n1581), .ZN(n1836)
         );
  XNOR2_X1 U1467 ( .A(n1606), .B(n1837), .ZN(n832) );
  AOI221_X1 U1468 ( .B1(n1579), .B2(b[20]), .C1(n1580), .C2(b[19]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1469 ( .A1(n1724), .A2(n1578), .B1(n1725), .B2(n1581), .ZN(n1838)
         );
  XNOR2_X1 U1470 ( .A(a[11]), .B(n1839), .ZN(n831) );
  AOI221_X1 U1471 ( .B1(n1579), .B2(b[21]), .C1(n1580), .C2(b[20]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1472 ( .A1(n1728), .A2(n1578), .B1(n1729), .B2(n1581), .ZN(n1840)
         );
  XNOR2_X1 U1473 ( .A(a[11]), .B(n1841), .ZN(n830) );
  AOI221_X1 U1474 ( .B1(n1579), .B2(b[22]), .C1(n1546), .C2(n1376), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1475 ( .A1(n1640), .A2(n1582), .B1(n1643), .B2(n1537), .ZN(n1842)
         );
  XNOR2_X1 U1476 ( .A(a[11]), .B(n1843), .ZN(n829) );
  AOI221_X1 U1477 ( .B1(n1580), .B2(b[22]), .C1(n1546), .C2(n1375), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1478 ( .A1(n1617), .A2(n1542), .B1(n1643), .B2(n1581), .ZN(n1844)
         );
  XNOR2_X1 U1479 ( .A(a[11]), .B(n1845), .ZN(n828) );
  AOI221_X1 U1480 ( .B1(n1579), .B2(n1614), .C1(n1580), .C2(n1614), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1481 ( .A1(n1633), .A2(n1578), .B1(n1634), .B2(n1581), .ZN(n1846)
         );
  XNOR2_X1 U1482 ( .A(a[11]), .B(n1847), .ZN(n827) );
  OAI221_X1 U1483 ( .B1(n1616), .B2(n1582), .C1(n1617), .C2(n1578), .A(n1848), 
        .ZN(n1847) );
  OAI21_X1 U1484 ( .B1(n1579), .B2(n1580), .A(n1614), .ZN(n1848) );
  INV_X1 U1485 ( .A(n1852), .ZN(n1849) );
  NAND3_X1 U1486 ( .A1(n1852), .A2(n1851), .A3(n1850), .ZN(n1802) );
  XNOR2_X1 U1487 ( .A(a[10]), .B(a[9]), .ZN(n1850) );
  XNOR2_X1 U1488 ( .A(a[10]), .B(n1607), .ZN(n1851) );
  XOR2_X1 U1489 ( .A(a[9]), .B(n1609), .Z(n1852) );
  XNOR2_X1 U1490 ( .A(n1853), .B(n1605), .ZN(n826) );
  OAI22_X1 U1491 ( .A1(n1565), .A2(n1541), .B1(n1565), .B2(n1583), .ZN(n1853)
         );
  XNOR2_X1 U1492 ( .A(n1854), .B(n1605), .ZN(n825) );
  OAI222_X1 U1493 ( .A1(n1649), .A2(n1541), .B1(n1566), .B2(n1550), .C1(n1650), 
        .C2(n1583), .ZN(n1854) );
  XNOR2_X1 U1494 ( .A(n1604), .B(n1855), .ZN(n824) );
  AOI221_X1 U1495 ( .B1(n1584), .B2(b[2]), .C1(n1585), .C2(b[1]), .A(n1856), 
        .ZN(n1855) );
  OAI22_X1 U1496 ( .A1(n1653), .A2(n1583), .B1(n1565), .B2(n1586), .ZN(n1856)
         );
  XNOR2_X1 U1497 ( .A(n1604), .B(n1858), .ZN(n823) );
  AOI221_X1 U1498 ( .B1(n1584), .B2(b[3]), .C1(n1585), .C2(b[2]), .A(n1859), 
        .ZN(n1858) );
  OAI22_X1 U1499 ( .A1(n1657), .A2(n1583), .B1(n1649), .B2(n1587), .ZN(n1859)
         );
  XNOR2_X1 U1500 ( .A(n1604), .B(n1860), .ZN(n822) );
  AOI221_X1 U1501 ( .B1(n1584), .B2(b[4]), .C1(n1585), .C2(b[3]), .A(n1861), 
        .ZN(n1860) );
  OAI22_X1 U1502 ( .A1(n1660), .A2(n1583), .B1(n1661), .B2(n1587), .ZN(n1861)
         );
  XNOR2_X1 U1503 ( .A(n1604), .B(n1862), .ZN(n821) );
  AOI221_X1 U1504 ( .B1(n1584), .B2(b[5]), .C1(n1585), .C2(b[4]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1505 ( .A1(n1664), .A2(n1583), .B1(n1665), .B2(n1587), .ZN(n1863)
         );
  XNOR2_X1 U1506 ( .A(n1604), .B(n1864), .ZN(n820) );
  AOI221_X1 U1507 ( .B1(n1584), .B2(b[6]), .C1(n1585), .C2(b[5]), .A(n1865), 
        .ZN(n1864) );
  OAI22_X1 U1508 ( .A1(n1668), .A2(n1583), .B1(n1669), .B2(n1587), .ZN(n1865)
         );
  XNOR2_X1 U1509 ( .A(n1604), .B(n1866), .ZN(n819) );
  AOI221_X1 U1510 ( .B1(n1584), .B2(b[7]), .C1(n1585), .C2(b[6]), .A(n1867), 
        .ZN(n1866) );
  OAI22_X1 U1511 ( .A1(n1672), .A2(n1583), .B1(n1673), .B2(n1587), .ZN(n1867)
         );
  XNOR2_X1 U1512 ( .A(n1604), .B(n1868), .ZN(n818) );
  AOI221_X1 U1513 ( .B1(n1584), .B2(b[8]), .C1(n1585), .C2(b[7]), .A(n1869), 
        .ZN(n1868) );
  OAI22_X1 U1514 ( .A1(n1676), .A2(n1583), .B1(n1677), .B2(n1587), .ZN(n1869)
         );
  XNOR2_X1 U1515 ( .A(n1604), .B(n1870), .ZN(n817) );
  AOI221_X1 U1516 ( .B1(n1584), .B2(b[9]), .C1(n1585), .C2(b[8]), .A(n1871), 
        .ZN(n1870) );
  OAI22_X1 U1517 ( .A1(n1680), .A2(n1583), .B1(n1681), .B2(n1587), .ZN(n1871)
         );
  XNOR2_X1 U1518 ( .A(n1604), .B(n1872), .ZN(n816) );
  AOI221_X1 U1519 ( .B1(n1584), .B2(b[10]), .C1(n1585), .C2(b[9]), .A(n1873), 
        .ZN(n1872) );
  OAI22_X1 U1520 ( .A1(n1684), .A2(n1583), .B1(n1685), .B2(n1587), .ZN(n1873)
         );
  XNOR2_X1 U1521 ( .A(n1604), .B(n1874), .ZN(n815) );
  AOI221_X1 U1522 ( .B1(n1584), .B2(b[11]), .C1(n1585), .C2(b[10]), .A(n1875), 
        .ZN(n1874) );
  OAI22_X1 U1523 ( .A1(n1688), .A2(n1583), .B1(n1689), .B2(n1587), .ZN(n1875)
         );
  XNOR2_X1 U1524 ( .A(n1604), .B(n1876), .ZN(n814) );
  AOI221_X1 U1525 ( .B1(n1584), .B2(b[12]), .C1(n1585), .C2(b[11]), .A(n1877), 
        .ZN(n1876) );
  OAI22_X1 U1526 ( .A1(n1692), .A2(n1583), .B1(n1693), .B2(n1587), .ZN(n1877)
         );
  XNOR2_X1 U1527 ( .A(n1604), .B(n1878), .ZN(n813) );
  AOI221_X1 U1528 ( .B1(n1584), .B2(b[13]), .C1(n1585), .C2(b[12]), .A(n1879), 
        .ZN(n1878) );
  OAI22_X1 U1529 ( .A1(n1696), .A2(n1583), .B1(n1697), .B2(n1586), .ZN(n1879)
         );
  XNOR2_X1 U1530 ( .A(n1604), .B(n1880), .ZN(n812) );
  AOI221_X1 U1531 ( .B1(n1584), .B2(b[14]), .C1(n1585), .C2(b[13]), .A(n1881), 
        .ZN(n1880) );
  OAI22_X1 U1532 ( .A1(n1700), .A2(n1583), .B1(n1701), .B2(n1586), .ZN(n1881)
         );
  XNOR2_X1 U1533 ( .A(n1604), .B(n1882), .ZN(n811) );
  AOI221_X1 U1534 ( .B1(n1584), .B2(b[15]), .C1(n1585), .C2(b[14]), .A(n1883), 
        .ZN(n1882) );
  OAI22_X1 U1535 ( .A1(n1704), .A2(n1583), .B1(n1705), .B2(n1586), .ZN(n1883)
         );
  XNOR2_X1 U1536 ( .A(n1604), .B(n1884), .ZN(n810) );
  AOI221_X1 U1537 ( .B1(n1584), .B2(b[16]), .C1(n1585), .C2(b[15]), .A(n1885), 
        .ZN(n1884) );
  OAI22_X1 U1538 ( .A1(n1708), .A2(n1583), .B1(n1709), .B2(n1586), .ZN(n1885)
         );
  XNOR2_X1 U1539 ( .A(n1604), .B(n1886), .ZN(n809) );
  AOI221_X1 U1540 ( .B1(n1584), .B2(b[17]), .C1(n1585), .C2(b[16]), .A(n1887), 
        .ZN(n1886) );
  OAI22_X1 U1541 ( .A1(n1712), .A2(n1583), .B1(n1713), .B2(n1586), .ZN(n1887)
         );
  XNOR2_X1 U1542 ( .A(n1604), .B(n1888), .ZN(n808) );
  AOI221_X1 U1543 ( .B1(n1584), .B2(b[18]), .C1(n1585), .C2(b[17]), .A(n1889), 
        .ZN(n1888) );
  OAI22_X1 U1544 ( .A1(n1716), .A2(n1583), .B1(n1717), .B2(n1586), .ZN(n1889)
         );
  XNOR2_X1 U1545 ( .A(n1604), .B(n1890), .ZN(n807) );
  AOI221_X1 U1546 ( .B1(n1584), .B2(b[19]), .C1(n1585), .C2(b[18]), .A(n1891), 
        .ZN(n1890) );
  OAI22_X1 U1547 ( .A1(n1720), .A2(n1583), .B1(n1721), .B2(n1586), .ZN(n1891)
         );
  XNOR2_X1 U1548 ( .A(n1604), .B(n1892), .ZN(n806) );
  AOI221_X1 U1549 ( .B1(n1584), .B2(b[20]), .C1(n1585), .C2(b[19]), .A(n1893), 
        .ZN(n1892) );
  OAI22_X1 U1550 ( .A1(n1724), .A2(n1583), .B1(n1725), .B2(n1586), .ZN(n1893)
         );
  XNOR2_X1 U1551 ( .A(a[14]), .B(n1894), .ZN(n805) );
  AOI221_X1 U1552 ( .B1(n1584), .B2(b[21]), .C1(n1585), .C2(b[20]), .A(n1895), 
        .ZN(n1894) );
  OAI22_X1 U1553 ( .A1(n1728), .A2(n1583), .B1(n1729), .B2(n1586), .ZN(n1895)
         );
  XNOR2_X1 U1554 ( .A(a[14]), .B(n1896), .ZN(n804) );
  AOI221_X1 U1555 ( .B1(n1584), .B2(b[22]), .C1(n1553), .C2(n1376), .A(n1897), 
        .ZN(n1896) );
  OAI22_X1 U1556 ( .A1(n1640), .A2(n1587), .B1(n1643), .B2(n1550), .ZN(n1897)
         );
  XNOR2_X1 U1557 ( .A(a[14]), .B(n1898), .ZN(n803) );
  AOI221_X1 U1558 ( .B1(n1585), .B2(b[22]), .C1(n1553), .C2(n1375), .A(n1899), 
        .ZN(n1898) );
  OAI22_X1 U1559 ( .A1(n1617), .A2(n1541), .B1(n1643), .B2(n1586), .ZN(n1899)
         );
  XNOR2_X1 U1560 ( .A(a[14]), .B(n1900), .ZN(n802) );
  AOI221_X1 U1561 ( .B1(n1584), .B2(n1614), .C1(n1585), .C2(n1614), .A(n1901), 
        .ZN(n1900) );
  OAI22_X1 U1562 ( .A1(n1633), .A2(n1583), .B1(n1634), .B2(n1586), .ZN(n1901)
         );
  XNOR2_X1 U1563 ( .A(a[14]), .B(n1902), .ZN(n801) );
  OAI221_X1 U1564 ( .B1(n1617), .B2(n1587), .C1(n1619), .C2(n1583), .A(n1903), 
        .ZN(n1902) );
  OAI21_X1 U1565 ( .B1(n1584), .B2(n1585), .A(n1614), .ZN(n1903) );
  INV_X1 U1566 ( .A(n1907), .ZN(n1904) );
  NAND3_X1 U1567 ( .A1(n1907), .A2(n1906), .A3(n1905), .ZN(n1857) );
  XNOR2_X1 U1568 ( .A(a[12]), .B(a[13]), .ZN(n1905) );
  XNOR2_X1 U1569 ( .A(a[13]), .B(n1605), .ZN(n1906) );
  XOR2_X1 U1570 ( .A(a[12]), .B(n1607), .Z(n1907) );
  XNOR2_X1 U1571 ( .A(n1908), .B(n1603), .ZN(n800) );
  OAI22_X1 U1572 ( .A1(n1565), .A2(n1540), .B1(n1566), .B2(n1588), .ZN(n1908)
         );
  XNOR2_X1 U1573 ( .A(n1909), .B(n1603), .ZN(n799) );
  OAI222_X1 U1574 ( .A1(n1649), .A2(n1540), .B1(n1566), .B2(n1549), .C1(n1650), 
        .C2(n1588), .ZN(n1909) );
  XNOR2_X1 U1575 ( .A(n1602), .B(n1910), .ZN(n798) );
  AOI221_X1 U1576 ( .B1(n1589), .B2(b[2]), .C1(n1590), .C2(b[1]), .A(n1911), 
        .ZN(n1910) );
  OAI22_X1 U1577 ( .A1(n1653), .A2(n1588), .B1(n1566), .B2(n1591), .ZN(n1911)
         );
  XNOR2_X1 U1578 ( .A(n1602), .B(n1913), .ZN(n797) );
  AOI221_X1 U1579 ( .B1(n1589), .B2(b[3]), .C1(n1590), .C2(b[2]), .A(n1914), 
        .ZN(n1913) );
  OAI22_X1 U1580 ( .A1(n1657), .A2(n1588), .B1(n1649), .B2(n1592), .ZN(n1914)
         );
  XNOR2_X1 U1581 ( .A(n1602), .B(n1915), .ZN(n796) );
  AOI221_X1 U1582 ( .B1(n1589), .B2(b[4]), .C1(n1590), .C2(b[3]), .A(n1916), 
        .ZN(n1915) );
  OAI22_X1 U1583 ( .A1(n1660), .A2(n1588), .B1(n1661), .B2(n1592), .ZN(n1916)
         );
  XNOR2_X1 U1584 ( .A(n1602), .B(n1917), .ZN(n795) );
  AOI221_X1 U1585 ( .B1(n1589), .B2(b[5]), .C1(n1590), .C2(b[4]), .A(n1918), 
        .ZN(n1917) );
  OAI22_X1 U1586 ( .A1(n1664), .A2(n1588), .B1(n1665), .B2(n1592), .ZN(n1918)
         );
  XNOR2_X1 U1587 ( .A(n1602), .B(n1919), .ZN(n794) );
  AOI221_X1 U1588 ( .B1(n1589), .B2(b[6]), .C1(n1590), .C2(b[5]), .A(n1920), 
        .ZN(n1919) );
  OAI22_X1 U1589 ( .A1(n1668), .A2(n1588), .B1(n1669), .B2(n1592), .ZN(n1920)
         );
  XNOR2_X1 U1590 ( .A(n1602), .B(n1921), .ZN(n793) );
  AOI221_X1 U1591 ( .B1(n1589), .B2(b[7]), .C1(n1590), .C2(b[6]), .A(n1922), 
        .ZN(n1921) );
  OAI22_X1 U1592 ( .A1(n1672), .A2(n1588), .B1(n1673), .B2(n1592), .ZN(n1922)
         );
  XNOR2_X1 U1593 ( .A(n1602), .B(n1923), .ZN(n792) );
  AOI221_X1 U1594 ( .B1(n1589), .B2(b[8]), .C1(n1590), .C2(b[7]), .A(n1924), 
        .ZN(n1923) );
  OAI22_X1 U1595 ( .A1(n1676), .A2(n1588), .B1(n1677), .B2(n1592), .ZN(n1924)
         );
  XNOR2_X1 U1596 ( .A(n1602), .B(n1925), .ZN(n791) );
  AOI221_X1 U1597 ( .B1(n1589), .B2(b[9]), .C1(n1590), .C2(b[8]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1598 ( .A1(n1680), .A2(n1588), .B1(n1681), .B2(n1592), .ZN(n1926)
         );
  XNOR2_X1 U1599 ( .A(n1602), .B(n1927), .ZN(n790) );
  AOI221_X1 U1600 ( .B1(n1589), .B2(b[10]), .C1(n1590), .C2(b[9]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1601 ( .A1(n1684), .A2(n1588), .B1(n1685), .B2(n1592), .ZN(n1928)
         );
  XNOR2_X1 U1602 ( .A(n1602), .B(n1929), .ZN(n789) );
  AOI221_X1 U1603 ( .B1(n1589), .B2(b[11]), .C1(n1590), .C2(b[10]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1604 ( .A1(n1688), .A2(n1588), .B1(n1689), .B2(n1592), .ZN(n1930)
         );
  XNOR2_X1 U1605 ( .A(n1602), .B(n1931), .ZN(n788) );
  AOI221_X1 U1606 ( .B1(n1589), .B2(b[12]), .C1(n1590), .C2(b[11]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1607 ( .A1(n1692), .A2(n1588), .B1(n1693), .B2(n1592), .ZN(n1932)
         );
  XNOR2_X1 U1608 ( .A(n1602), .B(n1933), .ZN(n787) );
  AOI221_X1 U1609 ( .B1(n1589), .B2(b[13]), .C1(n1590), .C2(b[12]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1610 ( .A1(n1696), .A2(n1588), .B1(n1697), .B2(n1591), .ZN(n1934)
         );
  XNOR2_X1 U1611 ( .A(n1602), .B(n1935), .ZN(n786) );
  AOI221_X1 U1612 ( .B1(n1589), .B2(b[14]), .C1(n1590), .C2(b[13]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1613 ( .A1(n1700), .A2(n1588), .B1(n1701), .B2(n1591), .ZN(n1936)
         );
  XNOR2_X1 U1614 ( .A(n1602), .B(n1937), .ZN(n785) );
  AOI221_X1 U1615 ( .B1(n1589), .B2(b[15]), .C1(n1590), .C2(b[14]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1616 ( .A1(n1704), .A2(n1588), .B1(n1705), .B2(n1591), .ZN(n1938)
         );
  XNOR2_X1 U1617 ( .A(n1602), .B(n1939), .ZN(n784) );
  AOI221_X1 U1618 ( .B1(n1589), .B2(b[16]), .C1(n1590), .C2(b[15]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1619 ( .A1(n1708), .A2(n1588), .B1(n1709), .B2(n1591), .ZN(n1940)
         );
  XNOR2_X1 U1620 ( .A(n1602), .B(n1941), .ZN(n783) );
  AOI221_X1 U1621 ( .B1(n1589), .B2(b[17]), .C1(n1590), .C2(b[16]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1622 ( .A1(n1712), .A2(n1588), .B1(n1713), .B2(n1591), .ZN(n1942)
         );
  XNOR2_X1 U1623 ( .A(n1602), .B(n1943), .ZN(n782) );
  AOI221_X1 U1624 ( .B1(n1589), .B2(b[18]), .C1(n1590), .C2(b[17]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1625 ( .A1(n1716), .A2(n1588), .B1(n1717), .B2(n1591), .ZN(n1944)
         );
  XNOR2_X1 U1626 ( .A(n1602), .B(n1945), .ZN(n781) );
  AOI221_X1 U1627 ( .B1(n1589), .B2(b[19]), .C1(n1590), .C2(b[18]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1628 ( .A1(n1720), .A2(n1588), .B1(n1721), .B2(n1591), .ZN(n1946)
         );
  XNOR2_X1 U1629 ( .A(n1602), .B(n1947), .ZN(n780) );
  AOI221_X1 U1630 ( .B1(n1589), .B2(b[20]), .C1(n1590), .C2(b[19]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1631 ( .A1(n1724), .A2(n1588), .B1(n1725), .B2(n1591), .ZN(n1948)
         );
  XNOR2_X1 U1632 ( .A(a[17]), .B(n1949), .ZN(n779) );
  AOI221_X1 U1633 ( .B1(n1589), .B2(b[21]), .C1(n1590), .C2(b[20]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1634 ( .A1(n1728), .A2(n1588), .B1(n1729), .B2(n1591), .ZN(n1950)
         );
  XNOR2_X1 U1635 ( .A(a[17]), .B(n1951), .ZN(n778) );
  AOI221_X1 U1636 ( .B1(n1589), .B2(b[22]), .C1(n1552), .C2(n1376), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1637 ( .A1(n1640), .A2(n1592), .B1(n1643), .B2(n1549), .ZN(n1952)
         );
  XNOR2_X1 U1638 ( .A(a[17]), .B(n1953), .ZN(n777) );
  AOI221_X1 U1639 ( .B1(n1590), .B2(b[22]), .C1(n1552), .C2(n1375), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1640 ( .A1(n1617), .A2(n1540), .B1(n1643), .B2(n1591), .ZN(n1954)
         );
  XNOR2_X1 U1641 ( .A(a[17]), .B(n1955), .ZN(n776) );
  AOI221_X1 U1642 ( .B1(n1589), .B2(n1613), .C1(n1590), .C2(n1614), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1643 ( .A1(n1633), .A2(n1588), .B1(n1634), .B2(n1591), .ZN(n1956)
         );
  XNOR2_X1 U1644 ( .A(a[17]), .B(n1957), .ZN(n775) );
  OAI221_X1 U1645 ( .B1(n1618), .B2(n1592), .C1(n1617), .C2(n1588), .A(n1958), 
        .ZN(n1957) );
  OAI21_X1 U1646 ( .B1(n1589), .B2(n1590), .A(n1614), .ZN(n1958) );
  INV_X1 U1647 ( .A(n1962), .ZN(n1959) );
  NAND3_X1 U1648 ( .A1(n1962), .A2(n1961), .A3(n1960), .ZN(n1912) );
  XNOR2_X1 U1649 ( .A(a[15]), .B(a[16]), .ZN(n1960) );
  XNOR2_X1 U1650 ( .A(a[16]), .B(n1603), .ZN(n1961) );
  XOR2_X1 U1651 ( .A(a[15]), .B(n1605), .Z(n1962) );
  XOR2_X1 U1652 ( .A(n1963), .B(n1600), .Z(n774) );
  OAI22_X1 U1653 ( .A1(n1565), .A2(n1539), .B1(n1566), .B2(n1593), .ZN(n1963)
         );
  XOR2_X1 U1654 ( .A(n1964), .B(n1600), .Z(n773) );
  OAI222_X1 U1655 ( .A1(n1649), .A2(n1539), .B1(n1566), .B2(n1548), .C1(n1650), 
        .C2(n1593), .ZN(n1964) );
  XNOR2_X1 U1656 ( .A(n1600), .B(n1965), .ZN(n772) );
  AOI221_X1 U1657 ( .B1(n1594), .B2(b[2]), .C1(n1595), .C2(b[1]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1658 ( .A1(n1653), .A2(n1593), .B1(n1566), .B2(n1596), .ZN(n1966)
         );
  XNOR2_X1 U1659 ( .A(n1600), .B(n1968), .ZN(n771) );
  AOI221_X1 U1660 ( .B1(n1594), .B2(b[3]), .C1(n1595), .C2(b[2]), .A(n1969), 
        .ZN(n1968) );
  OAI22_X1 U1661 ( .A1(n1657), .A2(n1593), .B1(n1649), .B2(n1597), .ZN(n1969)
         );
  XNOR2_X1 U1662 ( .A(n1600), .B(n1970), .ZN(n770) );
  AOI221_X1 U1663 ( .B1(n1594), .B2(b[4]), .C1(n1595), .C2(b[3]), .A(n1971), 
        .ZN(n1970) );
  OAI22_X1 U1664 ( .A1(n1660), .A2(n1593), .B1(n1661), .B2(n1597), .ZN(n1971)
         );
  XNOR2_X1 U1665 ( .A(n1600), .B(n1972), .ZN(n769) );
  AOI221_X1 U1666 ( .B1(n1594), .B2(b[5]), .C1(n1595), .C2(b[4]), .A(n1973), 
        .ZN(n1972) );
  OAI22_X1 U1667 ( .A1(n1664), .A2(n1593), .B1(n1665), .B2(n1597), .ZN(n1973)
         );
  XNOR2_X1 U1668 ( .A(n1600), .B(n1974), .ZN(n768) );
  AOI221_X1 U1669 ( .B1(n1594), .B2(b[6]), .C1(n1595), .C2(b[5]), .A(n1975), 
        .ZN(n1974) );
  OAI22_X1 U1670 ( .A1(n1668), .A2(n1593), .B1(n1669), .B2(n1597), .ZN(n1975)
         );
  XNOR2_X1 U1671 ( .A(n1600), .B(n1976), .ZN(n767) );
  AOI221_X1 U1672 ( .B1(n1594), .B2(b[7]), .C1(n1595), .C2(b[6]), .A(n1977), 
        .ZN(n1976) );
  OAI22_X1 U1673 ( .A1(n1672), .A2(n1593), .B1(n1673), .B2(n1597), .ZN(n1977)
         );
  XNOR2_X1 U1674 ( .A(n1600), .B(n1978), .ZN(n766) );
  AOI221_X1 U1675 ( .B1(n1594), .B2(b[8]), .C1(n1595), .C2(b[7]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1676 ( .A1(n1676), .A2(n1593), .B1(n1677), .B2(n1597), .ZN(n1979)
         );
  XNOR2_X1 U1677 ( .A(n1600), .B(n1980), .ZN(n765) );
  AOI221_X1 U1678 ( .B1(n1594), .B2(b[9]), .C1(n1595), .C2(b[8]), .A(n1981), 
        .ZN(n1980) );
  OAI22_X1 U1679 ( .A1(n1680), .A2(n1593), .B1(n1681), .B2(n1597), .ZN(n1981)
         );
  XNOR2_X1 U1680 ( .A(n1600), .B(n1982), .ZN(n764) );
  AOI221_X1 U1681 ( .B1(n1594), .B2(b[10]), .C1(n1595), .C2(b[9]), .A(n1983), 
        .ZN(n1982) );
  OAI22_X1 U1682 ( .A1(n1684), .A2(n1593), .B1(n1685), .B2(n1597), .ZN(n1983)
         );
  XNOR2_X1 U1683 ( .A(n1600), .B(n1984), .ZN(n763) );
  AOI221_X1 U1684 ( .B1(n1594), .B2(b[11]), .C1(n1595), .C2(b[10]), .A(n1985), 
        .ZN(n1984) );
  OAI22_X1 U1685 ( .A1(n1688), .A2(n1593), .B1(n1689), .B2(n1597), .ZN(n1985)
         );
  XNOR2_X1 U1686 ( .A(n1601), .B(n1986), .ZN(n762) );
  AOI221_X1 U1687 ( .B1(n1594), .B2(b[12]), .C1(n1595), .C2(b[11]), .A(n1987), 
        .ZN(n1986) );
  OAI22_X1 U1688 ( .A1(n1692), .A2(n1593), .B1(n1693), .B2(n1597), .ZN(n1987)
         );
  XNOR2_X1 U1689 ( .A(n1601), .B(n1988), .ZN(n761) );
  AOI221_X1 U1690 ( .B1(n1594), .B2(b[13]), .C1(n1595), .C2(b[12]), .A(n1989), 
        .ZN(n1988) );
  OAI22_X1 U1691 ( .A1(n1696), .A2(n1593), .B1(n1697), .B2(n1596), .ZN(n1989)
         );
  XNOR2_X1 U1692 ( .A(n1601), .B(n1990), .ZN(n760) );
  AOI221_X1 U1693 ( .B1(n1594), .B2(b[14]), .C1(n1595), .C2(b[13]), .A(n1991), 
        .ZN(n1990) );
  OAI22_X1 U1694 ( .A1(n1700), .A2(n1593), .B1(n1701), .B2(n1596), .ZN(n1991)
         );
  XNOR2_X1 U1695 ( .A(n1601), .B(n1992), .ZN(n759) );
  AOI221_X1 U1696 ( .B1(n1594), .B2(b[15]), .C1(n1595), .C2(b[14]), .A(n1993), 
        .ZN(n1992) );
  OAI22_X1 U1697 ( .A1(n1704), .A2(n1593), .B1(n1705), .B2(n1596), .ZN(n1993)
         );
  XNOR2_X1 U1698 ( .A(n1601), .B(n1994), .ZN(n758) );
  AOI221_X1 U1699 ( .B1(n1594), .B2(b[16]), .C1(n1595), .C2(b[15]), .A(n1995), 
        .ZN(n1994) );
  OAI22_X1 U1700 ( .A1(n1708), .A2(n1593), .B1(n1709), .B2(n1596), .ZN(n1995)
         );
  XNOR2_X1 U1701 ( .A(n1601), .B(n1996), .ZN(n757) );
  AOI221_X1 U1702 ( .B1(n1594), .B2(b[17]), .C1(n1595), .C2(b[16]), .A(n1997), 
        .ZN(n1996) );
  OAI22_X1 U1703 ( .A1(n1712), .A2(n1593), .B1(n1713), .B2(n1596), .ZN(n1997)
         );
  XNOR2_X1 U1704 ( .A(n1601), .B(n1998), .ZN(n756) );
  AOI221_X1 U1705 ( .B1(n1594), .B2(b[18]), .C1(n1595), .C2(b[17]), .A(n1999), 
        .ZN(n1998) );
  OAI22_X1 U1706 ( .A1(n1716), .A2(n1593), .B1(n1717), .B2(n1596), .ZN(n1999)
         );
  XNOR2_X1 U1707 ( .A(n1601), .B(n2000), .ZN(n755) );
  AOI221_X1 U1708 ( .B1(n1594), .B2(b[19]), .C1(n1595), .C2(b[18]), .A(n2001), 
        .ZN(n2000) );
  OAI22_X1 U1709 ( .A1(n1720), .A2(n1593), .B1(n1721), .B2(n1596), .ZN(n2001)
         );
  XNOR2_X1 U1710 ( .A(n1601), .B(n2002), .ZN(n754) );
  AOI221_X1 U1711 ( .B1(n1594), .B2(b[20]), .C1(n1595), .C2(b[19]), .A(n2003), 
        .ZN(n2002) );
  OAI22_X1 U1712 ( .A1(n1724), .A2(n1593), .B1(n1725), .B2(n1596), .ZN(n2003)
         );
  XNOR2_X1 U1713 ( .A(n1601), .B(n2004), .ZN(n753) );
  AOI221_X1 U1714 ( .B1(n1594), .B2(b[21]), .C1(n1595), .C2(b[20]), .A(n2005), 
        .ZN(n2004) );
  OAI22_X1 U1715 ( .A1(n1728), .A2(n1593), .B1(n1729), .B2(n1596), .ZN(n2005)
         );
  XNOR2_X1 U1716 ( .A(n1601), .B(n2006), .ZN(n752) );
  AOI221_X1 U1717 ( .B1(n1594), .B2(b[22]), .C1(n1545), .C2(n1376), .A(n2007), 
        .ZN(n2006) );
  OAI22_X1 U1718 ( .A1(n1640), .A2(n1597), .B1(n1643), .B2(n1548), .ZN(n2007)
         );
  XNOR2_X1 U1719 ( .A(n1601), .B(n2008), .ZN(n751) );
  AOI221_X1 U1720 ( .B1(n1595), .B2(b[22]), .C1(n1545), .C2(n1375), .A(n2009), 
        .ZN(n2008) );
  OAI22_X1 U1721 ( .A1(n1617), .A2(n1539), .B1(n1643), .B2(n1596), .ZN(n2009)
         );
  XNOR2_X1 U1722 ( .A(n1601), .B(n2010), .ZN(n750) );
  AOI221_X1 U1723 ( .B1(n1594), .B2(n1612), .C1(n1595), .C2(n1614), .A(n2011), 
        .ZN(n2010) );
  OAI22_X1 U1724 ( .A1(n1633), .A2(n1593), .B1(n1634), .B2(n1596), .ZN(n2011)
         );
  INV_X1 U1725 ( .A(b[22]), .ZN(n1634) );
  INV_X1 U1726 ( .A(n1374), .ZN(n1633) );
  XNOR2_X1 U1727 ( .A(n1600), .B(n2012), .ZN(n749) );
  OAI221_X1 U1728 ( .B1(n1617), .B2(n1597), .C1(n1619), .C2(n1593), .A(n2013), 
        .ZN(n2012) );
  OAI21_X1 U1729 ( .B1(n1594), .B2(n1595), .A(n1614), .ZN(n2013) );
  INV_X1 U1730 ( .A(n2017), .ZN(n2014) );
  NAND3_X1 U1731 ( .A1(n2017), .A2(n2016), .A3(n2015), .ZN(n1967) );
  XNOR2_X1 U1732 ( .A(a[18]), .B(a[19]), .ZN(n2015) );
  XOR2_X1 U1733 ( .A(a[19]), .B(n1600), .Z(n2016) );
  XOR2_X1 U1734 ( .A(a[18]), .B(n1603), .Z(n2017) );
  XNOR2_X1 U1735 ( .A(n2018), .B(n1599), .ZN(n748) );
  OAI22_X1 U1736 ( .A1(n1538), .A2(n1567), .B1(n1558), .B2(n1567), .ZN(n2018)
         );
  XNOR2_X1 U1737 ( .A(n2019), .B(n1599), .ZN(n747) );
  OAI222_X1 U1738 ( .A1(n1538), .A2(n1649), .B1(n1547), .B2(n1566), .C1(n1558), 
        .C2(n1650), .ZN(n2019) );
  XNOR2_X1 U1739 ( .A(n1598), .B(n2020), .ZN(n746) );
  AOI221_X1 U1740 ( .B1(b[2]), .B2(n1559), .C1(b[1]), .C2(n1560), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1741 ( .A1(n1558), .A2(n1653), .B1(n1557), .B2(n1567), .ZN(n2021)
         );
  INV_X1 U1742 ( .A(b[0]), .ZN(n1647) );
  INV_X1 U1743 ( .A(n1396), .ZN(n1653) );
  XNOR2_X1 U1744 ( .A(n1598), .B(n2022), .ZN(n745) );
  AOI221_X1 U1745 ( .B1(b[3]), .B2(n1559), .C1(b[2]), .C2(n1560), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1746 ( .A1(n1558), .A2(n1657), .B1(n1557), .B2(n1649), .ZN(n2023)
         );
  XNOR2_X1 U1747 ( .A(n1598), .B(n2024), .ZN(n744) );
  AOI221_X1 U1748 ( .B1(b[4]), .B2(n1559), .C1(b[3]), .C2(n1560), .A(n2025), 
        .ZN(n2024) );
  OAI22_X1 U1749 ( .A1(n1558), .A2(n1660), .B1(n1557), .B2(n1661), .ZN(n2025)
         );
  XNOR2_X1 U1750 ( .A(n1598), .B(n2026), .ZN(n743) );
  AOI221_X1 U1751 ( .B1(b[5]), .B2(n1559), .C1(b[4]), .C2(n1560), .A(n2027), 
        .ZN(n2026) );
  OAI22_X1 U1752 ( .A1(n1558), .A2(n1664), .B1(n1557), .B2(n1665), .ZN(n2027)
         );
  XNOR2_X1 U1753 ( .A(n1598), .B(n2028), .ZN(n742) );
  AOI221_X1 U1754 ( .B1(b[6]), .B2(n1559), .C1(b[5]), .C2(n1560), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1755 ( .A1(n1558), .A2(n1668), .B1(n1557), .B2(n1669), .ZN(n2029)
         );
  XNOR2_X1 U1756 ( .A(n1598), .B(n2030), .ZN(n741) );
  AOI221_X1 U1757 ( .B1(b[7]), .B2(n1559), .C1(b[6]), .C2(n1560), .A(n2031), 
        .ZN(n2030) );
  OAI22_X1 U1758 ( .A1(n1558), .A2(n1672), .B1(n1557), .B2(n1673), .ZN(n2031)
         );
  XNOR2_X1 U1759 ( .A(n1598), .B(n2032), .ZN(n740) );
  AOI221_X1 U1760 ( .B1(b[9]), .B2(n1559), .C1(b[8]), .C2(n1560), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1761 ( .A1(n1558), .A2(n1680), .B1(n1557), .B2(n1681), .ZN(n2033)
         );
  XNOR2_X1 U1762 ( .A(n1598), .B(n2034), .ZN(n739) );
  AOI221_X1 U1763 ( .B1(b[10]), .B2(n1559), .C1(b[9]), .C2(n1560), .A(n2035), 
        .ZN(n2034) );
  OAI22_X1 U1764 ( .A1(n1558), .A2(n1684), .B1(n1557), .B2(n1685), .ZN(n2035)
         );
  XNOR2_X1 U1765 ( .A(n1598), .B(n2036), .ZN(n738) );
  AOI221_X1 U1766 ( .B1(b[12]), .B2(n1559), .C1(b[11]), .C2(n1560), .A(n2037), 
        .ZN(n2036) );
  OAI22_X1 U1767 ( .A1(n1558), .A2(n1692), .B1(n1557), .B2(n1693), .ZN(n2037)
         );
  XNOR2_X1 U1768 ( .A(n1598), .B(n2038), .ZN(n737) );
  AOI221_X1 U1769 ( .B1(b[13]), .B2(n1559), .C1(b[12]), .C2(n1560), .A(n2039), 
        .ZN(n2038) );
  OAI22_X1 U1770 ( .A1(n1558), .A2(n1696), .B1(n1557), .B2(n1697), .ZN(n2039)
         );
  XNOR2_X1 U1771 ( .A(n1598), .B(n2040), .ZN(n736) );
  AOI221_X1 U1772 ( .B1(b[14]), .B2(n1559), .C1(b[13]), .C2(n1560), .A(n2041), 
        .ZN(n2040) );
  OAI22_X1 U1773 ( .A1(n1558), .A2(n1700), .B1(n1556), .B2(n1701), .ZN(n2041)
         );
  XNOR2_X1 U1774 ( .A(n1598), .B(n2042), .ZN(n735) );
  AOI221_X1 U1775 ( .B1(b[15]), .B2(n1559), .C1(b[14]), .C2(n1560), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1776 ( .A1(n1558), .A2(n1704), .B1(n1556), .B2(n1705), .ZN(n2043)
         );
  XNOR2_X1 U1777 ( .A(n1598), .B(n2044), .ZN(n734) );
  AOI221_X1 U1778 ( .B1(b[16]), .B2(n1559), .C1(b[15]), .C2(n1560), .A(n2045), 
        .ZN(n2044) );
  OAI22_X1 U1779 ( .A1(n1558), .A2(n1708), .B1(n1556), .B2(n1709), .ZN(n2045)
         );
  XNOR2_X1 U1780 ( .A(n1598), .B(n2046), .ZN(n733) );
  AOI221_X1 U1781 ( .B1(b[18]), .B2(n1559), .C1(b[17]), .C2(n1560), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1782 ( .A1(n1558), .A2(n1716), .B1(n1556), .B2(n1717), .ZN(n2047)
         );
  XNOR2_X1 U1783 ( .A(n1598), .B(n2048), .ZN(n732) );
  AOI221_X1 U1784 ( .B1(b[19]), .B2(n1559), .C1(b[18]), .C2(n1560), .A(n2049), 
        .ZN(n2048) );
  OAI22_X1 U1785 ( .A1(n1558), .A2(n1720), .B1(n1556), .B2(n1721), .ZN(n2049)
         );
  XNOR2_X1 U1786 ( .A(n1598), .B(n2050), .ZN(n731) );
  AOI221_X1 U1787 ( .B1(b[20]), .B2(n1559), .C1(b[19]), .C2(n1560), .A(n2051), 
        .ZN(n2050) );
  OAI22_X1 U1788 ( .A1(n1558), .A2(n1724), .B1(n1556), .B2(n1725), .ZN(n2051)
         );
  XNOR2_X1 U1789 ( .A(a[23]), .B(n2052), .ZN(n730) );
  AOI221_X1 U1790 ( .B1(b[21]), .B2(n1559), .C1(b[20]), .C2(n1560), .A(n2053), 
        .ZN(n2052) );
  OAI22_X1 U1791 ( .A1(n1558), .A2(n1728), .B1(n1556), .B2(n1729), .ZN(n2053)
         );
  XNOR2_X1 U1792 ( .A(a[23]), .B(n2054), .ZN(n729) );
  AOI221_X1 U1793 ( .B1(b[22]), .B2(n1559), .C1(n1376), .C2(n1544), .A(n2055), 
        .ZN(n2054) );
  OAI22_X1 U1794 ( .A1(n1556), .A2(n1640), .B1(n1547), .B2(n1643), .ZN(n2055)
         );
  INV_X1 U1795 ( .A(b[20]), .ZN(n1640) );
  XNOR2_X1 U1796 ( .A(n519), .B(n2056), .ZN(n506) );
  INV_X1 U1797 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1798 ( .A1(n2056), .A2(n519), .ZN(n493) );
  XOR2_X1 U1799 ( .A(n2057), .B(n1742), .Z(n2056) );
  OAI221_X1 U1800 ( .B1(n1618), .B2(n1639), .C1(n1619), .C2(n1564), .A(n2058), 
        .ZN(n2057) );
  OAI21_X1 U1801 ( .B1(n1561), .B2(n1563), .A(n1614), .ZN(n2058) );
  INV_X1 U1802 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1803 ( .A(n1598), .B(n2059), .Z(n454) );
  AOI221_X1 U1804 ( .B1(b[8]), .B2(n1559), .C1(b[7]), .C2(n1560), .A(n2060), 
        .ZN(n2059) );
  OAI22_X1 U1805 ( .A1(n1558), .A2(n1676), .B1(n1556), .B2(n1677), .ZN(n2060)
         );
  INV_X1 U1806 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1807 ( .A(n1598), .B(n2061), .Z(n421) );
  AOI221_X1 U1808 ( .B1(b[11]), .B2(n1559), .C1(b[10]), .C2(n1560), .A(n2062), 
        .ZN(n2061) );
  OAI22_X1 U1809 ( .A1(n1558), .A2(n1688), .B1(n1556), .B2(n1689), .ZN(n2062)
         );
  INV_X1 U1810 ( .A(n387), .ZN(n395) );
  INV_X1 U1811 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1812 ( .A(n1598), .B(n2063), .Z(n374) );
  AOI221_X1 U1813 ( .B1(b[17]), .B2(n1559), .C1(b[16]), .C2(n1560), .A(n2064), 
        .ZN(n2063) );
  OAI22_X1 U1814 ( .A1(n1558), .A2(n1712), .B1(n1556), .B2(n1713), .ZN(n2064)
         );
  INV_X1 U1815 ( .A(n356), .ZN(n360) );
  INV_X1 U1816 ( .A(n1627), .ZN(n351) );
  XOR2_X1 U1817 ( .A(n1599), .B(n2065), .Z(n1627) );
  AOI221_X1 U1818 ( .B1(b[22]), .B2(n1560), .C1(n1375), .C2(n1544), .A(n2066), 
        .ZN(n2065) );
  OAI22_X1 U1819 ( .A1(n1538), .A2(n1618), .B1(n1556), .B2(n1643), .ZN(n2066)
         );
  INV_X1 U1820 ( .A(b[21]), .ZN(n1643) );
  NAND3_X1 U1821 ( .A1(n2067), .A2(n2068), .A3(n2069), .ZN(n1629) );
  XNOR2_X1 U1822 ( .A(a[22]), .B(n1599), .ZN(n2068) );
  XNOR2_X1 U1823 ( .A(a[21]), .B(a[22]), .ZN(n2069) );
  INV_X1 U1824 ( .A(n2067), .ZN(n2070) );
  XNOR2_X1 U1825 ( .A(a[21]), .B(n1600), .ZN(n2067) );
  OAI222_X1 U1826 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n2073), .C1(n2073), 
        .C2(n2072), .ZN(n326) );
  INV_X1 U1827 ( .A(n550), .ZN(n2073) );
  XNOR2_X1 U1828 ( .A(n1742), .B(n2074), .ZN(n2072) );
  AOI221_X1 U1829 ( .B1(n1561), .B2(b[21]), .C1(b[20]), .C2(n1562), .A(n2075), 
        .ZN(n2074) );
  OAI22_X1 U1830 ( .A1(n1564), .A2(n1728), .B1(n1639), .B2(n1729), .ZN(n2075)
         );
  INV_X1 U1831 ( .A(b[19]), .ZN(n1729) );
  INV_X1 U1832 ( .A(n1377), .ZN(n1728) );
  AOI222_X1 U1833 ( .A1(n2076), .A2(n2077), .B1(n2076), .B2(n564), .C1(n564), 
        .C2(n2077), .ZN(n2071) );
  XNOR2_X1 U1834 ( .A(a[2]), .B(n2078), .ZN(n2077) );
  AOI221_X1 U1835 ( .B1(b[20]), .B2(n1561), .C1(b[19]), .C2(n1562), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1836 ( .A1(n1564), .A2(n1724), .B1(n1639), .B2(n1725), .ZN(n2079)
         );
  INV_X1 U1837 ( .A(b[18]), .ZN(n1725) );
  INV_X1 U1838 ( .A(n1378), .ZN(n1724) );
  INV_X1 U1839 ( .A(n2080), .ZN(n2076) );
  AOI222_X1 U1840 ( .A1(n2081), .A2(n2082), .B1(n2081), .B2(n576), .C1(n576), 
        .C2(n2082), .ZN(n2080) );
  XNOR2_X1 U1841 ( .A(a[2]), .B(n2083), .ZN(n2082) );
  AOI221_X1 U1842 ( .B1(b[19]), .B2(n1561), .C1(b[18]), .C2(n1562), .A(n2084), 
        .ZN(n2083) );
  OAI22_X1 U1843 ( .A1(n1564), .A2(n1720), .B1(n1639), .B2(n1721), .ZN(n2084)
         );
  INV_X1 U1844 ( .A(b[17]), .ZN(n1721) );
  INV_X1 U1845 ( .A(n1379), .ZN(n1720) );
  OAI222_X1 U1846 ( .A1(n2085), .A2(n2086), .B1(n2085), .B2(n2087), .C1(n2087), 
        .C2(n2086), .ZN(n2081) );
  INV_X1 U1847 ( .A(n588), .ZN(n2087) );
  XNOR2_X1 U1848 ( .A(n1742), .B(n2088), .ZN(n2086) );
  AOI221_X1 U1849 ( .B1(b[18]), .B2(n1561), .C1(b[17]), .C2(n1562), .A(n2089), 
        .ZN(n2088) );
  OAI22_X1 U1850 ( .A1(n1564), .A2(n1716), .B1(n1639), .B2(n1717), .ZN(n2089)
         );
  INV_X1 U1851 ( .A(b[16]), .ZN(n1717) );
  INV_X1 U1852 ( .A(n1380), .ZN(n1716) );
  AOI222_X1 U1853 ( .A1(n2090), .A2(n2091), .B1(n2090), .B2(n600), .C1(n600), 
        .C2(n2091), .ZN(n2085) );
  XNOR2_X1 U1854 ( .A(a[2]), .B(n2092), .ZN(n2091) );
  AOI221_X1 U1855 ( .B1(b[17]), .B2(n1561), .C1(b[16]), .C2(n1562), .A(n2093), 
        .ZN(n2092) );
  OAI22_X1 U1856 ( .A1(n1564), .A2(n1712), .B1(n1639), .B2(n1713), .ZN(n2093)
         );
  INV_X1 U1857 ( .A(b[15]), .ZN(n1713) );
  INV_X1 U1858 ( .A(n1381), .ZN(n1712) );
  OAI222_X1 U1859 ( .A1(n2094), .A2(n2095), .B1(n2094), .B2(n2096), .C1(n2096), 
        .C2(n2095), .ZN(n2090) );
  INV_X1 U1860 ( .A(n610), .ZN(n2096) );
  XNOR2_X1 U1861 ( .A(n1742), .B(n2097), .ZN(n2095) );
  AOI221_X1 U1862 ( .B1(b[16]), .B2(n1561), .C1(b[15]), .C2(n1562), .A(n2098), 
        .ZN(n2097) );
  OAI22_X1 U1863 ( .A1(n1564), .A2(n1708), .B1(n1639), .B2(n1709), .ZN(n2098)
         );
  INV_X1 U1864 ( .A(b[14]), .ZN(n1709) );
  INV_X1 U1865 ( .A(n1382), .ZN(n1708) );
  AOI222_X1 U1866 ( .A1(n2099), .A2(n2100), .B1(n2099), .B2(n620), .C1(n620), 
        .C2(n2100), .ZN(n2094) );
  XNOR2_X1 U1867 ( .A(a[2]), .B(n2101), .ZN(n2100) );
  AOI221_X1 U1868 ( .B1(b[15]), .B2(n1561), .C1(b[14]), .C2(n1562), .A(n2102), 
        .ZN(n2101) );
  OAI22_X1 U1869 ( .A1(n1564), .A2(n1704), .B1(n1639), .B2(n1705), .ZN(n2102)
         );
  INV_X1 U1870 ( .A(b[13]), .ZN(n1705) );
  INV_X1 U1871 ( .A(n1383), .ZN(n1704) );
  OAI222_X1 U1872 ( .A1(n2103), .A2(n2104), .B1(n2103), .B2(n2105), .C1(n2105), 
        .C2(n2104), .ZN(n2099) );
  INV_X1 U1873 ( .A(n630), .ZN(n2105) );
  XNOR2_X1 U1874 ( .A(n1742), .B(n2106), .ZN(n2104) );
  AOI221_X1 U1875 ( .B1(b[14]), .B2(n1561), .C1(b[13]), .C2(n1562), .A(n2107), 
        .ZN(n2106) );
  OAI22_X1 U1876 ( .A1(n1564), .A2(n1700), .B1(n1639), .B2(n1701), .ZN(n2107)
         );
  INV_X1 U1877 ( .A(b[12]), .ZN(n1701) );
  INV_X1 U1878 ( .A(n1384), .ZN(n1700) );
  AOI222_X1 U1879 ( .A1(n2108), .A2(n2109), .B1(n2108), .B2(n638), .C1(n638), 
        .C2(n2109), .ZN(n2103) );
  XNOR2_X1 U1880 ( .A(a[2]), .B(n2110), .ZN(n2109) );
  AOI221_X1 U1881 ( .B1(b[13]), .B2(n1561), .C1(b[12]), .C2(n1562), .A(n2111), 
        .ZN(n2110) );
  OAI22_X1 U1882 ( .A1(n1564), .A2(n1696), .B1(n1639), .B2(n1697), .ZN(n2111)
         );
  INV_X1 U1883 ( .A(b[11]), .ZN(n1697) );
  INV_X1 U1884 ( .A(n1385), .ZN(n1696) );
  OAI222_X1 U1885 ( .A1(n2112), .A2(n2113), .B1(n2112), .B2(n2114), .C1(n2114), 
        .C2(n2113), .ZN(n2108) );
  INV_X1 U1886 ( .A(n646), .ZN(n2114) );
  XNOR2_X1 U1887 ( .A(n1742), .B(n2115), .ZN(n2113) );
  AOI221_X1 U1888 ( .B1(b[12]), .B2(n1561), .C1(b[11]), .C2(n1562), .A(n2116), 
        .ZN(n2115) );
  OAI22_X1 U1889 ( .A1(n1564), .A2(n1692), .B1(n1639), .B2(n1693), .ZN(n2116)
         );
  INV_X1 U1890 ( .A(b[10]), .ZN(n1693) );
  INV_X1 U1891 ( .A(n1386), .ZN(n1692) );
  AOI222_X1 U1892 ( .A1(n2117), .A2(n2118), .B1(n2117), .B2(n654), .C1(n654), 
        .C2(n2118), .ZN(n2112) );
  XNOR2_X1 U1893 ( .A(a[2]), .B(n2119), .ZN(n2118) );
  AOI221_X1 U1894 ( .B1(b[11]), .B2(n1561), .C1(b[10]), .C2(n1562), .A(n2120), 
        .ZN(n2119) );
  OAI22_X1 U1895 ( .A1(n1564), .A2(n1688), .B1(n1639), .B2(n1689), .ZN(n2120)
         );
  INV_X1 U1896 ( .A(b[9]), .ZN(n1689) );
  INV_X1 U1897 ( .A(n1387), .ZN(n1688) );
  OAI222_X1 U1898 ( .A1(n2121), .A2(n2122), .B1(n2121), .B2(n2123), .C1(n2123), 
        .C2(n2122), .ZN(n2117) );
  INV_X1 U1899 ( .A(n660), .ZN(n2123) );
  XNOR2_X1 U1900 ( .A(n1742), .B(n2124), .ZN(n2122) );
  AOI221_X1 U1901 ( .B1(b[10]), .B2(n1561), .C1(b[9]), .C2(n1563), .A(n2125), 
        .ZN(n2124) );
  OAI22_X1 U1902 ( .A1(n1564), .A2(n1684), .B1(n1639), .B2(n1685), .ZN(n2125)
         );
  INV_X1 U1903 ( .A(b[8]), .ZN(n1685) );
  INV_X1 U1904 ( .A(n1388), .ZN(n1684) );
  AOI222_X1 U1905 ( .A1(n2126), .A2(n2127), .B1(n2126), .B2(n666), .C1(n666), 
        .C2(n2127), .ZN(n2121) );
  XNOR2_X1 U1906 ( .A(a[2]), .B(n2128), .ZN(n2127) );
  AOI221_X1 U1907 ( .B1(b[9]), .B2(n1561), .C1(b[8]), .C2(n1563), .A(n2129), 
        .ZN(n2128) );
  OAI22_X1 U1908 ( .A1(n1564), .A2(n1680), .B1(n1639), .B2(n1681), .ZN(n2129)
         );
  INV_X1 U1909 ( .A(b[7]), .ZN(n1681) );
  INV_X1 U1910 ( .A(n1389), .ZN(n1680) );
  OAI222_X1 U1911 ( .A1(n2130), .A2(n2131), .B1(n2130), .B2(n2132), .C1(n2132), 
        .C2(n2131), .ZN(n2126) );
  INV_X1 U1912 ( .A(n672), .ZN(n2132) );
  XNOR2_X1 U1913 ( .A(n1742), .B(n2133), .ZN(n2131) );
  AOI221_X1 U1914 ( .B1(b[8]), .B2(n1561), .C1(b[7]), .C2(n1562), .A(n2134), 
        .ZN(n2133) );
  OAI22_X1 U1915 ( .A1(n1564), .A2(n1676), .B1(n1639), .B2(n1677), .ZN(n2134)
         );
  INV_X1 U1916 ( .A(b[6]), .ZN(n1677) );
  INV_X1 U1917 ( .A(n1390), .ZN(n1676) );
  AOI222_X1 U1918 ( .A1(n2135), .A2(n2136), .B1(n2135), .B2(n676), .C1(n676), 
        .C2(n2136), .ZN(n2130) );
  XNOR2_X1 U1919 ( .A(a[2]), .B(n2137), .ZN(n2136) );
  AOI221_X1 U1920 ( .B1(b[7]), .B2(n1561), .C1(b[6]), .C2(n1563), .A(n2138), 
        .ZN(n2137) );
  OAI22_X1 U1921 ( .A1(n1564), .A2(n1672), .B1(n1639), .B2(n1673), .ZN(n2138)
         );
  INV_X1 U1922 ( .A(b[5]), .ZN(n1673) );
  INV_X1 U1923 ( .A(n1391), .ZN(n1672) );
  OAI222_X1 U1924 ( .A1(n2139), .A2(n2140), .B1(n2139), .B2(n2141), .C1(n2141), 
        .C2(n2140), .ZN(n2135) );
  INV_X1 U1925 ( .A(n680), .ZN(n2141) );
  XNOR2_X1 U1926 ( .A(n1742), .B(n2142), .ZN(n2140) );
  AOI221_X1 U1927 ( .B1(b[6]), .B2(n1561), .C1(b[5]), .C2(n1563), .A(n2143), 
        .ZN(n2142) );
  OAI22_X1 U1928 ( .A1(n1564), .A2(n1668), .B1(n1639), .B2(n1669), .ZN(n2143)
         );
  INV_X1 U1929 ( .A(b[4]), .ZN(n1669) );
  INV_X1 U1930 ( .A(n1392), .ZN(n1668) );
  AOI222_X1 U1931 ( .A1(n2144), .A2(n2145), .B1(n2144), .B2(n684), .C1(n684), 
        .C2(n2145), .ZN(n2139) );
  XNOR2_X1 U1932 ( .A(a[2]), .B(n2146), .ZN(n2145) );
  AOI221_X1 U1933 ( .B1(b[5]), .B2(n1561), .C1(b[4]), .C2(n1563), .A(n2147), 
        .ZN(n2146) );
  OAI22_X1 U1934 ( .A1(n1564), .A2(n1664), .B1(n1639), .B2(n1665), .ZN(n2147)
         );
  INV_X1 U1935 ( .A(b[3]), .ZN(n1665) );
  INV_X1 U1936 ( .A(n1393), .ZN(n1664) );
  OAI222_X1 U1937 ( .A1(n2148), .A2(n2149), .B1(n2148), .B2(n2150), .C1(n2150), 
        .C2(n2149), .ZN(n2144) );
  INV_X1 U1938 ( .A(n686), .ZN(n2150) );
  XNOR2_X1 U1939 ( .A(n1742), .B(n2151), .ZN(n2149) );
  AOI221_X1 U1940 ( .B1(b[4]), .B2(n1561), .C1(b[3]), .C2(n1563), .A(n2152), 
        .ZN(n2151) );
  OAI22_X1 U1941 ( .A1(n1564), .A2(n1660), .B1(n1639), .B2(n1661), .ZN(n2152)
         );
  INV_X1 U1942 ( .A(n1394), .ZN(n1660) );
  AOI222_X1 U1943 ( .A1(n2153), .A2(n2154), .B1(n2153), .B2(n688), .C1(n688), 
        .C2(n2154), .ZN(n2148) );
  XNOR2_X1 U1944 ( .A(a[2]), .B(n2155), .ZN(n2154) );
  AOI221_X1 U1945 ( .B1(b[3]), .B2(n1561), .C1(b[2]), .C2(n1563), .A(n2156), 
        .ZN(n2155) );
  OAI22_X1 U1946 ( .A1(n1564), .A2(n1657), .B1(n1639), .B2(n1649), .ZN(n2156)
         );
  INV_X1 U1947 ( .A(b[1]), .ZN(n1649) );
  INV_X1 U1948 ( .A(n1395), .ZN(n1657) );
  AND2_X1 U1949 ( .A1(n2160), .A2(n2161), .ZN(n2153) );
  AOI211_X1 U1950 ( .C1(b[1]), .C2(n1561), .A(n2162), .B(b[0]), .ZN(n2161) );
  OAI22_X1 U1951 ( .A1(n1535), .A2(n1661), .B1(n1564), .B2(n1650), .ZN(n2162)
         );
  INV_X1 U1952 ( .A(n1397), .ZN(n1650) );
  INV_X1 U1953 ( .A(b[2]), .ZN(n1661) );
  INV_X1 U1954 ( .A(a[0]), .ZN(n2158) );
  AOI221_X1 U1955 ( .B1(b[1]), .B2(n1563), .C1(n1396), .C2(n1555), .A(n1742), 
        .ZN(n2160) );
  XNOR2_X1 U1956 ( .A(a[1]), .B(n1742), .ZN(n2157) );
  INV_X1 U1957 ( .A(a[2]), .ZN(n1742) );
  NOR2_X1 U1958 ( .A1(n2159), .A2(a[0]), .ZN(n1636) );
  INV_X1 U1959 ( .A(a[1]), .ZN(n2159) );
endmodule


module iir_filter_DW_mult_tc_0 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(product[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(product[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(product[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(product[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(product[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(product[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(product[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(product[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(product[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(product[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(product[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(product[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(product[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(product[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(product[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(product[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(product[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(product[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(product[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(product[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(product[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(product[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(product[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1598), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1600), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1602), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1604), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1606), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1608), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1610), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(b[22]), .B(n1614), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(b[21]), .B(b[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(b[20]), .B(b[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(b[19]), .B(b[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(b[18]), .B(b[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(b[17]), .B(b[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(b[16]), .B(b[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(b[15]), .B(b[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(b[14]), .B(b[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(b[13]), .B(b[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(b[12]), .B(b[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(b[11]), .B(b[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(b[10]), .B(b[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(b[9]), .B(b[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(b[8]), .B(b[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(b[7]), .B(b[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(b[6]), .B(b[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(b[5]), .B(b[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(b[4]), .B(b[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(b[3]), .B(b[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(b[2]), .B(b[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(b[1]), .B(b[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(b[0]), .B(b[1]), .CO(n727), .S(n1397) );
  INV_X1 U1137 ( .A(n1533), .ZN(n1570) );
  INV_X1 U1138 ( .A(n1536), .ZN(n1568) );
  INV_X1 U1139 ( .A(n1535), .ZN(n1561) );
  INV_X1 U1140 ( .A(n1534), .ZN(n1569) );
  BUF_X1 U1141 ( .A(n1654), .Z(n1572) );
  INV_X1 U1142 ( .A(n1547), .ZN(n1560) );
  INV_X1 U1143 ( .A(n1544), .ZN(n1558) );
  INV_X1 U1144 ( .A(n1537), .ZN(n1580) );
  INV_X1 U1145 ( .A(n1551), .ZN(n1575) );
  INV_X1 U1146 ( .A(n1550), .ZN(n1585) );
  INV_X1 U1147 ( .A(n1548), .ZN(n1595) );
  INV_X1 U1148 ( .A(n1549), .ZN(n1590) );
  INV_X1 U1149 ( .A(n1538), .ZN(n1559) );
  INV_X1 U1150 ( .A(n1545), .ZN(n1593) );
  INV_X1 U1151 ( .A(n1553), .ZN(n1583) );
  INV_X1 U1152 ( .A(n1552), .ZN(n1588) );
  INV_X1 U1153 ( .A(n1546), .ZN(n1578) );
  INV_X1 U1154 ( .A(n1554), .ZN(n1573) );
  BUF_X1 U1155 ( .A(n1654), .Z(n1571) );
  BUF_X1 U1156 ( .A(n1629), .Z(n1557) );
  BUF_X1 U1157 ( .A(n1967), .Z(n1596) );
  BUF_X1 U1158 ( .A(n1912), .Z(n1591) );
  BUF_X1 U1159 ( .A(n1857), .Z(n1586) );
  BUF_X1 U1160 ( .A(n1802), .Z(n1581) );
  BUF_X1 U1161 ( .A(n1747), .Z(n1576) );
  BUF_X1 U1162 ( .A(n1912), .Z(n1592) );
  BUF_X1 U1163 ( .A(n1857), .Z(n1587) );
  BUF_X1 U1164 ( .A(n1802), .Z(n1582) );
  BUF_X1 U1165 ( .A(n1747), .Z(n1577) );
  BUF_X1 U1166 ( .A(n1967), .Z(n1597) );
  INV_X1 U1167 ( .A(n1615), .ZN(n1614) );
  INV_X1 U1168 ( .A(n1540), .ZN(n1589) );
  INV_X1 U1169 ( .A(n1541), .ZN(n1584) );
  INV_X1 U1170 ( .A(n1542), .ZN(n1579) );
  INV_X1 U1171 ( .A(n1543), .ZN(n1574) );
  BUF_X1 U1172 ( .A(n1629), .Z(n1556) );
  INV_X1 U1173 ( .A(n1539), .ZN(n1594) );
  NAND3_X1 U1174 ( .A1(n2157), .A2(n2158), .A3(n2159), .ZN(n1639) );
  INV_X1 U1175 ( .A(n1555), .ZN(n1564) );
  OR2_X1 U1176 ( .A1(n1738), .A2(n1739), .ZN(n1533) );
  OR2_X1 U1177 ( .A1(n1740), .A2(n1741), .ZN(n1534) );
  OR2_X1 U1178 ( .A1(n2158), .A2(n2157), .ZN(n1535) );
  AND2_X1 U1179 ( .A1(n1738), .A2(n1740), .ZN(n1536) );
  INV_X1 U1180 ( .A(n1611), .ZN(n1610) );
  INV_X1 U1181 ( .A(n1607), .ZN(n1606) );
  INV_X1 U1182 ( .A(n1609), .ZN(n1608) );
  INV_X1 U1183 ( .A(n1603), .ZN(n1602) );
  INV_X1 U1184 ( .A(n1605), .ZN(n1604) );
  OR2_X1 U1185 ( .A1(n1849), .A2(n1850), .ZN(n1537) );
  BUF_X1 U1186 ( .A(n1636), .Z(n1562) );
  BUF_X1 U1187 ( .A(n1636), .Z(n1563) );
  BUF_X1 U1188 ( .A(n1647), .Z(n1565) );
  BUF_X1 U1189 ( .A(n1647), .Z(n1566) );
  OR2_X1 U1190 ( .A1(n2068), .A2(n2067), .ZN(n1538) );
  OR2_X1 U1191 ( .A1(n2016), .A2(n2017), .ZN(n1539) );
  OR2_X1 U1192 ( .A1(n1961), .A2(n1962), .ZN(n1540) );
  OR2_X1 U1193 ( .A1(n1906), .A2(n1907), .ZN(n1541) );
  OR2_X1 U1194 ( .A1(n1851), .A2(n1852), .ZN(n1542) );
  OR2_X1 U1195 ( .A1(n1796), .A2(n1797), .ZN(n1543) );
  AND2_X1 U1196 ( .A1(n2070), .A2(n2068), .ZN(n1544) );
  AND2_X1 U1197 ( .A1(n2014), .A2(n2016), .ZN(n1545) );
  AND2_X1 U1198 ( .A1(n1849), .A2(n1851), .ZN(n1546) );
  OR2_X1 U1199 ( .A1(n2070), .A2(n2069), .ZN(n1547) );
  OR2_X1 U1200 ( .A1(n2014), .A2(n2015), .ZN(n1548) );
  OR2_X1 U1201 ( .A1(n1959), .A2(n1960), .ZN(n1549) );
  OR2_X1 U1202 ( .A1(n1904), .A2(n1905), .ZN(n1550) );
  OR2_X1 U1203 ( .A1(n1794), .A2(n1795), .ZN(n1551) );
  AND2_X1 U1204 ( .A1(n1959), .A2(n1961), .ZN(n1552) );
  AND2_X1 U1205 ( .A1(n1904), .A2(n1906), .ZN(n1553) );
  AND2_X1 U1206 ( .A1(n1794), .A2(n1796), .ZN(n1554) );
  BUF_X1 U1207 ( .A(n1647), .Z(n1567) );
  INV_X1 U1208 ( .A(n1599), .ZN(n1598) );
  AND2_X1 U1209 ( .A1(a[0]), .A2(n2157), .ZN(n1555) );
  BUF_X1 U1210 ( .A(a[20]), .Z(n1600) );
  INV_X1 U1211 ( .A(a[23]), .ZN(n1599) );
  INV_X1 U1212 ( .A(a[5]), .ZN(n1611) );
  INV_X1 U1213 ( .A(a[11]), .ZN(n1607) );
  INV_X1 U1214 ( .A(a[8]), .ZN(n1609) );
  INV_X1 U1215 ( .A(a[17]), .ZN(n1603) );
  INV_X1 U1216 ( .A(a[14]), .ZN(n1605) );
  BUF_X1 U1217 ( .A(a[20]), .Z(n1601) );
  CLKBUF_X1 U1218 ( .A(b[23]), .Z(n1612) );
  CLKBUF_X1 U1219 ( .A(b[23]), .Z(n1613) );
  INV_X1 U1220 ( .A(b[23]), .ZN(n1615) );
  INV_X1 U1221 ( .A(n1612), .ZN(n1616) );
  INV_X1 U1222 ( .A(n1612), .ZN(n1617) );
  INV_X1 U1223 ( .A(n1612), .ZN(n1618) );
  INV_X1 U1224 ( .A(n1613), .ZN(n1619) );
  INV_X1 U1225 ( .A(n1613), .ZN(n1620) );
  AOI21_X1 U1226 ( .B1(n1621), .B2(n1622), .A(n1623), .ZN(product[47]) );
  OAI22_X1 U1227 ( .A1(n1624), .A2(n1625), .B1(n1624), .B2(n1626), .ZN(n1623)
         );
  INV_X1 U1228 ( .A(n1622), .ZN(n1626) );
  AOI222_X1 U1229 ( .A1(n1627), .A2(n303), .B1(n1625), .B2(n303), .C1(n1627), 
        .C2(n1625), .ZN(n1624) );
  XOR2_X1 U1230 ( .A(n1628), .B(n1599), .Z(n1622) );
  OAI221_X1 U1231 ( .B1(n1617), .B2(n1557), .C1(n1620), .C2(n1558), .A(n1630), 
        .ZN(n1628) );
  OAI21_X1 U1232 ( .B1(n1559), .B2(n1560), .A(n1614), .ZN(n1630) );
  INV_X1 U1233 ( .A(n1625), .ZN(n1621) );
  XOR2_X1 U1234 ( .A(a[23]), .B(n1631), .Z(n1625) );
  AOI221_X1 U1235 ( .B1(n1613), .B2(n1559), .C1(n1560), .C2(n1614), .A(n1632), 
        .ZN(n1631) );
  OAI22_X1 U1236 ( .A1(n1558), .A2(n1633), .B1(n1557), .B2(n1634), .ZN(n1632)
         );
  XNOR2_X1 U1237 ( .A(a[2]), .B(n1635), .ZN(n908) );
  AOI221_X1 U1238 ( .B1(n1561), .B2(b[22]), .C1(n1563), .C2(b[21]), .A(n1637), 
        .ZN(n1635) );
  OAI22_X1 U1239 ( .A1(n1564), .A2(n1638), .B1(n1639), .B2(n1640), .ZN(n1637)
         );
  INV_X1 U1240 ( .A(n1376), .ZN(n1638) );
  XNOR2_X1 U1241 ( .A(a[2]), .B(n1641), .ZN(n907) );
  AOI221_X1 U1242 ( .B1(n1563), .B2(b[22]), .C1(n1555), .C2(n1375), .A(n1642), 
        .ZN(n1641) );
  OAI22_X1 U1243 ( .A1(n1643), .A2(n1639), .B1(n1617), .B2(n1535), .ZN(n1642)
         );
  XNOR2_X1 U1244 ( .A(a[2]), .B(n1644), .ZN(n906) );
  AOI221_X1 U1245 ( .B1(n1561), .B2(n1613), .C1(n1563), .C2(n1614), .A(n1645), 
        .ZN(n1644) );
  OAI22_X1 U1246 ( .A1(n1633), .A2(n1564), .B1(n1634), .B2(n1639), .ZN(n1645)
         );
  XNOR2_X1 U1247 ( .A(n1646), .B(n1611), .ZN(n904) );
  OAI22_X1 U1248 ( .A1(n1565), .A2(n1534), .B1(n1568), .B2(n1567), .ZN(n1646)
         );
  XNOR2_X1 U1249 ( .A(n1648), .B(n1611), .ZN(n903) );
  OAI222_X1 U1250 ( .A1(n1534), .A2(n1649), .B1(n1566), .B2(n1533), .C1(n1568), 
        .C2(n1650), .ZN(n1648) );
  XNOR2_X1 U1251 ( .A(n1610), .B(n1651), .ZN(n902) );
  AOI221_X1 U1252 ( .B1(b[2]), .B2(n1569), .C1(b[1]), .C2(n1570), .A(n1652), 
        .ZN(n1651) );
  OAI22_X1 U1253 ( .A1(n1568), .A2(n1653), .B1(n1565), .B2(n1572), .ZN(n1652)
         );
  XNOR2_X1 U1254 ( .A(n1610), .B(n1655), .ZN(n901) );
  AOI221_X1 U1255 ( .B1(b[3]), .B2(n1569), .C1(b[2]), .C2(n1570), .A(n1656), 
        .ZN(n1655) );
  OAI22_X1 U1256 ( .A1(n1568), .A2(n1657), .B1(n1649), .B2(n1572), .ZN(n1656)
         );
  XNOR2_X1 U1257 ( .A(n1610), .B(n1658), .ZN(n900) );
  AOI221_X1 U1258 ( .B1(b[4]), .B2(n1569), .C1(b[3]), .C2(n1570), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1259 ( .A1(n1568), .A2(n1660), .B1(n1661), .B2(n1572), .ZN(n1659)
         );
  XNOR2_X1 U1260 ( .A(n1610), .B(n1662), .ZN(n899) );
  AOI221_X1 U1261 ( .B1(b[5]), .B2(n1569), .C1(b[4]), .C2(n1570), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1262 ( .A1(n1568), .A2(n1664), .B1(n1572), .B2(n1665), .ZN(n1663)
         );
  XNOR2_X1 U1263 ( .A(n1610), .B(n1666), .ZN(n898) );
  AOI221_X1 U1264 ( .B1(b[6]), .B2(n1569), .C1(b[5]), .C2(n1570), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1265 ( .A1(n1568), .A2(n1668), .B1(n1572), .B2(n1669), .ZN(n1667)
         );
  XNOR2_X1 U1266 ( .A(n1610), .B(n1670), .ZN(n897) );
  AOI221_X1 U1267 ( .B1(b[7]), .B2(n1569), .C1(b[6]), .C2(n1570), .A(n1671), 
        .ZN(n1670) );
  OAI22_X1 U1268 ( .A1(n1568), .A2(n1672), .B1(n1572), .B2(n1673), .ZN(n1671)
         );
  XNOR2_X1 U1269 ( .A(n1610), .B(n1674), .ZN(n896) );
  AOI221_X1 U1270 ( .B1(b[8]), .B2(n1569), .C1(b[7]), .C2(n1570), .A(n1675), 
        .ZN(n1674) );
  OAI22_X1 U1271 ( .A1(n1568), .A2(n1676), .B1(n1571), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1272 ( .A(n1610), .B(n1678), .ZN(n895) );
  AOI221_X1 U1273 ( .B1(b[9]), .B2(n1569), .C1(b[8]), .C2(n1570), .A(n1679), 
        .ZN(n1678) );
  OAI22_X1 U1274 ( .A1(n1568), .A2(n1680), .B1(n1572), .B2(n1681), .ZN(n1679)
         );
  XNOR2_X1 U1275 ( .A(n1610), .B(n1682), .ZN(n894) );
  AOI221_X1 U1276 ( .B1(b[10]), .B2(n1569), .C1(b[9]), .C2(n1570), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1277 ( .A1(n1568), .A2(n1684), .B1(n1572), .B2(n1685), .ZN(n1683)
         );
  XNOR2_X1 U1278 ( .A(n1610), .B(n1686), .ZN(n893) );
  AOI221_X1 U1279 ( .B1(b[11]), .B2(n1569), .C1(b[10]), .C2(n1570), .A(n1687), 
        .ZN(n1686) );
  OAI22_X1 U1280 ( .A1(n1568), .A2(n1688), .B1(n1571), .B2(n1689), .ZN(n1687)
         );
  XNOR2_X1 U1281 ( .A(n1610), .B(n1690), .ZN(n892) );
  AOI221_X1 U1282 ( .B1(b[12]), .B2(n1569), .C1(b[11]), .C2(n1570), .A(n1691), 
        .ZN(n1690) );
  OAI22_X1 U1283 ( .A1(n1568), .A2(n1692), .B1(n1571), .B2(n1693), .ZN(n1691)
         );
  XNOR2_X1 U1284 ( .A(n1610), .B(n1694), .ZN(n891) );
  AOI221_X1 U1285 ( .B1(b[13]), .B2(n1569), .C1(b[12]), .C2(n1570), .A(n1695), 
        .ZN(n1694) );
  OAI22_X1 U1286 ( .A1(n1568), .A2(n1696), .B1(n1571), .B2(n1697), .ZN(n1695)
         );
  XNOR2_X1 U1287 ( .A(n1610), .B(n1698), .ZN(n890) );
  AOI221_X1 U1288 ( .B1(b[14]), .B2(n1569), .C1(b[13]), .C2(n1570), .A(n1699), 
        .ZN(n1698) );
  OAI22_X1 U1289 ( .A1(n1568), .A2(n1700), .B1(n1571), .B2(n1701), .ZN(n1699)
         );
  XNOR2_X1 U1290 ( .A(n1610), .B(n1702), .ZN(n889) );
  AOI221_X1 U1291 ( .B1(b[15]), .B2(n1569), .C1(b[14]), .C2(n1570), .A(n1703), 
        .ZN(n1702) );
  OAI22_X1 U1292 ( .A1(n1568), .A2(n1704), .B1(n1571), .B2(n1705), .ZN(n1703)
         );
  XNOR2_X1 U1293 ( .A(n1610), .B(n1706), .ZN(n888) );
  AOI221_X1 U1294 ( .B1(b[16]), .B2(n1569), .C1(b[15]), .C2(n1570), .A(n1707), 
        .ZN(n1706) );
  OAI22_X1 U1295 ( .A1(n1568), .A2(n1708), .B1(n1571), .B2(n1709), .ZN(n1707)
         );
  XNOR2_X1 U1296 ( .A(n1610), .B(n1710), .ZN(n887) );
  AOI221_X1 U1297 ( .B1(b[17]), .B2(n1569), .C1(b[16]), .C2(n1570), .A(n1711), 
        .ZN(n1710) );
  OAI22_X1 U1298 ( .A1(n1568), .A2(n1712), .B1(n1571), .B2(n1713), .ZN(n1711)
         );
  XNOR2_X1 U1299 ( .A(n1610), .B(n1714), .ZN(n886) );
  AOI221_X1 U1300 ( .B1(b[18]), .B2(n1569), .C1(b[17]), .C2(n1570), .A(n1715), 
        .ZN(n1714) );
  OAI22_X1 U1301 ( .A1(n1568), .A2(n1716), .B1(n1571), .B2(n1717), .ZN(n1715)
         );
  XNOR2_X1 U1302 ( .A(n1610), .B(n1718), .ZN(n885) );
  AOI221_X1 U1303 ( .B1(b[19]), .B2(n1569), .C1(b[18]), .C2(n1570), .A(n1719), 
        .ZN(n1718) );
  OAI22_X1 U1304 ( .A1(n1568), .A2(n1720), .B1(n1571), .B2(n1721), .ZN(n1719)
         );
  XNOR2_X1 U1305 ( .A(a[5]), .B(n1722), .ZN(n884) );
  AOI221_X1 U1306 ( .B1(n1569), .B2(b[20]), .C1(b[19]), .C2(n1570), .A(n1723), 
        .ZN(n1722) );
  OAI22_X1 U1307 ( .A1(n1568), .A2(n1724), .B1(n1571), .B2(n1725), .ZN(n1723)
         );
  XNOR2_X1 U1308 ( .A(a[5]), .B(n1726), .ZN(n883) );
  AOI221_X1 U1309 ( .B1(n1569), .B2(b[21]), .C1(n1570), .C2(b[20]), .A(n1727), 
        .ZN(n1726) );
  OAI22_X1 U1310 ( .A1(n1568), .A2(n1728), .B1(n1571), .B2(n1729), .ZN(n1727)
         );
  XNOR2_X1 U1311 ( .A(a[5]), .B(n1730), .ZN(n882) );
  AOI221_X1 U1312 ( .B1(n1569), .B2(b[22]), .C1(n1536), .C2(n1376), .A(n1731), 
        .ZN(n1730) );
  OAI22_X1 U1313 ( .A1(n1640), .A2(n1572), .B1(n1643), .B2(n1533), .ZN(n1731)
         );
  XNOR2_X1 U1314 ( .A(a[5]), .B(n1732), .ZN(n881) );
  AOI221_X1 U1315 ( .B1(n1570), .B2(b[22]), .C1(n1536), .C2(n1375), .A(n1733), 
        .ZN(n1732) );
  OAI22_X1 U1316 ( .A1(n1615), .A2(n1534), .B1(n1643), .B2(n1572), .ZN(n1733)
         );
  XNOR2_X1 U1317 ( .A(a[5]), .B(n1734), .ZN(n880) );
  AOI221_X1 U1318 ( .B1(n1569), .B2(n1613), .C1(n1570), .C2(n1614), .A(n1735), 
        .ZN(n1734) );
  OAI22_X1 U1319 ( .A1(n1633), .A2(n1568), .B1(n1634), .B2(n1572), .ZN(n1735)
         );
  XNOR2_X1 U1320 ( .A(n1610), .B(n1736), .ZN(n879) );
  OAI221_X1 U1321 ( .B1(n1616), .B2(n1572), .C1(n1620), .C2(n1568), .A(n1737), 
        .ZN(n1736) );
  OAI21_X1 U1322 ( .B1(n1569), .B2(n1570), .A(n1614), .ZN(n1737) );
  INV_X1 U1323 ( .A(n1741), .ZN(n1738) );
  NAND3_X1 U1324 ( .A1(n1741), .A2(n1740), .A3(n1739), .ZN(n1654) );
  XNOR2_X1 U1325 ( .A(a[3]), .B(a[4]), .ZN(n1739) );
  XNOR2_X1 U1326 ( .A(a[4]), .B(n1611), .ZN(n1740) );
  XOR2_X1 U1327 ( .A(a[3]), .B(n1742), .Z(n1741) );
  XNOR2_X1 U1328 ( .A(n1743), .B(n1609), .ZN(n878) );
  OAI22_X1 U1329 ( .A1(n1565), .A2(n1543), .B1(n1565), .B2(n1573), .ZN(n1743)
         );
  XNOR2_X1 U1330 ( .A(n1744), .B(n1609), .ZN(n877) );
  OAI222_X1 U1331 ( .A1(n1649), .A2(n1543), .B1(n1566), .B2(n1551), .C1(n1650), 
        .C2(n1573), .ZN(n1744) );
  XNOR2_X1 U1332 ( .A(n1608), .B(n1745), .ZN(n876) );
  AOI221_X1 U1333 ( .B1(n1574), .B2(b[2]), .C1(n1575), .C2(b[1]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1334 ( .A1(n1653), .A2(n1573), .B1(n1565), .B2(n1576), .ZN(n1746)
         );
  XNOR2_X1 U1335 ( .A(n1608), .B(n1748), .ZN(n875) );
  AOI221_X1 U1336 ( .B1(n1574), .B2(b[3]), .C1(n1575), .C2(b[2]), .A(n1749), 
        .ZN(n1748) );
  OAI22_X1 U1337 ( .A1(n1657), .A2(n1573), .B1(n1649), .B2(n1577), .ZN(n1749)
         );
  XNOR2_X1 U1338 ( .A(n1608), .B(n1750), .ZN(n874) );
  AOI221_X1 U1339 ( .B1(n1574), .B2(b[4]), .C1(n1575), .C2(b[3]), .A(n1751), 
        .ZN(n1750) );
  OAI22_X1 U1340 ( .A1(n1660), .A2(n1573), .B1(n1661), .B2(n1577), .ZN(n1751)
         );
  XNOR2_X1 U1341 ( .A(n1608), .B(n1752), .ZN(n873) );
  AOI221_X1 U1342 ( .B1(n1574), .B2(b[5]), .C1(n1575), .C2(b[4]), .A(n1753), 
        .ZN(n1752) );
  OAI22_X1 U1343 ( .A1(n1664), .A2(n1573), .B1(n1665), .B2(n1577), .ZN(n1753)
         );
  XNOR2_X1 U1344 ( .A(n1608), .B(n1754), .ZN(n872) );
  AOI221_X1 U1345 ( .B1(n1574), .B2(b[6]), .C1(n1575), .C2(b[5]), .A(n1755), 
        .ZN(n1754) );
  OAI22_X1 U1346 ( .A1(n1668), .A2(n1573), .B1(n1669), .B2(n1577), .ZN(n1755)
         );
  XNOR2_X1 U1347 ( .A(n1608), .B(n1756), .ZN(n871) );
  AOI221_X1 U1348 ( .B1(n1574), .B2(b[7]), .C1(n1575), .C2(b[6]), .A(n1757), 
        .ZN(n1756) );
  OAI22_X1 U1349 ( .A1(n1672), .A2(n1573), .B1(n1673), .B2(n1577), .ZN(n1757)
         );
  XNOR2_X1 U1350 ( .A(n1608), .B(n1758), .ZN(n870) );
  AOI221_X1 U1351 ( .B1(n1574), .B2(b[8]), .C1(n1575), .C2(b[7]), .A(n1759), 
        .ZN(n1758) );
  OAI22_X1 U1352 ( .A1(n1676), .A2(n1573), .B1(n1677), .B2(n1577), .ZN(n1759)
         );
  XNOR2_X1 U1353 ( .A(n1608), .B(n1760), .ZN(n869) );
  AOI221_X1 U1354 ( .B1(n1574), .B2(b[9]), .C1(n1575), .C2(b[8]), .A(n1761), 
        .ZN(n1760) );
  OAI22_X1 U1355 ( .A1(n1680), .A2(n1573), .B1(n1681), .B2(n1577), .ZN(n1761)
         );
  XNOR2_X1 U1356 ( .A(n1608), .B(n1762), .ZN(n868) );
  AOI221_X1 U1357 ( .B1(n1574), .B2(b[10]), .C1(n1575), .C2(b[9]), .A(n1763), 
        .ZN(n1762) );
  OAI22_X1 U1358 ( .A1(n1684), .A2(n1573), .B1(n1685), .B2(n1577), .ZN(n1763)
         );
  XNOR2_X1 U1359 ( .A(n1608), .B(n1764), .ZN(n867) );
  AOI221_X1 U1360 ( .B1(n1574), .B2(b[11]), .C1(n1575), .C2(b[10]), .A(n1765), 
        .ZN(n1764) );
  OAI22_X1 U1361 ( .A1(n1688), .A2(n1573), .B1(n1689), .B2(n1577), .ZN(n1765)
         );
  XNOR2_X1 U1362 ( .A(n1608), .B(n1766), .ZN(n866) );
  AOI221_X1 U1363 ( .B1(n1574), .B2(b[12]), .C1(n1575), .C2(b[11]), .A(n1767), 
        .ZN(n1766) );
  OAI22_X1 U1364 ( .A1(n1692), .A2(n1573), .B1(n1693), .B2(n1577), .ZN(n1767)
         );
  XNOR2_X1 U1365 ( .A(n1608), .B(n1768), .ZN(n865) );
  AOI221_X1 U1366 ( .B1(n1574), .B2(b[13]), .C1(n1575), .C2(b[12]), .A(n1769), 
        .ZN(n1768) );
  OAI22_X1 U1367 ( .A1(n1696), .A2(n1573), .B1(n1697), .B2(n1576), .ZN(n1769)
         );
  XNOR2_X1 U1368 ( .A(n1608), .B(n1770), .ZN(n864) );
  AOI221_X1 U1369 ( .B1(n1574), .B2(b[14]), .C1(n1575), .C2(b[13]), .A(n1771), 
        .ZN(n1770) );
  OAI22_X1 U1370 ( .A1(n1700), .A2(n1573), .B1(n1701), .B2(n1576), .ZN(n1771)
         );
  XNOR2_X1 U1371 ( .A(n1608), .B(n1772), .ZN(n863) );
  AOI221_X1 U1372 ( .B1(n1574), .B2(b[15]), .C1(n1575), .C2(b[14]), .A(n1773), 
        .ZN(n1772) );
  OAI22_X1 U1373 ( .A1(n1704), .A2(n1573), .B1(n1705), .B2(n1576), .ZN(n1773)
         );
  XNOR2_X1 U1374 ( .A(n1608), .B(n1774), .ZN(n862) );
  AOI221_X1 U1375 ( .B1(n1574), .B2(b[16]), .C1(n1575), .C2(b[15]), .A(n1775), 
        .ZN(n1774) );
  OAI22_X1 U1376 ( .A1(n1708), .A2(n1573), .B1(n1709), .B2(n1576), .ZN(n1775)
         );
  XNOR2_X1 U1377 ( .A(n1608), .B(n1776), .ZN(n861) );
  AOI221_X1 U1378 ( .B1(n1574), .B2(b[17]), .C1(n1575), .C2(b[16]), .A(n1777), 
        .ZN(n1776) );
  OAI22_X1 U1379 ( .A1(n1712), .A2(n1573), .B1(n1713), .B2(n1576), .ZN(n1777)
         );
  XNOR2_X1 U1380 ( .A(n1608), .B(n1778), .ZN(n860) );
  AOI221_X1 U1381 ( .B1(n1574), .B2(b[18]), .C1(n1575), .C2(b[17]), .A(n1779), 
        .ZN(n1778) );
  OAI22_X1 U1382 ( .A1(n1716), .A2(n1573), .B1(n1717), .B2(n1576), .ZN(n1779)
         );
  XNOR2_X1 U1383 ( .A(n1608), .B(n1780), .ZN(n859) );
  AOI221_X1 U1384 ( .B1(n1574), .B2(b[19]), .C1(n1575), .C2(b[18]), .A(n1781), 
        .ZN(n1780) );
  OAI22_X1 U1385 ( .A1(n1720), .A2(n1573), .B1(n1721), .B2(n1576), .ZN(n1781)
         );
  XNOR2_X1 U1386 ( .A(a[8]), .B(n1782), .ZN(n858) );
  AOI221_X1 U1387 ( .B1(n1574), .B2(b[20]), .C1(n1575), .C2(b[19]), .A(n1783), 
        .ZN(n1782) );
  OAI22_X1 U1388 ( .A1(n1724), .A2(n1573), .B1(n1725), .B2(n1576), .ZN(n1783)
         );
  XNOR2_X1 U1389 ( .A(a[8]), .B(n1784), .ZN(n857) );
  AOI221_X1 U1390 ( .B1(n1574), .B2(b[21]), .C1(n1575), .C2(b[20]), .A(n1785), 
        .ZN(n1784) );
  OAI22_X1 U1391 ( .A1(n1728), .A2(n1573), .B1(n1729), .B2(n1576), .ZN(n1785)
         );
  XNOR2_X1 U1392 ( .A(a[8]), .B(n1786), .ZN(n856) );
  AOI221_X1 U1393 ( .B1(n1574), .B2(b[22]), .C1(n1554), .C2(n1376), .A(n1787), 
        .ZN(n1786) );
  OAI22_X1 U1394 ( .A1(n1640), .A2(n1577), .B1(n1643), .B2(n1551), .ZN(n1787)
         );
  XNOR2_X1 U1395 ( .A(a[8]), .B(n1788), .ZN(n855) );
  AOI221_X1 U1396 ( .B1(n1575), .B2(b[22]), .C1(n1554), .C2(n1375), .A(n1789), 
        .ZN(n1788) );
  OAI22_X1 U1397 ( .A1(n1617), .A2(n1543), .B1(n1643), .B2(n1576), .ZN(n1789)
         );
  XNOR2_X1 U1398 ( .A(a[8]), .B(n1790), .ZN(n854) );
  AOI221_X1 U1399 ( .B1(n1574), .B2(n1613), .C1(n1575), .C2(n1614), .A(n1791), 
        .ZN(n1790) );
  OAI22_X1 U1400 ( .A1(n1633), .A2(n1573), .B1(n1634), .B2(n1576), .ZN(n1791)
         );
  XNOR2_X1 U1401 ( .A(n1608), .B(n1792), .ZN(n853) );
  OAI221_X1 U1402 ( .B1(n1616), .B2(n1577), .C1(n1617), .C2(n1573), .A(n1793), 
        .ZN(n1792) );
  OAI21_X1 U1403 ( .B1(n1574), .B2(n1575), .A(n1614), .ZN(n1793) );
  INV_X1 U1404 ( .A(n1797), .ZN(n1794) );
  NAND3_X1 U1405 ( .A1(n1797), .A2(n1796), .A3(n1795), .ZN(n1747) );
  XNOR2_X1 U1406 ( .A(a[6]), .B(a[7]), .ZN(n1795) );
  XNOR2_X1 U1407 ( .A(a[7]), .B(n1609), .ZN(n1796) );
  XOR2_X1 U1408 ( .A(a[6]), .B(n1611), .Z(n1797) );
  XNOR2_X1 U1409 ( .A(n1798), .B(n1607), .ZN(n852) );
  OAI22_X1 U1410 ( .A1(n1565), .A2(n1542), .B1(n1565), .B2(n1578), .ZN(n1798)
         );
  XNOR2_X1 U1411 ( .A(n1799), .B(n1607), .ZN(n851) );
  OAI222_X1 U1412 ( .A1(n1649), .A2(n1542), .B1(n1566), .B2(n1537), .C1(n1650), 
        .C2(n1578), .ZN(n1799) );
  XNOR2_X1 U1413 ( .A(n1606), .B(n1800), .ZN(n850) );
  AOI221_X1 U1414 ( .B1(n1579), .B2(b[2]), .C1(n1580), .C2(b[1]), .A(n1801), 
        .ZN(n1800) );
  OAI22_X1 U1415 ( .A1(n1653), .A2(n1578), .B1(n1566), .B2(n1581), .ZN(n1801)
         );
  XNOR2_X1 U1416 ( .A(n1606), .B(n1803), .ZN(n849) );
  AOI221_X1 U1417 ( .B1(n1579), .B2(b[3]), .C1(n1580), .C2(b[2]), .A(n1804), 
        .ZN(n1803) );
  OAI22_X1 U1418 ( .A1(n1657), .A2(n1578), .B1(n1649), .B2(n1582), .ZN(n1804)
         );
  XNOR2_X1 U1419 ( .A(n1606), .B(n1805), .ZN(n848) );
  AOI221_X1 U1420 ( .B1(n1579), .B2(b[4]), .C1(n1580), .C2(b[3]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1421 ( .A1(n1660), .A2(n1578), .B1(n1661), .B2(n1582), .ZN(n1806)
         );
  XNOR2_X1 U1422 ( .A(n1606), .B(n1807), .ZN(n847) );
  AOI221_X1 U1423 ( .B1(n1579), .B2(b[5]), .C1(n1580), .C2(b[4]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1424 ( .A1(n1664), .A2(n1578), .B1(n1665), .B2(n1582), .ZN(n1808)
         );
  XNOR2_X1 U1425 ( .A(n1606), .B(n1809), .ZN(n846) );
  AOI221_X1 U1426 ( .B1(n1579), .B2(b[6]), .C1(n1580), .C2(b[5]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1427 ( .A1(n1668), .A2(n1578), .B1(n1669), .B2(n1582), .ZN(n1810)
         );
  XNOR2_X1 U1428 ( .A(n1606), .B(n1811), .ZN(n845) );
  AOI221_X1 U1429 ( .B1(n1579), .B2(b[7]), .C1(n1580), .C2(b[6]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1430 ( .A1(n1672), .A2(n1578), .B1(n1673), .B2(n1582), .ZN(n1812)
         );
  XNOR2_X1 U1431 ( .A(n1606), .B(n1813), .ZN(n844) );
  AOI221_X1 U1432 ( .B1(n1579), .B2(b[8]), .C1(n1580), .C2(b[7]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1433 ( .A1(n1676), .A2(n1578), .B1(n1677), .B2(n1582), .ZN(n1814)
         );
  XNOR2_X1 U1434 ( .A(n1606), .B(n1815), .ZN(n843) );
  AOI221_X1 U1435 ( .B1(n1579), .B2(b[9]), .C1(n1580), .C2(b[8]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1436 ( .A1(n1680), .A2(n1578), .B1(n1681), .B2(n1582), .ZN(n1816)
         );
  XNOR2_X1 U1437 ( .A(n1606), .B(n1817), .ZN(n842) );
  AOI221_X1 U1438 ( .B1(n1579), .B2(b[10]), .C1(n1580), .C2(b[9]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1439 ( .A1(n1684), .A2(n1578), .B1(n1685), .B2(n1582), .ZN(n1818)
         );
  XNOR2_X1 U1440 ( .A(n1606), .B(n1819), .ZN(n841) );
  AOI221_X1 U1441 ( .B1(n1579), .B2(b[11]), .C1(n1580), .C2(b[10]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1442 ( .A1(n1688), .A2(n1578), .B1(n1689), .B2(n1582), .ZN(n1820)
         );
  XNOR2_X1 U1443 ( .A(n1606), .B(n1821), .ZN(n840) );
  AOI221_X1 U1444 ( .B1(n1579), .B2(b[12]), .C1(n1580), .C2(b[11]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1445 ( .A1(n1692), .A2(n1578), .B1(n1693), .B2(n1582), .ZN(n1822)
         );
  XNOR2_X1 U1446 ( .A(n1606), .B(n1823), .ZN(n839) );
  AOI221_X1 U1447 ( .B1(n1579), .B2(b[13]), .C1(n1580), .C2(b[12]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1448 ( .A1(n1696), .A2(n1578), .B1(n1697), .B2(n1581), .ZN(n1824)
         );
  XNOR2_X1 U1449 ( .A(n1606), .B(n1825), .ZN(n838) );
  AOI221_X1 U1450 ( .B1(n1579), .B2(b[14]), .C1(n1580), .C2(b[13]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1451 ( .A1(n1700), .A2(n1578), .B1(n1701), .B2(n1581), .ZN(n1826)
         );
  XNOR2_X1 U1452 ( .A(n1606), .B(n1827), .ZN(n837) );
  AOI221_X1 U1453 ( .B1(n1579), .B2(b[15]), .C1(n1580), .C2(b[14]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1454 ( .A1(n1704), .A2(n1578), .B1(n1705), .B2(n1581), .ZN(n1828)
         );
  XNOR2_X1 U1455 ( .A(n1606), .B(n1829), .ZN(n836) );
  AOI221_X1 U1456 ( .B1(n1579), .B2(b[16]), .C1(n1580), .C2(b[15]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1457 ( .A1(n1708), .A2(n1578), .B1(n1709), .B2(n1581), .ZN(n1830)
         );
  XNOR2_X1 U1458 ( .A(n1606), .B(n1831), .ZN(n835) );
  AOI221_X1 U1459 ( .B1(n1579), .B2(b[17]), .C1(n1580), .C2(b[16]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1460 ( .A1(n1712), .A2(n1578), .B1(n1713), .B2(n1581), .ZN(n1832)
         );
  XNOR2_X1 U1461 ( .A(n1606), .B(n1833), .ZN(n834) );
  AOI221_X1 U1462 ( .B1(n1579), .B2(b[18]), .C1(n1580), .C2(b[17]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1463 ( .A1(n1716), .A2(n1578), .B1(n1717), .B2(n1581), .ZN(n1834)
         );
  XNOR2_X1 U1464 ( .A(n1606), .B(n1835), .ZN(n833) );
  AOI221_X1 U1465 ( .B1(n1579), .B2(b[19]), .C1(n1580), .C2(b[18]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1466 ( .A1(n1720), .A2(n1578), .B1(n1721), .B2(n1581), .ZN(n1836)
         );
  XNOR2_X1 U1467 ( .A(n1606), .B(n1837), .ZN(n832) );
  AOI221_X1 U1468 ( .B1(n1579), .B2(b[20]), .C1(n1580), .C2(b[19]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1469 ( .A1(n1724), .A2(n1578), .B1(n1725), .B2(n1581), .ZN(n1838)
         );
  XNOR2_X1 U1470 ( .A(a[11]), .B(n1839), .ZN(n831) );
  AOI221_X1 U1471 ( .B1(n1579), .B2(b[21]), .C1(n1580), .C2(b[20]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1472 ( .A1(n1728), .A2(n1578), .B1(n1729), .B2(n1581), .ZN(n1840)
         );
  XNOR2_X1 U1473 ( .A(a[11]), .B(n1841), .ZN(n830) );
  AOI221_X1 U1474 ( .B1(n1579), .B2(b[22]), .C1(n1546), .C2(n1376), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1475 ( .A1(n1640), .A2(n1582), .B1(n1643), .B2(n1537), .ZN(n1842)
         );
  XNOR2_X1 U1476 ( .A(a[11]), .B(n1843), .ZN(n829) );
  AOI221_X1 U1477 ( .B1(n1580), .B2(b[22]), .C1(n1546), .C2(n1375), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1478 ( .A1(n1617), .A2(n1542), .B1(n1643), .B2(n1581), .ZN(n1844)
         );
  XNOR2_X1 U1479 ( .A(a[11]), .B(n1845), .ZN(n828) );
  AOI221_X1 U1480 ( .B1(n1579), .B2(n1614), .C1(n1580), .C2(n1614), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1481 ( .A1(n1633), .A2(n1578), .B1(n1634), .B2(n1581), .ZN(n1846)
         );
  XNOR2_X1 U1482 ( .A(a[11]), .B(n1847), .ZN(n827) );
  OAI221_X1 U1483 ( .B1(n1616), .B2(n1582), .C1(n1617), .C2(n1578), .A(n1848), 
        .ZN(n1847) );
  OAI21_X1 U1484 ( .B1(n1579), .B2(n1580), .A(n1614), .ZN(n1848) );
  INV_X1 U1485 ( .A(n1852), .ZN(n1849) );
  NAND3_X1 U1486 ( .A1(n1852), .A2(n1851), .A3(n1850), .ZN(n1802) );
  XNOR2_X1 U1487 ( .A(a[10]), .B(a[9]), .ZN(n1850) );
  XNOR2_X1 U1488 ( .A(a[10]), .B(n1607), .ZN(n1851) );
  XOR2_X1 U1489 ( .A(a[9]), .B(n1609), .Z(n1852) );
  XNOR2_X1 U1490 ( .A(n1853), .B(n1605), .ZN(n826) );
  OAI22_X1 U1491 ( .A1(n1565), .A2(n1541), .B1(n1565), .B2(n1583), .ZN(n1853)
         );
  XNOR2_X1 U1492 ( .A(n1854), .B(n1605), .ZN(n825) );
  OAI222_X1 U1493 ( .A1(n1649), .A2(n1541), .B1(n1566), .B2(n1550), .C1(n1650), 
        .C2(n1583), .ZN(n1854) );
  XNOR2_X1 U1494 ( .A(n1604), .B(n1855), .ZN(n824) );
  AOI221_X1 U1495 ( .B1(n1584), .B2(b[2]), .C1(n1585), .C2(b[1]), .A(n1856), 
        .ZN(n1855) );
  OAI22_X1 U1496 ( .A1(n1653), .A2(n1583), .B1(n1565), .B2(n1586), .ZN(n1856)
         );
  XNOR2_X1 U1497 ( .A(n1604), .B(n1858), .ZN(n823) );
  AOI221_X1 U1498 ( .B1(n1584), .B2(b[3]), .C1(n1585), .C2(b[2]), .A(n1859), 
        .ZN(n1858) );
  OAI22_X1 U1499 ( .A1(n1657), .A2(n1583), .B1(n1649), .B2(n1587), .ZN(n1859)
         );
  XNOR2_X1 U1500 ( .A(n1604), .B(n1860), .ZN(n822) );
  AOI221_X1 U1501 ( .B1(n1584), .B2(b[4]), .C1(n1585), .C2(b[3]), .A(n1861), 
        .ZN(n1860) );
  OAI22_X1 U1502 ( .A1(n1660), .A2(n1583), .B1(n1661), .B2(n1587), .ZN(n1861)
         );
  XNOR2_X1 U1503 ( .A(n1604), .B(n1862), .ZN(n821) );
  AOI221_X1 U1504 ( .B1(n1584), .B2(b[5]), .C1(n1585), .C2(b[4]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1505 ( .A1(n1664), .A2(n1583), .B1(n1665), .B2(n1587), .ZN(n1863)
         );
  XNOR2_X1 U1506 ( .A(n1604), .B(n1864), .ZN(n820) );
  AOI221_X1 U1507 ( .B1(n1584), .B2(b[6]), .C1(n1585), .C2(b[5]), .A(n1865), 
        .ZN(n1864) );
  OAI22_X1 U1508 ( .A1(n1668), .A2(n1583), .B1(n1669), .B2(n1587), .ZN(n1865)
         );
  XNOR2_X1 U1509 ( .A(n1604), .B(n1866), .ZN(n819) );
  AOI221_X1 U1510 ( .B1(n1584), .B2(b[7]), .C1(n1585), .C2(b[6]), .A(n1867), 
        .ZN(n1866) );
  OAI22_X1 U1511 ( .A1(n1672), .A2(n1583), .B1(n1673), .B2(n1587), .ZN(n1867)
         );
  XNOR2_X1 U1512 ( .A(n1604), .B(n1868), .ZN(n818) );
  AOI221_X1 U1513 ( .B1(n1584), .B2(b[8]), .C1(n1585), .C2(b[7]), .A(n1869), 
        .ZN(n1868) );
  OAI22_X1 U1514 ( .A1(n1676), .A2(n1583), .B1(n1677), .B2(n1587), .ZN(n1869)
         );
  XNOR2_X1 U1515 ( .A(n1604), .B(n1870), .ZN(n817) );
  AOI221_X1 U1516 ( .B1(n1584), .B2(b[9]), .C1(n1585), .C2(b[8]), .A(n1871), 
        .ZN(n1870) );
  OAI22_X1 U1517 ( .A1(n1680), .A2(n1583), .B1(n1681), .B2(n1587), .ZN(n1871)
         );
  XNOR2_X1 U1518 ( .A(n1604), .B(n1872), .ZN(n816) );
  AOI221_X1 U1519 ( .B1(n1584), .B2(b[10]), .C1(n1585), .C2(b[9]), .A(n1873), 
        .ZN(n1872) );
  OAI22_X1 U1520 ( .A1(n1684), .A2(n1583), .B1(n1685), .B2(n1587), .ZN(n1873)
         );
  XNOR2_X1 U1521 ( .A(n1604), .B(n1874), .ZN(n815) );
  AOI221_X1 U1522 ( .B1(n1584), .B2(b[11]), .C1(n1585), .C2(b[10]), .A(n1875), 
        .ZN(n1874) );
  OAI22_X1 U1523 ( .A1(n1688), .A2(n1583), .B1(n1689), .B2(n1587), .ZN(n1875)
         );
  XNOR2_X1 U1524 ( .A(n1604), .B(n1876), .ZN(n814) );
  AOI221_X1 U1525 ( .B1(n1584), .B2(b[12]), .C1(n1585), .C2(b[11]), .A(n1877), 
        .ZN(n1876) );
  OAI22_X1 U1526 ( .A1(n1692), .A2(n1583), .B1(n1693), .B2(n1587), .ZN(n1877)
         );
  XNOR2_X1 U1527 ( .A(n1604), .B(n1878), .ZN(n813) );
  AOI221_X1 U1528 ( .B1(n1584), .B2(b[13]), .C1(n1585), .C2(b[12]), .A(n1879), 
        .ZN(n1878) );
  OAI22_X1 U1529 ( .A1(n1696), .A2(n1583), .B1(n1697), .B2(n1586), .ZN(n1879)
         );
  XNOR2_X1 U1530 ( .A(n1604), .B(n1880), .ZN(n812) );
  AOI221_X1 U1531 ( .B1(n1584), .B2(b[14]), .C1(n1585), .C2(b[13]), .A(n1881), 
        .ZN(n1880) );
  OAI22_X1 U1532 ( .A1(n1700), .A2(n1583), .B1(n1701), .B2(n1586), .ZN(n1881)
         );
  XNOR2_X1 U1533 ( .A(n1604), .B(n1882), .ZN(n811) );
  AOI221_X1 U1534 ( .B1(n1584), .B2(b[15]), .C1(n1585), .C2(b[14]), .A(n1883), 
        .ZN(n1882) );
  OAI22_X1 U1535 ( .A1(n1704), .A2(n1583), .B1(n1705), .B2(n1586), .ZN(n1883)
         );
  XNOR2_X1 U1536 ( .A(n1604), .B(n1884), .ZN(n810) );
  AOI221_X1 U1537 ( .B1(n1584), .B2(b[16]), .C1(n1585), .C2(b[15]), .A(n1885), 
        .ZN(n1884) );
  OAI22_X1 U1538 ( .A1(n1708), .A2(n1583), .B1(n1709), .B2(n1586), .ZN(n1885)
         );
  XNOR2_X1 U1539 ( .A(n1604), .B(n1886), .ZN(n809) );
  AOI221_X1 U1540 ( .B1(n1584), .B2(b[17]), .C1(n1585), .C2(b[16]), .A(n1887), 
        .ZN(n1886) );
  OAI22_X1 U1541 ( .A1(n1712), .A2(n1583), .B1(n1713), .B2(n1586), .ZN(n1887)
         );
  XNOR2_X1 U1542 ( .A(n1604), .B(n1888), .ZN(n808) );
  AOI221_X1 U1543 ( .B1(n1584), .B2(b[18]), .C1(n1585), .C2(b[17]), .A(n1889), 
        .ZN(n1888) );
  OAI22_X1 U1544 ( .A1(n1716), .A2(n1583), .B1(n1717), .B2(n1586), .ZN(n1889)
         );
  XNOR2_X1 U1545 ( .A(n1604), .B(n1890), .ZN(n807) );
  AOI221_X1 U1546 ( .B1(n1584), .B2(b[19]), .C1(n1585), .C2(b[18]), .A(n1891), 
        .ZN(n1890) );
  OAI22_X1 U1547 ( .A1(n1720), .A2(n1583), .B1(n1721), .B2(n1586), .ZN(n1891)
         );
  XNOR2_X1 U1548 ( .A(n1604), .B(n1892), .ZN(n806) );
  AOI221_X1 U1549 ( .B1(n1584), .B2(b[20]), .C1(n1585), .C2(b[19]), .A(n1893), 
        .ZN(n1892) );
  OAI22_X1 U1550 ( .A1(n1724), .A2(n1583), .B1(n1725), .B2(n1586), .ZN(n1893)
         );
  XNOR2_X1 U1551 ( .A(a[14]), .B(n1894), .ZN(n805) );
  AOI221_X1 U1552 ( .B1(n1584), .B2(b[21]), .C1(n1585), .C2(b[20]), .A(n1895), 
        .ZN(n1894) );
  OAI22_X1 U1553 ( .A1(n1728), .A2(n1583), .B1(n1729), .B2(n1586), .ZN(n1895)
         );
  XNOR2_X1 U1554 ( .A(a[14]), .B(n1896), .ZN(n804) );
  AOI221_X1 U1555 ( .B1(n1584), .B2(b[22]), .C1(n1553), .C2(n1376), .A(n1897), 
        .ZN(n1896) );
  OAI22_X1 U1556 ( .A1(n1640), .A2(n1587), .B1(n1643), .B2(n1550), .ZN(n1897)
         );
  XNOR2_X1 U1557 ( .A(a[14]), .B(n1898), .ZN(n803) );
  AOI221_X1 U1558 ( .B1(n1585), .B2(b[22]), .C1(n1553), .C2(n1375), .A(n1899), 
        .ZN(n1898) );
  OAI22_X1 U1559 ( .A1(n1617), .A2(n1541), .B1(n1643), .B2(n1586), .ZN(n1899)
         );
  XNOR2_X1 U1560 ( .A(a[14]), .B(n1900), .ZN(n802) );
  AOI221_X1 U1561 ( .B1(n1584), .B2(n1614), .C1(n1585), .C2(n1614), .A(n1901), 
        .ZN(n1900) );
  OAI22_X1 U1562 ( .A1(n1633), .A2(n1583), .B1(n1634), .B2(n1586), .ZN(n1901)
         );
  XNOR2_X1 U1563 ( .A(a[14]), .B(n1902), .ZN(n801) );
  OAI221_X1 U1564 ( .B1(n1617), .B2(n1587), .C1(n1619), .C2(n1583), .A(n1903), 
        .ZN(n1902) );
  OAI21_X1 U1565 ( .B1(n1584), .B2(n1585), .A(n1614), .ZN(n1903) );
  INV_X1 U1566 ( .A(n1907), .ZN(n1904) );
  NAND3_X1 U1567 ( .A1(n1907), .A2(n1906), .A3(n1905), .ZN(n1857) );
  XNOR2_X1 U1568 ( .A(a[12]), .B(a[13]), .ZN(n1905) );
  XNOR2_X1 U1569 ( .A(a[13]), .B(n1605), .ZN(n1906) );
  XOR2_X1 U1570 ( .A(a[12]), .B(n1607), .Z(n1907) );
  XNOR2_X1 U1571 ( .A(n1908), .B(n1603), .ZN(n800) );
  OAI22_X1 U1572 ( .A1(n1565), .A2(n1540), .B1(n1566), .B2(n1588), .ZN(n1908)
         );
  XNOR2_X1 U1573 ( .A(n1909), .B(n1603), .ZN(n799) );
  OAI222_X1 U1574 ( .A1(n1649), .A2(n1540), .B1(n1566), .B2(n1549), .C1(n1650), 
        .C2(n1588), .ZN(n1909) );
  XNOR2_X1 U1575 ( .A(n1602), .B(n1910), .ZN(n798) );
  AOI221_X1 U1576 ( .B1(n1589), .B2(b[2]), .C1(n1590), .C2(b[1]), .A(n1911), 
        .ZN(n1910) );
  OAI22_X1 U1577 ( .A1(n1653), .A2(n1588), .B1(n1566), .B2(n1591), .ZN(n1911)
         );
  XNOR2_X1 U1578 ( .A(n1602), .B(n1913), .ZN(n797) );
  AOI221_X1 U1579 ( .B1(n1589), .B2(b[3]), .C1(n1590), .C2(b[2]), .A(n1914), 
        .ZN(n1913) );
  OAI22_X1 U1580 ( .A1(n1657), .A2(n1588), .B1(n1649), .B2(n1592), .ZN(n1914)
         );
  XNOR2_X1 U1581 ( .A(n1602), .B(n1915), .ZN(n796) );
  AOI221_X1 U1582 ( .B1(n1589), .B2(b[4]), .C1(n1590), .C2(b[3]), .A(n1916), 
        .ZN(n1915) );
  OAI22_X1 U1583 ( .A1(n1660), .A2(n1588), .B1(n1661), .B2(n1592), .ZN(n1916)
         );
  XNOR2_X1 U1584 ( .A(n1602), .B(n1917), .ZN(n795) );
  AOI221_X1 U1585 ( .B1(n1589), .B2(b[5]), .C1(n1590), .C2(b[4]), .A(n1918), 
        .ZN(n1917) );
  OAI22_X1 U1586 ( .A1(n1664), .A2(n1588), .B1(n1665), .B2(n1592), .ZN(n1918)
         );
  XNOR2_X1 U1587 ( .A(n1602), .B(n1919), .ZN(n794) );
  AOI221_X1 U1588 ( .B1(n1589), .B2(b[6]), .C1(n1590), .C2(b[5]), .A(n1920), 
        .ZN(n1919) );
  OAI22_X1 U1589 ( .A1(n1668), .A2(n1588), .B1(n1669), .B2(n1592), .ZN(n1920)
         );
  XNOR2_X1 U1590 ( .A(n1602), .B(n1921), .ZN(n793) );
  AOI221_X1 U1591 ( .B1(n1589), .B2(b[7]), .C1(n1590), .C2(b[6]), .A(n1922), 
        .ZN(n1921) );
  OAI22_X1 U1592 ( .A1(n1672), .A2(n1588), .B1(n1673), .B2(n1592), .ZN(n1922)
         );
  XNOR2_X1 U1593 ( .A(n1602), .B(n1923), .ZN(n792) );
  AOI221_X1 U1594 ( .B1(n1589), .B2(b[8]), .C1(n1590), .C2(b[7]), .A(n1924), 
        .ZN(n1923) );
  OAI22_X1 U1595 ( .A1(n1676), .A2(n1588), .B1(n1677), .B2(n1592), .ZN(n1924)
         );
  XNOR2_X1 U1596 ( .A(n1602), .B(n1925), .ZN(n791) );
  AOI221_X1 U1597 ( .B1(n1589), .B2(b[9]), .C1(n1590), .C2(b[8]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1598 ( .A1(n1680), .A2(n1588), .B1(n1681), .B2(n1592), .ZN(n1926)
         );
  XNOR2_X1 U1599 ( .A(n1602), .B(n1927), .ZN(n790) );
  AOI221_X1 U1600 ( .B1(n1589), .B2(b[10]), .C1(n1590), .C2(b[9]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1601 ( .A1(n1684), .A2(n1588), .B1(n1685), .B2(n1592), .ZN(n1928)
         );
  XNOR2_X1 U1602 ( .A(n1602), .B(n1929), .ZN(n789) );
  AOI221_X1 U1603 ( .B1(n1589), .B2(b[11]), .C1(n1590), .C2(b[10]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1604 ( .A1(n1688), .A2(n1588), .B1(n1689), .B2(n1592), .ZN(n1930)
         );
  XNOR2_X1 U1605 ( .A(n1602), .B(n1931), .ZN(n788) );
  AOI221_X1 U1606 ( .B1(n1589), .B2(b[12]), .C1(n1590), .C2(b[11]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1607 ( .A1(n1692), .A2(n1588), .B1(n1693), .B2(n1592), .ZN(n1932)
         );
  XNOR2_X1 U1608 ( .A(n1602), .B(n1933), .ZN(n787) );
  AOI221_X1 U1609 ( .B1(n1589), .B2(b[13]), .C1(n1590), .C2(b[12]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1610 ( .A1(n1696), .A2(n1588), .B1(n1697), .B2(n1591), .ZN(n1934)
         );
  XNOR2_X1 U1611 ( .A(n1602), .B(n1935), .ZN(n786) );
  AOI221_X1 U1612 ( .B1(n1589), .B2(b[14]), .C1(n1590), .C2(b[13]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1613 ( .A1(n1700), .A2(n1588), .B1(n1701), .B2(n1591), .ZN(n1936)
         );
  XNOR2_X1 U1614 ( .A(n1602), .B(n1937), .ZN(n785) );
  AOI221_X1 U1615 ( .B1(n1589), .B2(b[15]), .C1(n1590), .C2(b[14]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1616 ( .A1(n1704), .A2(n1588), .B1(n1705), .B2(n1591), .ZN(n1938)
         );
  XNOR2_X1 U1617 ( .A(n1602), .B(n1939), .ZN(n784) );
  AOI221_X1 U1618 ( .B1(n1589), .B2(b[16]), .C1(n1590), .C2(b[15]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1619 ( .A1(n1708), .A2(n1588), .B1(n1709), .B2(n1591), .ZN(n1940)
         );
  XNOR2_X1 U1620 ( .A(n1602), .B(n1941), .ZN(n783) );
  AOI221_X1 U1621 ( .B1(n1589), .B2(b[17]), .C1(n1590), .C2(b[16]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1622 ( .A1(n1712), .A2(n1588), .B1(n1713), .B2(n1591), .ZN(n1942)
         );
  XNOR2_X1 U1623 ( .A(n1602), .B(n1943), .ZN(n782) );
  AOI221_X1 U1624 ( .B1(n1589), .B2(b[18]), .C1(n1590), .C2(b[17]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1625 ( .A1(n1716), .A2(n1588), .B1(n1717), .B2(n1591), .ZN(n1944)
         );
  XNOR2_X1 U1626 ( .A(n1602), .B(n1945), .ZN(n781) );
  AOI221_X1 U1627 ( .B1(n1589), .B2(b[19]), .C1(n1590), .C2(b[18]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1628 ( .A1(n1720), .A2(n1588), .B1(n1721), .B2(n1591), .ZN(n1946)
         );
  XNOR2_X1 U1629 ( .A(n1602), .B(n1947), .ZN(n780) );
  AOI221_X1 U1630 ( .B1(n1589), .B2(b[20]), .C1(n1590), .C2(b[19]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1631 ( .A1(n1724), .A2(n1588), .B1(n1725), .B2(n1591), .ZN(n1948)
         );
  XNOR2_X1 U1632 ( .A(a[17]), .B(n1949), .ZN(n779) );
  AOI221_X1 U1633 ( .B1(n1589), .B2(b[21]), .C1(n1590), .C2(b[20]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1634 ( .A1(n1728), .A2(n1588), .B1(n1729), .B2(n1591), .ZN(n1950)
         );
  XNOR2_X1 U1635 ( .A(a[17]), .B(n1951), .ZN(n778) );
  AOI221_X1 U1636 ( .B1(n1589), .B2(b[22]), .C1(n1552), .C2(n1376), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1637 ( .A1(n1640), .A2(n1592), .B1(n1643), .B2(n1549), .ZN(n1952)
         );
  XNOR2_X1 U1638 ( .A(a[17]), .B(n1953), .ZN(n777) );
  AOI221_X1 U1639 ( .B1(n1590), .B2(b[22]), .C1(n1552), .C2(n1375), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1640 ( .A1(n1617), .A2(n1540), .B1(n1643), .B2(n1591), .ZN(n1954)
         );
  XNOR2_X1 U1641 ( .A(a[17]), .B(n1955), .ZN(n776) );
  AOI221_X1 U1642 ( .B1(n1589), .B2(n1613), .C1(n1590), .C2(n1614), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1643 ( .A1(n1633), .A2(n1588), .B1(n1634), .B2(n1591), .ZN(n1956)
         );
  XNOR2_X1 U1644 ( .A(a[17]), .B(n1957), .ZN(n775) );
  OAI221_X1 U1645 ( .B1(n1618), .B2(n1592), .C1(n1617), .C2(n1588), .A(n1958), 
        .ZN(n1957) );
  OAI21_X1 U1646 ( .B1(n1589), .B2(n1590), .A(n1614), .ZN(n1958) );
  INV_X1 U1647 ( .A(n1962), .ZN(n1959) );
  NAND3_X1 U1648 ( .A1(n1962), .A2(n1961), .A3(n1960), .ZN(n1912) );
  XNOR2_X1 U1649 ( .A(a[15]), .B(a[16]), .ZN(n1960) );
  XNOR2_X1 U1650 ( .A(a[16]), .B(n1603), .ZN(n1961) );
  XOR2_X1 U1651 ( .A(a[15]), .B(n1605), .Z(n1962) );
  XOR2_X1 U1652 ( .A(n1963), .B(n1600), .Z(n774) );
  OAI22_X1 U1653 ( .A1(n1565), .A2(n1539), .B1(n1566), .B2(n1593), .ZN(n1963)
         );
  XOR2_X1 U1654 ( .A(n1964), .B(n1600), .Z(n773) );
  OAI222_X1 U1655 ( .A1(n1649), .A2(n1539), .B1(n1566), .B2(n1548), .C1(n1650), 
        .C2(n1593), .ZN(n1964) );
  XNOR2_X1 U1656 ( .A(n1600), .B(n1965), .ZN(n772) );
  AOI221_X1 U1657 ( .B1(n1594), .B2(b[2]), .C1(n1595), .C2(b[1]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1658 ( .A1(n1653), .A2(n1593), .B1(n1566), .B2(n1596), .ZN(n1966)
         );
  XNOR2_X1 U1659 ( .A(n1600), .B(n1968), .ZN(n771) );
  AOI221_X1 U1660 ( .B1(n1594), .B2(b[3]), .C1(n1595), .C2(b[2]), .A(n1969), 
        .ZN(n1968) );
  OAI22_X1 U1661 ( .A1(n1657), .A2(n1593), .B1(n1649), .B2(n1597), .ZN(n1969)
         );
  XNOR2_X1 U1662 ( .A(n1600), .B(n1970), .ZN(n770) );
  AOI221_X1 U1663 ( .B1(n1594), .B2(b[4]), .C1(n1595), .C2(b[3]), .A(n1971), 
        .ZN(n1970) );
  OAI22_X1 U1664 ( .A1(n1660), .A2(n1593), .B1(n1661), .B2(n1597), .ZN(n1971)
         );
  XNOR2_X1 U1665 ( .A(n1600), .B(n1972), .ZN(n769) );
  AOI221_X1 U1666 ( .B1(n1594), .B2(b[5]), .C1(n1595), .C2(b[4]), .A(n1973), 
        .ZN(n1972) );
  OAI22_X1 U1667 ( .A1(n1664), .A2(n1593), .B1(n1665), .B2(n1597), .ZN(n1973)
         );
  XNOR2_X1 U1668 ( .A(n1600), .B(n1974), .ZN(n768) );
  AOI221_X1 U1669 ( .B1(n1594), .B2(b[6]), .C1(n1595), .C2(b[5]), .A(n1975), 
        .ZN(n1974) );
  OAI22_X1 U1670 ( .A1(n1668), .A2(n1593), .B1(n1669), .B2(n1597), .ZN(n1975)
         );
  XNOR2_X1 U1671 ( .A(n1600), .B(n1976), .ZN(n767) );
  AOI221_X1 U1672 ( .B1(n1594), .B2(b[7]), .C1(n1595), .C2(b[6]), .A(n1977), 
        .ZN(n1976) );
  OAI22_X1 U1673 ( .A1(n1672), .A2(n1593), .B1(n1673), .B2(n1597), .ZN(n1977)
         );
  XNOR2_X1 U1674 ( .A(n1600), .B(n1978), .ZN(n766) );
  AOI221_X1 U1675 ( .B1(n1594), .B2(b[8]), .C1(n1595), .C2(b[7]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1676 ( .A1(n1676), .A2(n1593), .B1(n1677), .B2(n1597), .ZN(n1979)
         );
  XNOR2_X1 U1677 ( .A(n1600), .B(n1980), .ZN(n765) );
  AOI221_X1 U1678 ( .B1(n1594), .B2(b[9]), .C1(n1595), .C2(b[8]), .A(n1981), 
        .ZN(n1980) );
  OAI22_X1 U1679 ( .A1(n1680), .A2(n1593), .B1(n1681), .B2(n1597), .ZN(n1981)
         );
  XNOR2_X1 U1680 ( .A(n1600), .B(n1982), .ZN(n764) );
  AOI221_X1 U1681 ( .B1(n1594), .B2(b[10]), .C1(n1595), .C2(b[9]), .A(n1983), 
        .ZN(n1982) );
  OAI22_X1 U1682 ( .A1(n1684), .A2(n1593), .B1(n1685), .B2(n1597), .ZN(n1983)
         );
  XNOR2_X1 U1683 ( .A(n1600), .B(n1984), .ZN(n763) );
  AOI221_X1 U1684 ( .B1(n1594), .B2(b[11]), .C1(n1595), .C2(b[10]), .A(n1985), 
        .ZN(n1984) );
  OAI22_X1 U1685 ( .A1(n1688), .A2(n1593), .B1(n1689), .B2(n1597), .ZN(n1985)
         );
  XNOR2_X1 U1686 ( .A(n1601), .B(n1986), .ZN(n762) );
  AOI221_X1 U1687 ( .B1(n1594), .B2(b[12]), .C1(n1595), .C2(b[11]), .A(n1987), 
        .ZN(n1986) );
  OAI22_X1 U1688 ( .A1(n1692), .A2(n1593), .B1(n1693), .B2(n1597), .ZN(n1987)
         );
  XNOR2_X1 U1689 ( .A(n1601), .B(n1988), .ZN(n761) );
  AOI221_X1 U1690 ( .B1(n1594), .B2(b[13]), .C1(n1595), .C2(b[12]), .A(n1989), 
        .ZN(n1988) );
  OAI22_X1 U1691 ( .A1(n1696), .A2(n1593), .B1(n1697), .B2(n1596), .ZN(n1989)
         );
  XNOR2_X1 U1692 ( .A(n1601), .B(n1990), .ZN(n760) );
  AOI221_X1 U1693 ( .B1(n1594), .B2(b[14]), .C1(n1595), .C2(b[13]), .A(n1991), 
        .ZN(n1990) );
  OAI22_X1 U1694 ( .A1(n1700), .A2(n1593), .B1(n1701), .B2(n1596), .ZN(n1991)
         );
  XNOR2_X1 U1695 ( .A(n1601), .B(n1992), .ZN(n759) );
  AOI221_X1 U1696 ( .B1(n1594), .B2(b[15]), .C1(n1595), .C2(b[14]), .A(n1993), 
        .ZN(n1992) );
  OAI22_X1 U1697 ( .A1(n1704), .A2(n1593), .B1(n1705), .B2(n1596), .ZN(n1993)
         );
  XNOR2_X1 U1698 ( .A(n1601), .B(n1994), .ZN(n758) );
  AOI221_X1 U1699 ( .B1(n1594), .B2(b[16]), .C1(n1595), .C2(b[15]), .A(n1995), 
        .ZN(n1994) );
  OAI22_X1 U1700 ( .A1(n1708), .A2(n1593), .B1(n1709), .B2(n1596), .ZN(n1995)
         );
  XNOR2_X1 U1701 ( .A(n1601), .B(n1996), .ZN(n757) );
  AOI221_X1 U1702 ( .B1(n1594), .B2(b[17]), .C1(n1595), .C2(b[16]), .A(n1997), 
        .ZN(n1996) );
  OAI22_X1 U1703 ( .A1(n1712), .A2(n1593), .B1(n1713), .B2(n1596), .ZN(n1997)
         );
  XNOR2_X1 U1704 ( .A(n1601), .B(n1998), .ZN(n756) );
  AOI221_X1 U1705 ( .B1(n1594), .B2(b[18]), .C1(n1595), .C2(b[17]), .A(n1999), 
        .ZN(n1998) );
  OAI22_X1 U1706 ( .A1(n1716), .A2(n1593), .B1(n1717), .B2(n1596), .ZN(n1999)
         );
  XNOR2_X1 U1707 ( .A(n1601), .B(n2000), .ZN(n755) );
  AOI221_X1 U1708 ( .B1(n1594), .B2(b[19]), .C1(n1595), .C2(b[18]), .A(n2001), 
        .ZN(n2000) );
  OAI22_X1 U1709 ( .A1(n1720), .A2(n1593), .B1(n1721), .B2(n1596), .ZN(n2001)
         );
  XNOR2_X1 U1710 ( .A(n1601), .B(n2002), .ZN(n754) );
  AOI221_X1 U1711 ( .B1(n1594), .B2(b[20]), .C1(n1595), .C2(b[19]), .A(n2003), 
        .ZN(n2002) );
  OAI22_X1 U1712 ( .A1(n1724), .A2(n1593), .B1(n1725), .B2(n1596), .ZN(n2003)
         );
  XNOR2_X1 U1713 ( .A(n1601), .B(n2004), .ZN(n753) );
  AOI221_X1 U1714 ( .B1(n1594), .B2(b[21]), .C1(n1595), .C2(b[20]), .A(n2005), 
        .ZN(n2004) );
  OAI22_X1 U1715 ( .A1(n1728), .A2(n1593), .B1(n1729), .B2(n1596), .ZN(n2005)
         );
  XNOR2_X1 U1716 ( .A(n1601), .B(n2006), .ZN(n752) );
  AOI221_X1 U1717 ( .B1(n1594), .B2(b[22]), .C1(n1545), .C2(n1376), .A(n2007), 
        .ZN(n2006) );
  OAI22_X1 U1718 ( .A1(n1640), .A2(n1597), .B1(n1643), .B2(n1548), .ZN(n2007)
         );
  XNOR2_X1 U1719 ( .A(n1601), .B(n2008), .ZN(n751) );
  AOI221_X1 U1720 ( .B1(n1595), .B2(b[22]), .C1(n1545), .C2(n1375), .A(n2009), 
        .ZN(n2008) );
  OAI22_X1 U1721 ( .A1(n1617), .A2(n1539), .B1(n1643), .B2(n1596), .ZN(n2009)
         );
  XNOR2_X1 U1722 ( .A(n1601), .B(n2010), .ZN(n750) );
  AOI221_X1 U1723 ( .B1(n1594), .B2(n1612), .C1(n1595), .C2(n1614), .A(n2011), 
        .ZN(n2010) );
  OAI22_X1 U1724 ( .A1(n1633), .A2(n1593), .B1(n1634), .B2(n1596), .ZN(n2011)
         );
  INV_X1 U1725 ( .A(b[22]), .ZN(n1634) );
  INV_X1 U1726 ( .A(n1374), .ZN(n1633) );
  XNOR2_X1 U1727 ( .A(n1600), .B(n2012), .ZN(n749) );
  OAI221_X1 U1728 ( .B1(n1617), .B2(n1597), .C1(n1619), .C2(n1593), .A(n2013), 
        .ZN(n2012) );
  OAI21_X1 U1729 ( .B1(n1594), .B2(n1595), .A(n1614), .ZN(n2013) );
  INV_X1 U1730 ( .A(n2017), .ZN(n2014) );
  NAND3_X1 U1731 ( .A1(n2017), .A2(n2016), .A3(n2015), .ZN(n1967) );
  XNOR2_X1 U1732 ( .A(a[18]), .B(a[19]), .ZN(n2015) );
  XOR2_X1 U1733 ( .A(a[19]), .B(n1600), .Z(n2016) );
  XOR2_X1 U1734 ( .A(a[18]), .B(n1603), .Z(n2017) );
  XNOR2_X1 U1735 ( .A(n2018), .B(n1599), .ZN(n748) );
  OAI22_X1 U1736 ( .A1(n1538), .A2(n1567), .B1(n1558), .B2(n1567), .ZN(n2018)
         );
  XNOR2_X1 U1737 ( .A(n2019), .B(n1599), .ZN(n747) );
  OAI222_X1 U1738 ( .A1(n1538), .A2(n1649), .B1(n1547), .B2(n1566), .C1(n1558), 
        .C2(n1650), .ZN(n2019) );
  XNOR2_X1 U1739 ( .A(n1598), .B(n2020), .ZN(n746) );
  AOI221_X1 U1740 ( .B1(b[2]), .B2(n1559), .C1(b[1]), .C2(n1560), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1741 ( .A1(n1558), .A2(n1653), .B1(n1557), .B2(n1567), .ZN(n2021)
         );
  INV_X1 U1742 ( .A(b[0]), .ZN(n1647) );
  INV_X1 U1743 ( .A(n1396), .ZN(n1653) );
  XNOR2_X1 U1744 ( .A(n1598), .B(n2022), .ZN(n745) );
  AOI221_X1 U1745 ( .B1(b[3]), .B2(n1559), .C1(b[2]), .C2(n1560), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1746 ( .A1(n1558), .A2(n1657), .B1(n1557), .B2(n1649), .ZN(n2023)
         );
  XNOR2_X1 U1747 ( .A(n1598), .B(n2024), .ZN(n744) );
  AOI221_X1 U1748 ( .B1(b[4]), .B2(n1559), .C1(b[3]), .C2(n1560), .A(n2025), 
        .ZN(n2024) );
  OAI22_X1 U1749 ( .A1(n1558), .A2(n1660), .B1(n1557), .B2(n1661), .ZN(n2025)
         );
  XNOR2_X1 U1750 ( .A(n1598), .B(n2026), .ZN(n743) );
  AOI221_X1 U1751 ( .B1(b[5]), .B2(n1559), .C1(b[4]), .C2(n1560), .A(n2027), 
        .ZN(n2026) );
  OAI22_X1 U1752 ( .A1(n1558), .A2(n1664), .B1(n1557), .B2(n1665), .ZN(n2027)
         );
  XNOR2_X1 U1753 ( .A(n1598), .B(n2028), .ZN(n742) );
  AOI221_X1 U1754 ( .B1(b[6]), .B2(n1559), .C1(b[5]), .C2(n1560), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1755 ( .A1(n1558), .A2(n1668), .B1(n1557), .B2(n1669), .ZN(n2029)
         );
  XNOR2_X1 U1756 ( .A(n1598), .B(n2030), .ZN(n741) );
  AOI221_X1 U1757 ( .B1(b[7]), .B2(n1559), .C1(b[6]), .C2(n1560), .A(n2031), 
        .ZN(n2030) );
  OAI22_X1 U1758 ( .A1(n1558), .A2(n1672), .B1(n1557), .B2(n1673), .ZN(n2031)
         );
  XNOR2_X1 U1759 ( .A(n1598), .B(n2032), .ZN(n740) );
  AOI221_X1 U1760 ( .B1(b[9]), .B2(n1559), .C1(b[8]), .C2(n1560), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1761 ( .A1(n1558), .A2(n1680), .B1(n1557), .B2(n1681), .ZN(n2033)
         );
  XNOR2_X1 U1762 ( .A(n1598), .B(n2034), .ZN(n739) );
  AOI221_X1 U1763 ( .B1(b[10]), .B2(n1559), .C1(b[9]), .C2(n1560), .A(n2035), 
        .ZN(n2034) );
  OAI22_X1 U1764 ( .A1(n1558), .A2(n1684), .B1(n1557), .B2(n1685), .ZN(n2035)
         );
  XNOR2_X1 U1765 ( .A(n1598), .B(n2036), .ZN(n738) );
  AOI221_X1 U1766 ( .B1(b[12]), .B2(n1559), .C1(b[11]), .C2(n1560), .A(n2037), 
        .ZN(n2036) );
  OAI22_X1 U1767 ( .A1(n1558), .A2(n1692), .B1(n1557), .B2(n1693), .ZN(n2037)
         );
  XNOR2_X1 U1768 ( .A(n1598), .B(n2038), .ZN(n737) );
  AOI221_X1 U1769 ( .B1(b[13]), .B2(n1559), .C1(b[12]), .C2(n1560), .A(n2039), 
        .ZN(n2038) );
  OAI22_X1 U1770 ( .A1(n1558), .A2(n1696), .B1(n1557), .B2(n1697), .ZN(n2039)
         );
  XNOR2_X1 U1771 ( .A(n1598), .B(n2040), .ZN(n736) );
  AOI221_X1 U1772 ( .B1(b[14]), .B2(n1559), .C1(b[13]), .C2(n1560), .A(n2041), 
        .ZN(n2040) );
  OAI22_X1 U1773 ( .A1(n1558), .A2(n1700), .B1(n1556), .B2(n1701), .ZN(n2041)
         );
  XNOR2_X1 U1774 ( .A(n1598), .B(n2042), .ZN(n735) );
  AOI221_X1 U1775 ( .B1(b[15]), .B2(n1559), .C1(b[14]), .C2(n1560), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1776 ( .A1(n1558), .A2(n1704), .B1(n1556), .B2(n1705), .ZN(n2043)
         );
  XNOR2_X1 U1777 ( .A(n1598), .B(n2044), .ZN(n734) );
  AOI221_X1 U1778 ( .B1(b[16]), .B2(n1559), .C1(b[15]), .C2(n1560), .A(n2045), 
        .ZN(n2044) );
  OAI22_X1 U1779 ( .A1(n1558), .A2(n1708), .B1(n1556), .B2(n1709), .ZN(n2045)
         );
  XNOR2_X1 U1780 ( .A(n1598), .B(n2046), .ZN(n733) );
  AOI221_X1 U1781 ( .B1(b[18]), .B2(n1559), .C1(b[17]), .C2(n1560), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1782 ( .A1(n1558), .A2(n1716), .B1(n1556), .B2(n1717), .ZN(n2047)
         );
  XNOR2_X1 U1783 ( .A(n1598), .B(n2048), .ZN(n732) );
  AOI221_X1 U1784 ( .B1(b[19]), .B2(n1559), .C1(b[18]), .C2(n1560), .A(n2049), 
        .ZN(n2048) );
  OAI22_X1 U1785 ( .A1(n1558), .A2(n1720), .B1(n1556), .B2(n1721), .ZN(n2049)
         );
  XNOR2_X1 U1786 ( .A(n1598), .B(n2050), .ZN(n731) );
  AOI221_X1 U1787 ( .B1(b[20]), .B2(n1559), .C1(b[19]), .C2(n1560), .A(n2051), 
        .ZN(n2050) );
  OAI22_X1 U1788 ( .A1(n1558), .A2(n1724), .B1(n1556), .B2(n1725), .ZN(n2051)
         );
  XNOR2_X1 U1789 ( .A(a[23]), .B(n2052), .ZN(n730) );
  AOI221_X1 U1790 ( .B1(b[21]), .B2(n1559), .C1(b[20]), .C2(n1560), .A(n2053), 
        .ZN(n2052) );
  OAI22_X1 U1791 ( .A1(n1558), .A2(n1728), .B1(n1556), .B2(n1729), .ZN(n2053)
         );
  XNOR2_X1 U1792 ( .A(a[23]), .B(n2054), .ZN(n729) );
  AOI221_X1 U1793 ( .B1(b[22]), .B2(n1559), .C1(n1376), .C2(n1544), .A(n2055), 
        .ZN(n2054) );
  OAI22_X1 U1794 ( .A1(n1556), .A2(n1640), .B1(n1547), .B2(n1643), .ZN(n2055)
         );
  INV_X1 U1795 ( .A(b[20]), .ZN(n1640) );
  XNOR2_X1 U1796 ( .A(n519), .B(n2056), .ZN(n506) );
  INV_X1 U1797 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1798 ( .A1(n2056), .A2(n519), .ZN(n493) );
  XOR2_X1 U1799 ( .A(n2057), .B(n1742), .Z(n2056) );
  OAI221_X1 U1800 ( .B1(n1618), .B2(n1639), .C1(n1619), .C2(n1564), .A(n2058), 
        .ZN(n2057) );
  OAI21_X1 U1801 ( .B1(n1561), .B2(n1563), .A(n1614), .ZN(n2058) );
  INV_X1 U1802 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1803 ( .A(n1598), .B(n2059), .Z(n454) );
  AOI221_X1 U1804 ( .B1(b[8]), .B2(n1559), .C1(b[7]), .C2(n1560), .A(n2060), 
        .ZN(n2059) );
  OAI22_X1 U1805 ( .A1(n1558), .A2(n1676), .B1(n1556), .B2(n1677), .ZN(n2060)
         );
  INV_X1 U1806 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1807 ( .A(n1598), .B(n2061), .Z(n421) );
  AOI221_X1 U1808 ( .B1(b[11]), .B2(n1559), .C1(b[10]), .C2(n1560), .A(n2062), 
        .ZN(n2061) );
  OAI22_X1 U1809 ( .A1(n1558), .A2(n1688), .B1(n1556), .B2(n1689), .ZN(n2062)
         );
  INV_X1 U1810 ( .A(n387), .ZN(n395) );
  INV_X1 U1811 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1812 ( .A(n1598), .B(n2063), .Z(n374) );
  AOI221_X1 U1813 ( .B1(b[17]), .B2(n1559), .C1(b[16]), .C2(n1560), .A(n2064), 
        .ZN(n2063) );
  OAI22_X1 U1814 ( .A1(n1558), .A2(n1712), .B1(n1556), .B2(n1713), .ZN(n2064)
         );
  INV_X1 U1815 ( .A(n356), .ZN(n360) );
  INV_X1 U1816 ( .A(n1627), .ZN(n351) );
  XOR2_X1 U1817 ( .A(n1599), .B(n2065), .Z(n1627) );
  AOI221_X1 U1818 ( .B1(b[22]), .B2(n1560), .C1(n1375), .C2(n1544), .A(n2066), 
        .ZN(n2065) );
  OAI22_X1 U1819 ( .A1(n1538), .A2(n1618), .B1(n1556), .B2(n1643), .ZN(n2066)
         );
  INV_X1 U1820 ( .A(b[21]), .ZN(n1643) );
  NAND3_X1 U1821 ( .A1(n2067), .A2(n2068), .A3(n2069), .ZN(n1629) );
  XNOR2_X1 U1822 ( .A(a[22]), .B(n1599), .ZN(n2068) );
  XNOR2_X1 U1823 ( .A(a[21]), .B(a[22]), .ZN(n2069) );
  INV_X1 U1824 ( .A(n2067), .ZN(n2070) );
  XNOR2_X1 U1825 ( .A(a[21]), .B(n1600), .ZN(n2067) );
  OAI222_X1 U1826 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n2073), .C1(n2073), 
        .C2(n2072), .ZN(n326) );
  INV_X1 U1827 ( .A(n550), .ZN(n2073) );
  XNOR2_X1 U1828 ( .A(n1742), .B(n2074), .ZN(n2072) );
  AOI221_X1 U1829 ( .B1(n1561), .B2(b[21]), .C1(b[20]), .C2(n1562), .A(n2075), 
        .ZN(n2074) );
  OAI22_X1 U1830 ( .A1(n1564), .A2(n1728), .B1(n1639), .B2(n1729), .ZN(n2075)
         );
  INV_X1 U1831 ( .A(b[19]), .ZN(n1729) );
  INV_X1 U1832 ( .A(n1377), .ZN(n1728) );
  AOI222_X1 U1833 ( .A1(n2076), .A2(n2077), .B1(n2076), .B2(n564), .C1(n564), 
        .C2(n2077), .ZN(n2071) );
  XNOR2_X1 U1834 ( .A(a[2]), .B(n2078), .ZN(n2077) );
  AOI221_X1 U1835 ( .B1(b[20]), .B2(n1561), .C1(b[19]), .C2(n1562), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1836 ( .A1(n1564), .A2(n1724), .B1(n1639), .B2(n1725), .ZN(n2079)
         );
  INV_X1 U1837 ( .A(b[18]), .ZN(n1725) );
  INV_X1 U1838 ( .A(n1378), .ZN(n1724) );
  INV_X1 U1839 ( .A(n2080), .ZN(n2076) );
  AOI222_X1 U1840 ( .A1(n2081), .A2(n2082), .B1(n2081), .B2(n576), .C1(n576), 
        .C2(n2082), .ZN(n2080) );
  XNOR2_X1 U1841 ( .A(a[2]), .B(n2083), .ZN(n2082) );
  AOI221_X1 U1842 ( .B1(b[19]), .B2(n1561), .C1(b[18]), .C2(n1562), .A(n2084), 
        .ZN(n2083) );
  OAI22_X1 U1843 ( .A1(n1564), .A2(n1720), .B1(n1639), .B2(n1721), .ZN(n2084)
         );
  INV_X1 U1844 ( .A(b[17]), .ZN(n1721) );
  INV_X1 U1845 ( .A(n1379), .ZN(n1720) );
  OAI222_X1 U1846 ( .A1(n2085), .A2(n2086), .B1(n2085), .B2(n2087), .C1(n2087), 
        .C2(n2086), .ZN(n2081) );
  INV_X1 U1847 ( .A(n588), .ZN(n2087) );
  XNOR2_X1 U1848 ( .A(n1742), .B(n2088), .ZN(n2086) );
  AOI221_X1 U1849 ( .B1(b[18]), .B2(n1561), .C1(b[17]), .C2(n1562), .A(n2089), 
        .ZN(n2088) );
  OAI22_X1 U1850 ( .A1(n1564), .A2(n1716), .B1(n1639), .B2(n1717), .ZN(n2089)
         );
  INV_X1 U1851 ( .A(b[16]), .ZN(n1717) );
  INV_X1 U1852 ( .A(n1380), .ZN(n1716) );
  AOI222_X1 U1853 ( .A1(n2090), .A2(n2091), .B1(n2090), .B2(n600), .C1(n600), 
        .C2(n2091), .ZN(n2085) );
  XNOR2_X1 U1854 ( .A(a[2]), .B(n2092), .ZN(n2091) );
  AOI221_X1 U1855 ( .B1(b[17]), .B2(n1561), .C1(b[16]), .C2(n1562), .A(n2093), 
        .ZN(n2092) );
  OAI22_X1 U1856 ( .A1(n1564), .A2(n1712), .B1(n1639), .B2(n1713), .ZN(n2093)
         );
  INV_X1 U1857 ( .A(b[15]), .ZN(n1713) );
  INV_X1 U1858 ( .A(n1381), .ZN(n1712) );
  OAI222_X1 U1859 ( .A1(n2094), .A2(n2095), .B1(n2094), .B2(n2096), .C1(n2096), 
        .C2(n2095), .ZN(n2090) );
  INV_X1 U1860 ( .A(n610), .ZN(n2096) );
  XNOR2_X1 U1861 ( .A(n1742), .B(n2097), .ZN(n2095) );
  AOI221_X1 U1862 ( .B1(b[16]), .B2(n1561), .C1(b[15]), .C2(n1562), .A(n2098), 
        .ZN(n2097) );
  OAI22_X1 U1863 ( .A1(n1564), .A2(n1708), .B1(n1639), .B2(n1709), .ZN(n2098)
         );
  INV_X1 U1864 ( .A(b[14]), .ZN(n1709) );
  INV_X1 U1865 ( .A(n1382), .ZN(n1708) );
  AOI222_X1 U1866 ( .A1(n2099), .A2(n2100), .B1(n2099), .B2(n620), .C1(n620), 
        .C2(n2100), .ZN(n2094) );
  XNOR2_X1 U1867 ( .A(a[2]), .B(n2101), .ZN(n2100) );
  AOI221_X1 U1868 ( .B1(b[15]), .B2(n1561), .C1(b[14]), .C2(n1562), .A(n2102), 
        .ZN(n2101) );
  OAI22_X1 U1869 ( .A1(n1564), .A2(n1704), .B1(n1639), .B2(n1705), .ZN(n2102)
         );
  INV_X1 U1870 ( .A(b[13]), .ZN(n1705) );
  INV_X1 U1871 ( .A(n1383), .ZN(n1704) );
  OAI222_X1 U1872 ( .A1(n2103), .A2(n2104), .B1(n2103), .B2(n2105), .C1(n2105), 
        .C2(n2104), .ZN(n2099) );
  INV_X1 U1873 ( .A(n630), .ZN(n2105) );
  XNOR2_X1 U1874 ( .A(n1742), .B(n2106), .ZN(n2104) );
  AOI221_X1 U1875 ( .B1(b[14]), .B2(n1561), .C1(b[13]), .C2(n1562), .A(n2107), 
        .ZN(n2106) );
  OAI22_X1 U1876 ( .A1(n1564), .A2(n1700), .B1(n1639), .B2(n1701), .ZN(n2107)
         );
  INV_X1 U1877 ( .A(b[12]), .ZN(n1701) );
  INV_X1 U1878 ( .A(n1384), .ZN(n1700) );
  AOI222_X1 U1879 ( .A1(n2108), .A2(n2109), .B1(n2108), .B2(n638), .C1(n638), 
        .C2(n2109), .ZN(n2103) );
  XNOR2_X1 U1880 ( .A(a[2]), .B(n2110), .ZN(n2109) );
  AOI221_X1 U1881 ( .B1(b[13]), .B2(n1561), .C1(b[12]), .C2(n1562), .A(n2111), 
        .ZN(n2110) );
  OAI22_X1 U1882 ( .A1(n1564), .A2(n1696), .B1(n1639), .B2(n1697), .ZN(n2111)
         );
  INV_X1 U1883 ( .A(b[11]), .ZN(n1697) );
  INV_X1 U1884 ( .A(n1385), .ZN(n1696) );
  OAI222_X1 U1885 ( .A1(n2112), .A2(n2113), .B1(n2112), .B2(n2114), .C1(n2114), 
        .C2(n2113), .ZN(n2108) );
  INV_X1 U1886 ( .A(n646), .ZN(n2114) );
  XNOR2_X1 U1887 ( .A(n1742), .B(n2115), .ZN(n2113) );
  AOI221_X1 U1888 ( .B1(b[12]), .B2(n1561), .C1(b[11]), .C2(n1562), .A(n2116), 
        .ZN(n2115) );
  OAI22_X1 U1889 ( .A1(n1564), .A2(n1692), .B1(n1639), .B2(n1693), .ZN(n2116)
         );
  INV_X1 U1890 ( .A(b[10]), .ZN(n1693) );
  INV_X1 U1891 ( .A(n1386), .ZN(n1692) );
  AOI222_X1 U1892 ( .A1(n2117), .A2(n2118), .B1(n2117), .B2(n654), .C1(n654), 
        .C2(n2118), .ZN(n2112) );
  XNOR2_X1 U1893 ( .A(a[2]), .B(n2119), .ZN(n2118) );
  AOI221_X1 U1894 ( .B1(b[11]), .B2(n1561), .C1(b[10]), .C2(n1562), .A(n2120), 
        .ZN(n2119) );
  OAI22_X1 U1895 ( .A1(n1564), .A2(n1688), .B1(n1639), .B2(n1689), .ZN(n2120)
         );
  INV_X1 U1896 ( .A(b[9]), .ZN(n1689) );
  INV_X1 U1897 ( .A(n1387), .ZN(n1688) );
  OAI222_X1 U1898 ( .A1(n2121), .A2(n2122), .B1(n2121), .B2(n2123), .C1(n2123), 
        .C2(n2122), .ZN(n2117) );
  INV_X1 U1899 ( .A(n660), .ZN(n2123) );
  XNOR2_X1 U1900 ( .A(n1742), .B(n2124), .ZN(n2122) );
  AOI221_X1 U1901 ( .B1(b[10]), .B2(n1561), .C1(b[9]), .C2(n1563), .A(n2125), 
        .ZN(n2124) );
  OAI22_X1 U1902 ( .A1(n1564), .A2(n1684), .B1(n1639), .B2(n1685), .ZN(n2125)
         );
  INV_X1 U1903 ( .A(b[8]), .ZN(n1685) );
  INV_X1 U1904 ( .A(n1388), .ZN(n1684) );
  AOI222_X1 U1905 ( .A1(n2126), .A2(n2127), .B1(n2126), .B2(n666), .C1(n666), 
        .C2(n2127), .ZN(n2121) );
  XNOR2_X1 U1906 ( .A(a[2]), .B(n2128), .ZN(n2127) );
  AOI221_X1 U1907 ( .B1(b[9]), .B2(n1561), .C1(b[8]), .C2(n1563), .A(n2129), 
        .ZN(n2128) );
  OAI22_X1 U1908 ( .A1(n1564), .A2(n1680), .B1(n1639), .B2(n1681), .ZN(n2129)
         );
  INV_X1 U1909 ( .A(b[7]), .ZN(n1681) );
  INV_X1 U1910 ( .A(n1389), .ZN(n1680) );
  OAI222_X1 U1911 ( .A1(n2130), .A2(n2131), .B1(n2130), .B2(n2132), .C1(n2132), 
        .C2(n2131), .ZN(n2126) );
  INV_X1 U1912 ( .A(n672), .ZN(n2132) );
  XNOR2_X1 U1913 ( .A(n1742), .B(n2133), .ZN(n2131) );
  AOI221_X1 U1914 ( .B1(b[8]), .B2(n1561), .C1(b[7]), .C2(n1562), .A(n2134), 
        .ZN(n2133) );
  OAI22_X1 U1915 ( .A1(n1564), .A2(n1676), .B1(n1639), .B2(n1677), .ZN(n2134)
         );
  INV_X1 U1916 ( .A(b[6]), .ZN(n1677) );
  INV_X1 U1917 ( .A(n1390), .ZN(n1676) );
  AOI222_X1 U1918 ( .A1(n2135), .A2(n2136), .B1(n2135), .B2(n676), .C1(n676), 
        .C2(n2136), .ZN(n2130) );
  XNOR2_X1 U1919 ( .A(a[2]), .B(n2137), .ZN(n2136) );
  AOI221_X1 U1920 ( .B1(b[7]), .B2(n1561), .C1(b[6]), .C2(n1563), .A(n2138), 
        .ZN(n2137) );
  OAI22_X1 U1921 ( .A1(n1564), .A2(n1672), .B1(n1639), .B2(n1673), .ZN(n2138)
         );
  INV_X1 U1922 ( .A(b[5]), .ZN(n1673) );
  INV_X1 U1923 ( .A(n1391), .ZN(n1672) );
  OAI222_X1 U1924 ( .A1(n2139), .A2(n2140), .B1(n2139), .B2(n2141), .C1(n2141), 
        .C2(n2140), .ZN(n2135) );
  INV_X1 U1925 ( .A(n680), .ZN(n2141) );
  XNOR2_X1 U1926 ( .A(n1742), .B(n2142), .ZN(n2140) );
  AOI221_X1 U1927 ( .B1(b[6]), .B2(n1561), .C1(b[5]), .C2(n1563), .A(n2143), 
        .ZN(n2142) );
  OAI22_X1 U1928 ( .A1(n1564), .A2(n1668), .B1(n1639), .B2(n1669), .ZN(n2143)
         );
  INV_X1 U1929 ( .A(b[4]), .ZN(n1669) );
  INV_X1 U1930 ( .A(n1392), .ZN(n1668) );
  AOI222_X1 U1931 ( .A1(n2144), .A2(n2145), .B1(n2144), .B2(n684), .C1(n684), 
        .C2(n2145), .ZN(n2139) );
  XNOR2_X1 U1932 ( .A(a[2]), .B(n2146), .ZN(n2145) );
  AOI221_X1 U1933 ( .B1(b[5]), .B2(n1561), .C1(b[4]), .C2(n1563), .A(n2147), 
        .ZN(n2146) );
  OAI22_X1 U1934 ( .A1(n1564), .A2(n1664), .B1(n1639), .B2(n1665), .ZN(n2147)
         );
  INV_X1 U1935 ( .A(b[3]), .ZN(n1665) );
  INV_X1 U1936 ( .A(n1393), .ZN(n1664) );
  OAI222_X1 U1937 ( .A1(n2148), .A2(n2149), .B1(n2148), .B2(n2150), .C1(n2150), 
        .C2(n2149), .ZN(n2144) );
  INV_X1 U1938 ( .A(n686), .ZN(n2150) );
  XNOR2_X1 U1939 ( .A(n1742), .B(n2151), .ZN(n2149) );
  AOI221_X1 U1940 ( .B1(b[4]), .B2(n1561), .C1(b[3]), .C2(n1563), .A(n2152), 
        .ZN(n2151) );
  OAI22_X1 U1941 ( .A1(n1564), .A2(n1660), .B1(n1639), .B2(n1661), .ZN(n2152)
         );
  INV_X1 U1942 ( .A(n1394), .ZN(n1660) );
  AOI222_X1 U1943 ( .A1(n2153), .A2(n2154), .B1(n2153), .B2(n688), .C1(n688), 
        .C2(n2154), .ZN(n2148) );
  XNOR2_X1 U1944 ( .A(a[2]), .B(n2155), .ZN(n2154) );
  AOI221_X1 U1945 ( .B1(b[3]), .B2(n1561), .C1(b[2]), .C2(n1563), .A(n2156), 
        .ZN(n2155) );
  OAI22_X1 U1946 ( .A1(n1564), .A2(n1657), .B1(n1639), .B2(n1649), .ZN(n2156)
         );
  INV_X1 U1947 ( .A(b[1]), .ZN(n1649) );
  INV_X1 U1948 ( .A(n1395), .ZN(n1657) );
  AND2_X1 U1949 ( .A1(n2160), .A2(n2161), .ZN(n2153) );
  AOI211_X1 U1950 ( .C1(b[1]), .C2(n1561), .A(n2162), .B(b[0]), .ZN(n2161) );
  OAI22_X1 U1951 ( .A1(n1535), .A2(n1661), .B1(n1564), .B2(n1650), .ZN(n2162)
         );
  INV_X1 U1952 ( .A(n1397), .ZN(n1650) );
  INV_X1 U1953 ( .A(b[2]), .ZN(n1661) );
  INV_X1 U1954 ( .A(a[0]), .ZN(n2158) );
  AOI221_X1 U1955 ( .B1(b[1]), .B2(n1563), .C1(n1396), .C2(n1555), .A(n1742), 
        .ZN(n2160) );
  XNOR2_X1 U1956 ( .A(a[1]), .B(n1742), .ZN(n2157) );
  INV_X1 U1957 ( .A(a[2]), .ZN(n1742) );
  NOR2_X1 U1958 ( .A1(n2159), .A2(a[0]), .ZN(n1636) );
  INV_X1 U1959 ( .A(a[1]), .ZN(n2159) );
endmodule


module iir_filter_DW01_add_2 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_add_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  OAI21_X1 U1 ( .B1(n1), .B2(n2), .A(n3), .ZN(carry_11_) );
  OAI21_X1 U2 ( .B1(A[10]), .B2(n4), .A(B[10]), .ZN(n3) );
  INV_X1 U3 ( .A(n1), .ZN(n4) );
  INV_X1 U4 ( .A(A[10]), .ZN(n2) );
  AOI21_X1 U5 ( .B1(n5), .B2(A[9]), .A(n6), .ZN(n1) );
  INV_X1 U6 ( .A(n7), .ZN(n6) );
  OAI21_X1 U7 ( .B1(A[9]), .B2(n5), .A(B[9]), .ZN(n7) );
  OAI21_X1 U8 ( .B1(n8), .B2(n9), .A(n10), .ZN(n5) );
  OAI21_X1 U9 ( .B1(A[8]), .B2(n11), .A(B[8]), .ZN(n10) );
  INV_X1 U10 ( .A(n8), .ZN(n11) );
  INV_X1 U11 ( .A(A[8]), .ZN(n9) );
  AOI21_X1 U12 ( .B1(n12), .B2(A[7]), .A(n13), .ZN(n8) );
  INV_X1 U13 ( .A(n14), .ZN(n13) );
  OAI21_X1 U14 ( .B1(A[7]), .B2(n12), .A(B[7]), .ZN(n14) );
  OAI21_X1 U15 ( .B1(n15), .B2(n16), .A(n17), .ZN(n12) );
  OAI21_X1 U16 ( .B1(A[6]), .B2(n18), .A(B[6]), .ZN(n17) );
  INV_X1 U17 ( .A(A[6]), .ZN(n16) );
  INV_X1 U18 ( .A(n18), .ZN(n15) );
  OAI21_X1 U19 ( .B1(n19), .B2(n20), .A(n21), .ZN(n18) );
  OAI21_X1 U20 ( .B1(A[5]), .B2(n22), .A(B[5]), .ZN(n21) );
  INV_X1 U21 ( .A(A[5]), .ZN(n20) );
  INV_X1 U22 ( .A(n22), .ZN(n19) );
  OAI21_X1 U23 ( .B1(n23), .B2(n24), .A(n25), .ZN(n22) );
  OAI21_X1 U24 ( .B1(A[4]), .B2(n26), .A(B[4]), .ZN(n25) );
  INV_X1 U25 ( .A(A[4]), .ZN(n24) );
  INV_X1 U26 ( .A(n26), .ZN(n23) );
  OAI21_X1 U27 ( .B1(n27), .B2(n28), .A(n29), .ZN(n26) );
  OAI21_X1 U28 ( .B1(A[3]), .B2(n30), .A(B[3]), .ZN(n29) );
  INV_X1 U29 ( .A(A[3]), .ZN(n28) );
  INV_X1 U30 ( .A(n30), .ZN(n27) );
  OAI21_X1 U31 ( .B1(n31), .B2(n32), .A(n33), .ZN(n30) );
  OAI21_X1 U32 ( .B1(A[2]), .B2(n34), .A(B[2]), .ZN(n33) );
  INV_X1 U33 ( .A(A[2]), .ZN(n32) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  OAI21_X1 U35 ( .B1(n35), .B2(n36), .A(n37), .ZN(n34) );
  OAI211_X1 U36 ( .C1(A[1]), .C2(B[1]), .A(A[0]), .B(B[0]), .ZN(n37) );
  INV_X1 U37 ( .A(B[1]), .ZN(n36) );
  INV_X1 U38 ( .A(A[1]), .ZN(n35) );
endmodule


module iir_filter ( clk, rst_n, vIn, dIn, coeffs_fb, coeffs_ff, dOut, vOut );
  input [11:0] dIn;
  input [47:0] coeffs_fb;
  input [95:0] coeffs_ff;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   delayed_controls_0__1_, delayed_controls_1__0_,
         delayed_controls_1__1_, delayed_controls_2__0_, DP_N4, DP_N2, DP_y_0_,
         DP_y_1_, DP_y_2_, DP_y_3_, DP_y_4_, DP_y_5_, DP_y_6_, DP_y_7_,
         DP_y_8_, DP_y_9_, DP_y_10_, DP_y_11_, DP_y_23, DP_sw1_0_, DP_sw1_1_,
         DP_sw1_2_, DP_sw1_3_, DP_sw1_4_, DP_sw1_5_, DP_sw1_6_, DP_sw1_7_,
         DP_sw1_8_, DP_sw1_9_, DP_sw1_10_, DP_sw1_11_, DP_sw1_12_, DP_sw1_13_,
         DP_sw1_14_, DP_sw1_15_, DP_sw1_16_, DP_sw1_17_, DP_sw1_18_,
         DP_sw1_19_, DP_sw1_20_, DP_sw1_21_, DP_sw1_22_, DP_sw0_0_, DP_sw0_1_,
         DP_sw0_2_, DP_sw0_3_, DP_sw0_4_, DP_sw0_5_, DP_sw0_6_, DP_sw0_7_,
         DP_sw0_8_, DP_sw0_9_, DP_sw0_10_, DP_sw0_11_, DP_sw0_12_, DP_sw0_13_,
         DP_sw0_14_, DP_sw0_15_, DP_sw0_16_, DP_sw0_17_, DP_sw0_18_,
         DP_sw0_19_, DP_sw0_20_, DP_sw0_21_, DP_sw0_22_, DP_sw0_23_, DP_w_0_,
         DP_w_1_, DP_w_2_, DP_w_3_, DP_w_4_, DP_w_5_, DP_w_6_, DP_w_7_,
         DP_w_8_, DP_w_9_, DP_w_10_, DP_w_11_, DP_w_12_, DP_w_13_, DP_w_14_,
         DP_w_15_, DP_w_16_, DP_w_17_, DP_w_18_, DP_w_19_, DP_w_20_, DP_w_21_,
         DP_w_22_, DP_w_23_, CU_nextState_0_, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n38, n39, n40, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n529, n531, n533, n535, n537, n539, n541, n543, n545, n547, n549,
         n551, n553, n555, n557, n559, n561, n563, n565, n567, n569, n571,
         n573, n575, n577, n579, n581, n583, n585, n587, n589, n591, n593,
         n595, n597, n599, n601, n603, n605, n607, n609, n611, n613, n615,
         n617, n619, n621, n623, n625, n627, n629, n631, n633, n635, n637,
         n639, n641, n643, n645, n647, n649, n651, n653, n655, n657, n659,
         n661, n663, n665, n667, n669, n671, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, DP_fb_9_, DP_fb_8_,
         DP_fb_7_, DP_fb_6_, DP_fb_5_, DP_fb_4_, DP_fb_3_, DP_fb_2_, DP_fb_23_,
         DP_fb_22_, DP_fb_21_, DP_fb_20_, DP_fb_1_, DP_fb_19_, DP_fb_18_,
         DP_fb_17_, DP_fb_16_, DP_fb_15_, DP_fb_14_, DP_fb_13_, DP_fb_12_,
         DP_fb_11_, DP_fb_10_, DP_fb_0_, DP_ff_part_9_, DP_ff_part_8_,
         DP_ff_part_7_, DP_ff_part_6_, DP_ff_part_5_, DP_ff_part_4_,
         DP_ff_part_3_, DP_ff_part_2_, DP_ff_part_23_, DP_ff_part_22_,
         DP_ff_part_21_, DP_ff_part_20_, DP_ff_part_1_, DP_ff_part_19_,
         DP_ff_part_18_, DP_ff_part_17_, DP_ff_part_16_, DP_ff_part_15_,
         DP_ff_part_14_, DP_ff_part_13_, DP_ff_part_12_, DP_ff_part_11_,
         DP_ff_part_10_, DP_ff_part_0_, DP_ff_9_, DP_ff_8_, DP_ff_7_, DP_ff_6_,
         DP_ff_5_, DP_ff_4_, DP_ff_3_, DP_ff_2_, DP_ff_23_, DP_ff_22_,
         DP_ff_21_, DP_ff_20_, DP_ff_1_, DP_ff_19_, DP_ff_18_, DP_ff_17_,
         DP_ff_16_, DP_ff_15_, DP_ff_14_, DP_ff_13_, DP_ff_12_, DP_ff_11_,
         DP_ff_10_, DP_ff_0_, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175;
  wire   [0:23] DP_pipe13;
  wire   [0:23] DP_pipe0_coeff_pipe03;
  wire   [0:23] DP_pipe12;
  wire   [0:23] DP_pipe0_coeff_pipe02;
  wire   [0:23] DP_pipe11;
  wire   [0:23] DP_pipe0_coeff_pipe01;
  wire   [0:23] DP_pipe10;
  wire   [0:23] DP_pipe0_coeff_pipe00;
  wire   [0:23] DP_pipe03;
  wire   [0:23] DP_pipe02;
  wire   [0:23] DP_pipe01;
  wire   [0:23] DP_pipe00;
  wire   [0:23] DP_ret1;
  wire   [0:23] DP_sw1_coeff_ret1;
  wire   [0:23] DP_ret0;
  wire   [0:23] DP_sw0_coeff_ret0;
  wire   [0:23] DP_sw2;
  wire   [95:0] DP_coeffs_ff_int;
  wire   [47:0] DP_coeffs_fb_int;
  wire   [0:11] DP_x;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154;

  DFFR_X1 DP_reg_in_Q_reg_0_ ( .D(n995), .CK(clk), .RN(n1122), .Q(DP_x[0]) );
  DFFR_X1 DP_reg_in_Q_reg_1_ ( .D(n994), .CK(clk), .RN(n1122), .Q(DP_x[1]) );
  DFFR_X1 DP_reg_in_Q_reg_2_ ( .D(n993), .CK(clk), .RN(n1122), .Q(DP_x[2]) );
  DFFR_X1 DP_reg_in_Q_reg_3_ ( .D(n992), .CK(clk), .RN(n1122), .Q(DP_x[3]) );
  DFFR_X1 DP_reg_in_Q_reg_4_ ( .D(n991), .CK(clk), .RN(n1122), .Q(DP_x[4]) );
  DFFR_X1 DP_reg_in_Q_reg_5_ ( .D(n990), .CK(clk), .RN(n1122), .Q(DP_x[5]) );
  DFFR_X1 DP_reg_in_Q_reg_6_ ( .D(n989), .CK(clk), .RN(n1122), .Q(DP_x[6]) );
  DFFR_X1 DP_reg_in_Q_reg_7_ ( .D(n988), .CK(clk), .RN(n1122), .Q(DP_x[7]) );
  DFFR_X1 DP_reg_in_Q_reg_8_ ( .D(n987), .CK(clk), .RN(n1122), .Q(DP_x[8]) );
  DFFR_X1 DP_reg_in_Q_reg_9_ ( .D(n986), .CK(clk), .RN(n1122), .Q(DP_x[9]) );
  DFFR_X1 DP_reg_in_Q_reg_10_ ( .D(n985), .CK(clk), .RN(n1122), .Q(DP_x[10])
         );
  DFFR_X1 DP_reg_in_Q_reg_11_ ( .D(n984), .CK(clk), .RN(n1122), .Q(DP_x[11])
         );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_0_ ( .D(n983), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[23]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_1_ ( .D(n982), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[22]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_2_ ( .D(n981), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[21]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_3_ ( .D(n980), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[20]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_4_ ( .D(n979), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[19]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_5_ ( .D(n978), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[18]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_6_ ( .D(n977), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[17]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_7_ ( .D(n976), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[16]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_8_ ( .D(n975), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[15]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_9_ ( .D(n974), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[14]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_10_ ( .D(n973), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[13]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_11_ ( .D(n972), .CK(clk), .RN(n1123), .Q(
        DP_coeffs_fb_int[12]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_12_ ( .D(n971), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[11]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_13_ ( .D(n970), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[10]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_14_ ( .D(n969), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[9]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_15_ ( .D(n968), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[8]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_16_ ( .D(n967), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[7]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_17_ ( .D(n966), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[6]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_18_ ( .D(n965), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[5]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_19_ ( .D(n964), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[4]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_20_ ( .D(n963), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[3]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_21_ ( .D(n962), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[2]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_22_ ( .D(n961), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[1]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_23_ ( .D(n960), .CK(clk), .RN(n1124), .Q(
        DP_coeffs_fb_int[0]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_0_ ( .D(n959), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[47]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_1_ ( .D(n958), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[46]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_2_ ( .D(n957), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[45]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_3_ ( .D(n956), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[44]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_4_ ( .D(n955), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[43]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_5_ ( .D(n954), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[42]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_6_ ( .D(n953), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[41]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_7_ ( .D(n952), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[40]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_8_ ( .D(n951), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[39]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_9_ ( .D(n950), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[38]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_10_ ( .D(n949), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[37]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_11_ ( .D(n948), .CK(clk), .RN(n1125), .Q(
        DP_coeffs_fb_int[36]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_12_ ( .D(n947), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[35]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_13_ ( .D(n946), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[34]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_14_ ( .D(n945), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[33]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_15_ ( .D(n944), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[32]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_16_ ( .D(n943), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[31]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_17_ ( .D(n942), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[30]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_18_ ( .D(n941), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[29]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_19_ ( .D(n940), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[28]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_20_ ( .D(n939), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[27]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_21_ ( .D(n938), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[26]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_22_ ( .D(n937), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[25]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_23_ ( .D(n936), .CK(clk), .RN(n1126), .Q(
        DP_coeffs_fb_int[24]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_0_ ( .D(n935), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[23]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_1_ ( .D(n934), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[22]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_2_ ( .D(n933), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[21]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_3_ ( .D(n932), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[20]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_4_ ( .D(n931), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[19]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_5_ ( .D(n930), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[18]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_6_ ( .D(n929), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[17]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_7_ ( .D(n928), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[16]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_8_ ( .D(n927), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[15]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_9_ ( .D(n926), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[14]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_10_ ( .D(n925), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[13]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_11_ ( .D(n924), .CK(clk), .RN(n1127), .Q(
        DP_coeffs_ff_int[12]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_12_ ( .D(n923), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[11]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_13_ ( .D(n922), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[10]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_14_ ( .D(n921), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[9]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_15_ ( .D(n920), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[8]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_16_ ( .D(n919), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[7]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_17_ ( .D(n918), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[6]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_18_ ( .D(n917), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[5]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_19_ ( .D(n916), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[4]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_20_ ( .D(n915), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[3]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_21_ ( .D(n914), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[2]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_22_ ( .D(n913), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[1]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_23_ ( .D(n912), .CK(clk), .RN(n1128), .Q(
        DP_coeffs_ff_int[0]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_0_ ( .D(n911), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[47]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_1_ ( .D(n910), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[46]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_2_ ( .D(n909), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[45]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_3_ ( .D(n908), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[44]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_4_ ( .D(n907), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[43]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_5_ ( .D(n906), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[42]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_6_ ( .D(n905), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[41]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_7_ ( .D(n904), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[40]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_8_ ( .D(n903), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[39]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_9_ ( .D(n902), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[38]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_10_ ( .D(n901), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[37]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_11_ ( .D(n900), .CK(clk), .RN(n1129), .Q(
        DP_coeffs_ff_int[36]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_12_ ( .D(n899), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[35]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_13_ ( .D(n898), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[34]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_14_ ( .D(n897), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[33]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_15_ ( .D(n896), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[32]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_16_ ( .D(n895), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[31]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_17_ ( .D(n894), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[30]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_18_ ( .D(n893), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[29]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_19_ ( .D(n892), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[28]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_20_ ( .D(n891), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[27]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_21_ ( .D(n890), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[26]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_22_ ( .D(n889), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[25]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_23_ ( .D(n888), .CK(clk), .RN(n1130), .Q(
        DP_coeffs_ff_int[24]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_0_ ( .D(n887), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[71]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_1_ ( .D(n886), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[70]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_2_ ( .D(n885), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[69]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_3_ ( .D(n884), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[68]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_4_ ( .D(n883), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[67]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_5_ ( .D(n882), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[66]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_6_ ( .D(n881), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[65]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_7_ ( .D(n880), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[64]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_8_ ( .D(n879), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[63]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_9_ ( .D(n878), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[62]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_10_ ( .D(n877), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[61]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_11_ ( .D(n876), .CK(clk), .RN(n1131), .Q(
        DP_coeffs_ff_int[60]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_12_ ( .D(n875), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[59]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_13_ ( .D(n874), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[58]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_14_ ( .D(n873), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[57]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_15_ ( .D(n872), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[56]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_16_ ( .D(n871), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[55]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_17_ ( .D(n870), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[54]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_18_ ( .D(n869), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[53]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_19_ ( .D(n868), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[52]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_20_ ( .D(n867), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[51]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_21_ ( .D(n866), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[50]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_22_ ( .D(n865), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[49]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_23_ ( .D(n864), .CK(clk), .RN(n1132), .Q(
        DP_coeffs_ff_int[48]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_0_ ( .D(n863), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[95]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_1_ ( .D(n862), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[94]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_2_ ( .D(n861), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[93]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_3_ ( .D(n860), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[92]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_4_ ( .D(n859), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[91]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_5_ ( .D(n858), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[90]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_6_ ( .D(n857), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[89]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_7_ ( .D(n856), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[88]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_8_ ( .D(n855), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[87]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_9_ ( .D(n854), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[86]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_10_ ( .D(n853), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[85]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_11_ ( .D(n852), .CK(clk), .RN(n1133), .Q(
        DP_coeffs_ff_int[84]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_12_ ( .D(n851), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[83]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_13_ ( .D(n850), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[82]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_14_ ( .D(n849), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[81]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_15_ ( .D(n848), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[80]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_16_ ( .D(n847), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[79]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_17_ ( .D(n846), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[78]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_18_ ( .D(n845), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[77]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_19_ ( .D(n844), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[76]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_20_ ( .D(n843), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[75]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_21_ ( .D(n842), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[74]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_22_ ( .D(n841), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[73]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_23_ ( .D(n840), .CK(clk), .RN(n1134), .Q(
        DP_coeffs_ff_int[72]) );
  DFFR_X1 DP_reg_ret0_Q_reg_0_ ( .D(DP_sw0_coeff_ret0[0]), .CK(clk), .RN(n1135), .Q(DP_ret0[0]) );
  DFFR_X1 DP_reg_ret0_Q_reg_1_ ( .D(DP_sw0_coeff_ret0[1]), .CK(clk), .RN(n1135), .Q(DP_ret0[1]) );
  DFFR_X1 DP_reg_ret0_Q_reg_2_ ( .D(DP_sw0_coeff_ret0[2]), .CK(clk), .RN(n1135), .Q(DP_ret0[2]) );
  DFFR_X1 DP_reg_ret0_Q_reg_3_ ( .D(DP_sw0_coeff_ret0[3]), .CK(clk), .RN(n1135), .Q(DP_ret0[3]) );
  DFFR_X1 DP_reg_ret0_Q_reg_4_ ( .D(DP_sw0_coeff_ret0[4]), .CK(clk), .RN(n1135), .Q(DP_ret0[4]) );
  DFFR_X1 DP_reg_ret0_Q_reg_5_ ( .D(DP_sw0_coeff_ret0[5]), .CK(clk), .RN(n1135), .Q(DP_ret0[5]) );
  DFFR_X1 DP_reg_ret0_Q_reg_6_ ( .D(DP_sw0_coeff_ret0[6]), .CK(clk), .RN(n1135), .Q(DP_ret0[6]) );
  DFFR_X1 DP_reg_ret0_Q_reg_7_ ( .D(DP_sw0_coeff_ret0[7]), .CK(clk), .RN(n1135), .Q(DP_ret0[7]) );
  DFFR_X1 DP_reg_ret0_Q_reg_8_ ( .D(DP_sw0_coeff_ret0[8]), .CK(clk), .RN(n1135), .Q(DP_ret0[8]) );
  DFFR_X1 DP_reg_ret0_Q_reg_9_ ( .D(DP_sw0_coeff_ret0[9]), .CK(clk), .RN(n1135), .Q(DP_ret0[9]) );
  DFFR_X1 DP_reg_ret0_Q_reg_10_ ( .D(DP_sw0_coeff_ret0[10]), .CK(clk), .RN(
        n1135), .Q(DP_ret0[10]) );
  DFFR_X1 DP_reg_ret0_Q_reg_11_ ( .D(DP_sw0_coeff_ret0[11]), .CK(clk), .RN(
        n1135), .Q(DP_ret0[11]) );
  DFFR_X1 DP_reg_ret0_Q_reg_12_ ( .D(DP_sw0_coeff_ret0[12]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[12]) );
  DFFR_X1 DP_reg_ret0_Q_reg_13_ ( .D(DP_sw0_coeff_ret0[13]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[13]) );
  DFFR_X1 DP_reg_ret0_Q_reg_14_ ( .D(DP_sw0_coeff_ret0[14]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[14]) );
  DFFR_X1 DP_reg_ret0_Q_reg_15_ ( .D(DP_sw0_coeff_ret0[15]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[15]) );
  DFFR_X1 DP_reg_ret0_Q_reg_16_ ( .D(DP_sw0_coeff_ret0[16]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[16]) );
  DFFR_X1 DP_reg_ret0_Q_reg_17_ ( .D(DP_sw0_coeff_ret0[17]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[17]) );
  DFFR_X1 DP_reg_ret0_Q_reg_18_ ( .D(DP_sw0_coeff_ret0[18]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[18]) );
  DFFR_X1 DP_reg_ret0_Q_reg_19_ ( .D(DP_sw0_coeff_ret0[19]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[19]) );
  DFFR_X1 DP_reg_ret0_Q_reg_20_ ( .D(DP_sw0_coeff_ret0[20]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[20]) );
  DFFR_X1 DP_reg_ret0_Q_reg_21_ ( .D(DP_sw0_coeff_ret0[21]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[21]) );
  DFFR_X1 DP_reg_ret0_Q_reg_22_ ( .D(DP_sw0_coeff_ret0[22]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[22]) );
  DFFR_X1 DP_reg_ret0_Q_reg_23_ ( .D(DP_sw0_coeff_ret0[23]), .CK(clk), .RN(
        n1136), .Q(DP_ret0[23]) );
  DFFR_X1 DP_reg_ret1_Q_reg_0_ ( .D(DP_sw1_coeff_ret1[0]), .CK(clk), .RN(n1137), .Q(DP_ret1[0]) );
  DFFR_X1 DP_reg_ret1_Q_reg_1_ ( .D(DP_sw1_coeff_ret1[1]), .CK(clk), .RN(n1137), .Q(DP_ret1[1]) );
  DFFR_X1 DP_reg_ret1_Q_reg_2_ ( .D(DP_sw1_coeff_ret1[2]), .CK(clk), .RN(n1137), .Q(DP_ret1[2]) );
  DFFR_X1 DP_reg_ret1_Q_reg_3_ ( .D(DP_sw1_coeff_ret1[3]), .CK(clk), .RN(n1137), .Q(DP_ret1[3]) );
  DFFR_X1 DP_reg_ret1_Q_reg_4_ ( .D(DP_sw1_coeff_ret1[4]), .CK(clk), .RN(n1137), .Q(DP_ret1[4]) );
  DFFR_X1 DP_reg_ret1_Q_reg_5_ ( .D(DP_sw1_coeff_ret1[5]), .CK(clk), .RN(n1137), .Q(DP_ret1[5]) );
  DFFR_X1 DP_reg_ret1_Q_reg_6_ ( .D(DP_sw1_coeff_ret1[6]), .CK(clk), .RN(n1137), .Q(DP_ret1[6]) );
  DFFR_X1 DP_reg_ret1_Q_reg_7_ ( .D(DP_sw1_coeff_ret1[7]), .CK(clk), .RN(n1137), .Q(DP_ret1[7]) );
  DFFR_X1 DP_reg_ret1_Q_reg_8_ ( .D(DP_sw1_coeff_ret1[8]), .CK(clk), .RN(n1137), .Q(DP_ret1[8]) );
  DFFR_X1 DP_reg_ret1_Q_reg_9_ ( .D(DP_sw1_coeff_ret1[9]), .CK(clk), .RN(n1137), .Q(DP_ret1[9]) );
  DFFR_X1 DP_reg_ret1_Q_reg_10_ ( .D(DP_sw1_coeff_ret1[10]), .CK(clk), .RN(
        n1137), .Q(DP_ret1[10]) );
  DFFR_X1 DP_reg_ret1_Q_reg_11_ ( .D(DP_sw1_coeff_ret1[11]), .CK(clk), .RN(
        n1137), .Q(DP_ret1[11]) );
  DFFR_X1 DP_reg_ret1_Q_reg_12_ ( .D(DP_sw1_coeff_ret1[12]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[12]) );
  DFFR_X1 DP_reg_ret1_Q_reg_13_ ( .D(DP_sw1_coeff_ret1[13]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[13]) );
  DFFR_X1 DP_reg_ret1_Q_reg_14_ ( .D(DP_sw1_coeff_ret1[14]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[14]) );
  DFFR_X1 DP_reg_ret1_Q_reg_15_ ( .D(DP_sw1_coeff_ret1[15]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[15]) );
  DFFR_X1 DP_reg_ret1_Q_reg_16_ ( .D(DP_sw1_coeff_ret1[16]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[16]) );
  DFFR_X1 DP_reg_ret1_Q_reg_17_ ( .D(DP_sw1_coeff_ret1[17]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[17]) );
  DFFR_X1 DP_reg_ret1_Q_reg_18_ ( .D(DP_sw1_coeff_ret1[18]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[18]) );
  DFFR_X1 DP_reg_ret1_Q_reg_19_ ( .D(DP_sw1_coeff_ret1[19]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[19]) );
  DFFR_X1 DP_reg_ret1_Q_reg_20_ ( .D(DP_sw1_coeff_ret1[20]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[20]) );
  DFFR_X1 DP_reg_ret1_Q_reg_21_ ( .D(DP_sw1_coeff_ret1[21]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[21]) );
  DFFR_X1 DP_reg_ret1_Q_reg_22_ ( .D(DP_sw1_coeff_ret1[22]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[22]) );
  DFFR_X1 DP_reg_ret1_Q_reg_23_ ( .D(DP_sw1_coeff_ret1[23]), .CK(clk), .RN(
        n1138), .Q(DP_ret1[23]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_0_ ( .D(DP_w_0_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[0]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_1_ ( .D(DP_w_1_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[1]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_2_ ( .D(DP_w_2_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[2]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_3_ ( .D(DP_w_3_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[3]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_4_ ( .D(DP_w_4_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[4]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_5_ ( .D(DP_w_5_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[5]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_6_ ( .D(DP_w_6_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[6]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_7_ ( .D(DP_w_7_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[7]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_8_ ( .D(DP_w_8_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[8]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_9_ ( .D(DP_w_9_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[9]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_10_ ( .D(DP_w_10_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[10]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_11_ ( .D(DP_w_11_), .CK(clk), .RN(n1139), .Q(
        DP_pipe00[11]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_12_ ( .D(DP_w_12_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[12]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_13_ ( .D(DP_w_13_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[13]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_14_ ( .D(DP_w_14_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[14]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_15_ ( .D(DP_w_15_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[15]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_16_ ( .D(DP_w_16_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[16]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_17_ ( .D(DP_w_17_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[17]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_18_ ( .D(DP_w_18_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[18]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_19_ ( .D(DP_w_19_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[19]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_20_ ( .D(DP_w_20_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[20]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_21_ ( .D(DP_w_21_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[21]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_22_ ( .D(DP_w_22_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[22]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_23_ ( .D(DP_w_23_), .CK(clk), .RN(n1140), .Q(
        DP_pipe00[23]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe00[0]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[0]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe00[1]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[1]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe00[2]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[2]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe00[3]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[3]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe00[4]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[4]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe00[5]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[5]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe00[6]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[6]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe00[7]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[7]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe00[8]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[8]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe00[9]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[9]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe00[10]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[10]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe00[11]), .CK(clk), 
        .RN(n1141), .Q(DP_pipe10[11]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe00[12]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[12]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe00[13]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[13]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe00[14]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[14]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe00[15]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[15]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe00[16]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[16]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe00[17]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[17]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe00[18]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[18]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe00[19]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[19]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe00[20]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[20]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe00[21]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[21]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe00[22]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[22]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe00[23]), .CK(clk), 
        .RN(n1142), .Q(DP_pipe10[23]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe01[0]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[0]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe01[1]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[1]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe01[2]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[2]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe01[3]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[3]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe01[4]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[4]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe01[5]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[5]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe01[6]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[6]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe01[7]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[7]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe01[8]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[8]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe01[9]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[9]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe01[10]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[10]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe01[11]), .CK(clk), 
        .RN(n1143), .Q(DP_pipe11[11]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe01[12]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[12]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe01[13]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[13]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe01[14]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[14]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe01[15]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[15]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe01[16]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[16]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe01[17]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[17]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe01[18]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[18]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe01[19]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[19]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe01[20]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[20]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe01[21]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[21]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe01[22]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[22]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe01[23]), .CK(clk), 
        .RN(n1144), .Q(DP_pipe11[23]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe02[0]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[0]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe02[1]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[1]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe02[2]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[2]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe02[3]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[3]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe02[4]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[4]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe02[5]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[5]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe02[6]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[6]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe02[7]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[7]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe02[8]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[8]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe02[9]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[9]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe02[10]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[10]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe02[11]), .CK(clk), 
        .RN(n1145), .Q(DP_pipe12[11]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe02[12]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[12]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe02[13]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[13]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe02[14]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[14]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe02[15]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[15]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe02[16]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[16]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe02[17]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[17]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe02[18]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[18]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe02[19]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[19]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe02[20]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[20]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe02[21]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[21]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe02[22]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[22]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe02[23]), .CK(clk), 
        .RN(n1146), .Q(DP_pipe12[23]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe03[0]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[0]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe03[1]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[1]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe03[2]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[2]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe03[3]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[3]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe03[4]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[4]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe03[5]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[5]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe03[6]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[6]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe03[7]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[7]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe03[8]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[8]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe03[9]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[9]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe03[10]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[10]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe03[11]), .CK(clk), 
        .RN(n1147), .Q(DP_pipe13[11]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe03[12]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[12]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe03[13]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[13]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe03[14]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[14]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe03[15]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[15]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe03[16]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[16]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe03[17]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[17]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe03[18]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[18]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe03[19]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[19]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe03[20]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[20]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe03[21]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[21]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe03[22]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[22]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe03[23]), .CK(clk), 
        .RN(n1148), .Q(DP_pipe13[23]) );
  DFFR_X1 CU_presentState_reg_1_ ( .D(n1026), .CK(clk), .RN(n1149), .Q(
        delayed_controls_0__1_) );
  DFFR_X1 DP_reg_sw0_Q_reg_23_ ( .D(n671), .CK(clk), .RN(n1149), .Q(DP_sw0_23_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_23_ ( .D(DP_sw0_23_), .CK(clk), .RN(n1149), .Q(
        DP_pipe01[23]) );
  DFFR_X1 DP_reg_sw0_Q_reg_22_ ( .D(n669), .CK(clk), .RN(n1149), .Q(DP_sw0_22_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_22_ ( .D(DP_sw0_22_), .CK(clk), .RN(n1149), .Q(
        DP_pipe01[22]) );
  DFFR_X1 DP_reg_sw0_Q_reg_21_ ( .D(n667), .CK(clk), .RN(n1149), .Q(DP_sw0_21_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_21_ ( .D(DP_sw0_21_), .CK(clk), .RN(n1149), .Q(
        DP_pipe01[21]) );
  DFFR_X1 DP_reg_sw0_Q_reg_20_ ( .D(n665), .CK(clk), .RN(n1149), .Q(DP_sw0_20_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_20_ ( .D(DP_sw0_20_), .CK(clk), .RN(n1149), .Q(
        DP_pipe01[20]) );
  DFFR_X1 DP_reg_sw0_Q_reg_19_ ( .D(n663), .CK(clk), .RN(n1149), .Q(DP_sw0_19_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_19_ ( .D(DP_sw0_19_), .CK(clk), .RN(n1149), .Q(
        DP_pipe01[19]) );
  DFFR_X1 DP_reg_sw0_Q_reg_18_ ( .D(n661), .CK(clk), .RN(n1149), .Q(DP_sw0_18_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_18_ ( .D(DP_sw0_18_), .CK(clk), .RN(n1150), .Q(
        DP_pipe01[18]) );
  DFFR_X1 DP_reg_sw0_Q_reg_17_ ( .D(n659), .CK(clk), .RN(n1150), .Q(DP_sw0_17_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_17_ ( .D(DP_sw0_17_), .CK(clk), .RN(n1150), .Q(
        DP_pipe01[17]) );
  DFFR_X1 DP_reg_sw0_Q_reg_16_ ( .D(n657), .CK(clk), .RN(n1150), .Q(DP_sw0_16_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_16_ ( .D(DP_sw0_16_), .CK(clk), .RN(n1150), .Q(
        DP_pipe01[16]) );
  DFFR_X1 DP_reg_sw0_Q_reg_15_ ( .D(n655), .CK(clk), .RN(n1150), .Q(DP_sw0_15_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_15_ ( .D(DP_sw0_15_), .CK(clk), .RN(n1150), .Q(
        DP_pipe01[15]) );
  DFFR_X1 DP_reg_sw0_Q_reg_14_ ( .D(n653), .CK(clk), .RN(n1150), .Q(DP_sw0_14_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_14_ ( .D(DP_sw0_14_), .CK(clk), .RN(n1150), .Q(
        DP_pipe01[14]) );
  DFFR_X1 DP_reg_sw0_Q_reg_13_ ( .D(n651), .CK(clk), .RN(n1150), .Q(DP_sw0_13_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_13_ ( .D(DP_sw0_13_), .CK(clk), .RN(n1150), .Q(
        DP_pipe01[13]) );
  DFFR_X1 DP_reg_sw0_Q_reg_12_ ( .D(n649), .CK(clk), .RN(n1150), .Q(DP_sw0_12_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_12_ ( .D(DP_sw0_12_), .CK(clk), .RN(n1151), .Q(
        DP_pipe01[12]) );
  DFFR_X1 DP_reg_sw0_Q_reg_11_ ( .D(n647), .CK(clk), .RN(n1151), .Q(DP_sw0_11_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_11_ ( .D(DP_sw0_11_), .CK(clk), .RN(n1151), .Q(
        DP_pipe01[11]) );
  DFFR_X1 DP_reg_sw0_Q_reg_10_ ( .D(n645), .CK(clk), .RN(n1151), .Q(DP_sw0_10_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_10_ ( .D(DP_sw0_10_), .CK(clk), .RN(n1151), .Q(
        DP_pipe01[10]) );
  DFFR_X1 DP_reg_sw0_Q_reg_9_ ( .D(n643), .CK(clk), .RN(n1151), .Q(DP_sw0_9_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_9_ ( .D(DP_sw0_9_), .CK(clk), .RN(n1151), .Q(
        DP_pipe01[9]) );
  DFFR_X1 DP_reg_sw0_Q_reg_8_ ( .D(n641), .CK(clk), .RN(n1151), .Q(DP_sw0_8_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_8_ ( .D(DP_sw0_8_), .CK(clk), .RN(n1151), .Q(
        DP_pipe01[8]) );
  DFFR_X1 DP_reg_sw0_Q_reg_7_ ( .D(n639), .CK(clk), .RN(n1151), .Q(DP_sw0_7_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_7_ ( .D(DP_sw0_7_), .CK(clk), .RN(n1151), .Q(
        DP_pipe01[7]) );
  DFFR_X1 DP_reg_sw0_Q_reg_6_ ( .D(n637), .CK(clk), .RN(n1151), .Q(DP_sw0_6_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_6_ ( .D(DP_sw0_6_), .CK(clk), .RN(n1152), .Q(
        DP_pipe01[6]) );
  DFFR_X1 DP_reg_sw0_Q_reg_5_ ( .D(n635), .CK(clk), .RN(n1152), .Q(DP_sw0_5_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_5_ ( .D(DP_sw0_5_), .CK(clk), .RN(n1152), .Q(
        DP_pipe01[5]) );
  DFFR_X1 DP_reg_sw0_Q_reg_4_ ( .D(n633), .CK(clk), .RN(n1152), .Q(DP_sw0_4_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_4_ ( .D(DP_sw0_4_), .CK(clk), .RN(n1152), .Q(
        DP_pipe01[4]) );
  DFFR_X1 DP_reg_sw0_Q_reg_3_ ( .D(n631), .CK(clk), .RN(n1152), .Q(DP_sw0_3_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_3_ ( .D(DP_sw0_3_), .CK(clk), .RN(n1152), .Q(
        DP_pipe01[3]) );
  DFFR_X1 DP_reg_sw0_Q_reg_2_ ( .D(n629), .CK(clk), .RN(n1152), .Q(DP_sw0_2_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_2_ ( .D(DP_sw0_2_), .CK(clk), .RN(n1152), .Q(
        DP_pipe01[2]) );
  DFFR_X1 DP_reg_sw0_Q_reg_1_ ( .D(n627), .CK(clk), .RN(n1152), .Q(DP_sw0_1_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_1_ ( .D(DP_sw0_1_), .CK(clk), .RN(n1152), .Q(
        DP_pipe01[1]) );
  DFFR_X1 DP_reg_sw0_Q_reg_0_ ( .D(n625), .CK(clk), .RN(n1152), .Q(DP_sw0_0_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_0_ ( .D(DP_sw0_0_), .CK(clk), .RN(n1153), .Q(
        DP_pipe01[0]) );
  DFFR_X1 DP_reg_sw1_Q_reg_23_ ( .D(n623), .CK(clk), .RN(n1153), .QN(n996) );
  DFFR_X1 DP_reg_pipe02_Q_reg_23_ ( .D(n1051), .CK(clk), .RN(n1153), .Q(
        DP_pipe02[23]) );
  DFFR_X1 DP_reg_sw1_Q_reg_22_ ( .D(n621), .CK(clk), .RN(n1153), .Q(DP_sw1_22_), .QN(n1015) );
  DFFR_X1 DP_reg_pipe02_Q_reg_22_ ( .D(DP_sw1_22_), .CK(clk), .RN(n1153), .Q(
        DP_pipe02[22]) );
  DFFR_X1 DP_reg_sw1_Q_reg_21_ ( .D(n619), .CK(clk), .RN(n1153), .Q(DP_sw1_21_), .QN(n1018) );
  DFFR_X1 DP_reg_pipe02_Q_reg_21_ ( .D(DP_sw1_21_), .CK(clk), .RN(n1153), .Q(
        DP_pipe02[21]) );
  DFFR_X1 DP_reg_sw1_Q_reg_20_ ( .D(n617), .CK(clk), .RN(n1153), .Q(DP_sw1_20_), .QN(n997) );
  DFFR_X1 DP_reg_pipe02_Q_reg_20_ ( .D(DP_sw1_20_), .CK(clk), .RN(n1153), .Q(
        DP_pipe02[20]) );
  DFFR_X1 DP_reg_sw1_Q_reg_19_ ( .D(n615), .CK(clk), .RN(n1153), .Q(DP_sw1_19_), .QN(n1014) );
  DFFR_X1 DP_reg_pipe02_Q_reg_19_ ( .D(DP_sw1_19_), .CK(clk), .RN(n1153), .Q(
        DP_pipe02[19]) );
  DFFR_X1 DP_reg_sw1_Q_reg_18_ ( .D(n613), .CK(clk), .RN(n1153), .Q(DP_sw1_18_), .QN(n1013) );
  DFFR_X1 DP_reg_pipe02_Q_reg_18_ ( .D(DP_sw1_18_), .CK(clk), .RN(n1154), .Q(
        DP_pipe02[18]) );
  DFFR_X1 DP_reg_sw1_Q_reg_17_ ( .D(n611), .CK(clk), .RN(n1154), .Q(DP_sw1_17_), .QN(n1012) );
  DFFR_X1 DP_reg_pipe02_Q_reg_17_ ( .D(DP_sw1_17_), .CK(clk), .RN(n1154), .Q(
        DP_pipe02[17]) );
  DFFR_X1 DP_reg_sw1_Q_reg_16_ ( .D(n609), .CK(clk), .RN(n1154), .Q(DP_sw1_16_), .QN(n1011) );
  DFFR_X1 DP_reg_pipe02_Q_reg_16_ ( .D(DP_sw1_16_), .CK(clk), .RN(n1154), .Q(
        DP_pipe02[16]) );
  DFFR_X1 DP_reg_sw1_Q_reg_15_ ( .D(n607), .CK(clk), .RN(n1154), .Q(DP_sw1_15_), .QN(n1010) );
  DFFR_X1 DP_reg_pipe02_Q_reg_15_ ( .D(DP_sw1_15_), .CK(clk), .RN(n1154), .Q(
        DP_pipe02[15]) );
  DFFR_X1 DP_reg_sw1_Q_reg_14_ ( .D(n605), .CK(clk), .RN(n1154), .Q(DP_sw1_14_), .QN(n1009) );
  DFFR_X1 DP_reg_pipe02_Q_reg_14_ ( .D(DP_sw1_14_), .CK(clk), .RN(n1154), .Q(
        DP_pipe02[14]) );
  DFFR_X1 DP_reg_sw1_Q_reg_13_ ( .D(n603), .CK(clk), .RN(n1154), .Q(DP_sw1_13_), .QN(n1008) );
  DFFR_X1 DP_reg_pipe02_Q_reg_13_ ( .D(DP_sw1_13_), .CK(clk), .RN(n1154), .Q(
        DP_pipe02[13]) );
  DFFR_X1 DP_reg_sw1_Q_reg_12_ ( .D(n601), .CK(clk), .RN(n1154), .Q(DP_sw1_12_), .QN(n1007) );
  DFFR_X1 DP_reg_pipe02_Q_reg_12_ ( .D(DP_sw1_12_), .CK(clk), .RN(n1155), .Q(
        DP_pipe02[12]) );
  DFFR_X1 DP_reg_sw1_Q_reg_11_ ( .D(n599), .CK(clk), .RN(n1155), .Q(DP_sw1_11_), .QN(n1006) );
  DFFR_X1 DP_reg_pipe02_Q_reg_11_ ( .D(DP_sw1_11_), .CK(clk), .RN(n1155), .Q(
        DP_pipe02[11]) );
  DFFR_X1 DP_reg_sw1_Q_reg_10_ ( .D(n597), .CK(clk), .RN(n1155), .Q(DP_sw1_10_), .QN(n1005) );
  DFFR_X1 DP_reg_pipe02_Q_reg_10_ ( .D(DP_sw1_10_), .CK(clk), .RN(n1155), .Q(
        DP_pipe02[10]) );
  DFFR_X1 DP_reg_sw1_Q_reg_9_ ( .D(n595), .CK(clk), .RN(n1155), .Q(DP_sw1_9_), 
        .QN(n1004) );
  DFFR_X1 DP_reg_pipe02_Q_reg_9_ ( .D(DP_sw1_9_), .CK(clk), .RN(n1155), .Q(
        DP_pipe02[9]) );
  DFFR_X1 DP_reg_sw1_Q_reg_8_ ( .D(n593), .CK(clk), .RN(n1155), .Q(DP_sw1_8_), 
        .QN(n1003) );
  DFFR_X1 DP_reg_pipe02_Q_reg_8_ ( .D(DP_sw1_8_), .CK(clk), .RN(n1155), .Q(
        DP_pipe02[8]) );
  DFFR_X1 DP_reg_sw1_Q_reg_7_ ( .D(n591), .CK(clk), .RN(n1155), .Q(DP_sw1_7_), 
        .QN(n1002) );
  DFFR_X1 DP_reg_pipe02_Q_reg_7_ ( .D(DP_sw1_7_), .CK(clk), .RN(n1155), .Q(
        DP_pipe02[7]) );
  DFFR_X1 DP_reg_sw1_Q_reg_6_ ( .D(n589), .CK(clk), .RN(n1155), .Q(DP_sw1_6_), 
        .QN(n1001) );
  DFFR_X1 DP_reg_pipe02_Q_reg_6_ ( .D(DP_sw1_6_), .CK(clk), .RN(n1156), .Q(
        DP_pipe02[6]) );
  DFFR_X1 DP_reg_sw1_Q_reg_5_ ( .D(n587), .CK(clk), .RN(n1156), .Q(DP_sw1_5_), 
        .QN(n1000) );
  DFFR_X1 DP_reg_pipe02_Q_reg_5_ ( .D(DP_sw1_5_), .CK(clk), .RN(n1156), .Q(
        DP_pipe02[5]) );
  DFFR_X1 DP_reg_sw1_Q_reg_4_ ( .D(n585), .CK(clk), .RN(n1156), .Q(DP_sw1_4_), 
        .QN(n999) );
  DFFR_X1 DP_reg_pipe02_Q_reg_4_ ( .D(DP_sw1_4_), .CK(clk), .RN(n1156), .Q(
        DP_pipe02[4]) );
  DFFR_X1 DP_reg_sw1_Q_reg_3_ ( .D(n583), .CK(clk), .RN(n1156), .Q(DP_sw1_3_), 
        .QN(n998) );
  DFFR_X1 DP_reg_pipe02_Q_reg_3_ ( .D(DP_sw1_3_), .CK(clk), .RN(n1156), .Q(
        DP_pipe02[3]) );
  DFFR_X1 DP_reg_sw1_Q_reg_2_ ( .D(n581), .CK(clk), .RN(n1156), .Q(DP_sw1_2_), 
        .QN(n1016) );
  DFFR_X1 DP_reg_pipe02_Q_reg_2_ ( .D(DP_sw1_2_), .CK(clk), .RN(n1156), .Q(
        DP_pipe02[2]) );
  DFFR_X1 DP_reg_sw1_Q_reg_1_ ( .D(n579), .CK(clk), .RN(n1156), .Q(DP_sw1_1_), 
        .QN(n1017) );
  DFFR_X1 DP_reg_pipe02_Q_reg_1_ ( .D(DP_sw1_1_), .CK(clk), .RN(n1156), .Q(
        DP_pipe02[1]) );
  DFFR_X1 DP_reg_sw1_Q_reg_0_ ( .D(n577), .CK(clk), .RN(n1156), .Q(DP_sw1_0_), 
        .QN(n1019) );
  DFFR_X1 DP_reg_pipe02_Q_reg_0_ ( .D(DP_sw1_0_), .CK(clk), .RN(n1157), .Q(
        DP_pipe02[0]) );
  DFFR_X1 DP_reg_sw2_Q_reg_23_ ( .D(n575), .CK(clk), .RN(n1157), .Q(DP_sw2[23]), .QN(n307) );
  DFFR_X1 DP_reg_pipe03_Q_reg_23_ ( .D(DP_sw2[23]), .CK(clk), .RN(n1157), .Q(
        DP_pipe03[23]) );
  DFFR_X1 DP_reg_sw2_Q_reg_22_ ( .D(n573), .CK(clk), .RN(n1157), .Q(DP_sw2[22]), .QN(n306) );
  DFFR_X1 DP_reg_pipe03_Q_reg_22_ ( .D(DP_sw2[22]), .CK(clk), .RN(n1157), .Q(
        DP_pipe03[22]) );
  DFFR_X1 DP_reg_sw2_Q_reg_21_ ( .D(n571), .CK(clk), .RN(n1157), .Q(DP_sw2[21]), .QN(n305) );
  DFFR_X1 DP_reg_pipe03_Q_reg_21_ ( .D(DP_sw2[21]), .CK(clk), .RN(n1157), .Q(
        DP_pipe03[21]) );
  DFFR_X1 DP_reg_sw2_Q_reg_20_ ( .D(n569), .CK(clk), .RN(n1157), .Q(DP_sw2[20]), .QN(n304) );
  DFFR_X1 DP_reg_pipe03_Q_reg_20_ ( .D(DP_sw2[20]), .CK(clk), .RN(n1157), .Q(
        DP_pipe03[20]) );
  DFFR_X1 DP_reg_sw2_Q_reg_19_ ( .D(n567), .CK(clk), .RN(n1157), .Q(DP_sw2[19]), .QN(n303) );
  DFFR_X1 DP_reg_pipe03_Q_reg_19_ ( .D(DP_sw2[19]), .CK(clk), .RN(n1157), .Q(
        DP_pipe03[19]) );
  DFFR_X1 DP_reg_sw2_Q_reg_18_ ( .D(n565), .CK(clk), .RN(n1157), .Q(DP_sw2[18]), .QN(n302) );
  DFFR_X1 DP_reg_pipe03_Q_reg_18_ ( .D(DP_sw2[18]), .CK(clk), .RN(n1158), .Q(
        DP_pipe03[18]) );
  DFFR_X1 DP_reg_sw2_Q_reg_17_ ( .D(n563), .CK(clk), .RN(n1158), .Q(DP_sw2[17]), .QN(n301) );
  DFFR_X1 DP_reg_pipe03_Q_reg_17_ ( .D(DP_sw2[17]), .CK(clk), .RN(n1158), .Q(
        DP_pipe03[17]) );
  DFFR_X1 DP_reg_sw2_Q_reg_16_ ( .D(n561), .CK(clk), .RN(n1158), .Q(DP_sw2[16]), .QN(n300) );
  DFFR_X1 DP_reg_pipe03_Q_reg_16_ ( .D(DP_sw2[16]), .CK(clk), .RN(n1158), .Q(
        DP_pipe03[16]) );
  DFFR_X1 DP_reg_sw2_Q_reg_15_ ( .D(n559), .CK(clk), .RN(n1158), .Q(DP_sw2[15]), .QN(n299) );
  DFFR_X1 DP_reg_pipe03_Q_reg_15_ ( .D(DP_sw2[15]), .CK(clk), .RN(n1158), .Q(
        DP_pipe03[15]) );
  DFFR_X1 DP_reg_sw2_Q_reg_14_ ( .D(n557), .CK(clk), .RN(n1158), .Q(DP_sw2[14]), .QN(n298) );
  DFFR_X1 DP_reg_pipe03_Q_reg_14_ ( .D(DP_sw2[14]), .CK(clk), .RN(n1158), .Q(
        DP_pipe03[14]) );
  DFFR_X1 DP_reg_sw2_Q_reg_13_ ( .D(n555), .CK(clk), .RN(n1158), .Q(DP_sw2[13]), .QN(n297) );
  DFFR_X1 DP_reg_pipe03_Q_reg_13_ ( .D(DP_sw2[13]), .CK(clk), .RN(n1158), .Q(
        DP_pipe03[13]) );
  DFFR_X1 DP_reg_sw2_Q_reg_12_ ( .D(n553), .CK(clk), .RN(n1158), .Q(DP_sw2[12]), .QN(n296) );
  DFFR_X1 DP_reg_pipe03_Q_reg_12_ ( .D(DP_sw2[12]), .CK(clk), .RN(n1159), .Q(
        DP_pipe03[12]) );
  DFFR_X1 DP_reg_sw2_Q_reg_11_ ( .D(n551), .CK(clk), .RN(n1159), .Q(DP_sw2[11]), .QN(n295) );
  DFFR_X1 DP_reg_pipe03_Q_reg_11_ ( .D(DP_sw2[11]), .CK(clk), .RN(n1159), .Q(
        DP_pipe03[11]) );
  DFFR_X1 DP_reg_sw2_Q_reg_10_ ( .D(n549), .CK(clk), .RN(n1159), .Q(DP_sw2[10]), .QN(n294) );
  DFFR_X1 DP_reg_pipe03_Q_reg_10_ ( .D(DP_sw2[10]), .CK(clk), .RN(n1159), .Q(
        DP_pipe03[10]) );
  DFFR_X1 DP_reg_sw2_Q_reg_9_ ( .D(n547), .CK(clk), .RN(n1159), .Q(DP_sw2[9]), 
        .QN(n293) );
  DFFR_X1 DP_reg_pipe03_Q_reg_9_ ( .D(DP_sw2[9]), .CK(clk), .RN(n1159), .Q(
        DP_pipe03[9]) );
  DFFR_X1 DP_reg_sw2_Q_reg_8_ ( .D(n545), .CK(clk), .RN(n1159), .Q(DP_sw2[8]), 
        .QN(n292) );
  DFFR_X1 DP_reg_pipe03_Q_reg_8_ ( .D(DP_sw2[8]), .CK(clk), .RN(n1159), .Q(
        DP_pipe03[8]) );
  DFFR_X1 DP_reg_sw2_Q_reg_7_ ( .D(n543), .CK(clk), .RN(n1159), .Q(DP_sw2[7]), 
        .QN(n291) );
  DFFR_X1 DP_reg_pipe03_Q_reg_7_ ( .D(DP_sw2[7]), .CK(clk), .RN(n1159), .Q(
        DP_pipe03[7]) );
  DFFR_X1 DP_reg_sw2_Q_reg_6_ ( .D(n541), .CK(clk), .RN(n1159), .Q(DP_sw2[6]), 
        .QN(n290) );
  DFFR_X1 DP_reg_pipe03_Q_reg_6_ ( .D(DP_sw2[6]), .CK(clk), .RN(n1160), .Q(
        DP_pipe03[6]) );
  DFFR_X1 DP_reg_sw2_Q_reg_5_ ( .D(n539), .CK(clk), .RN(n1160), .Q(DP_sw2[5]), 
        .QN(n289) );
  DFFR_X1 DP_reg_pipe03_Q_reg_5_ ( .D(DP_sw2[5]), .CK(clk), .RN(n1160), .Q(
        DP_pipe03[5]) );
  DFFR_X1 DP_reg_sw2_Q_reg_4_ ( .D(n537), .CK(clk), .RN(n1160), .Q(DP_sw2[4]), 
        .QN(n288) );
  DFFR_X1 DP_reg_pipe03_Q_reg_4_ ( .D(DP_sw2[4]), .CK(clk), .RN(n1160), .Q(
        DP_pipe03[4]) );
  DFFR_X1 DP_reg_sw2_Q_reg_3_ ( .D(n535), .CK(clk), .RN(n1160), .Q(DP_sw2[3]), 
        .QN(n287) );
  DFFR_X1 DP_reg_pipe03_Q_reg_3_ ( .D(DP_sw2[3]), .CK(clk), .RN(n1160), .Q(
        DP_pipe03[3]) );
  DFFR_X1 DP_reg_sw2_Q_reg_2_ ( .D(n533), .CK(clk), .RN(n1160), .Q(DP_sw2[2]), 
        .QN(n286) );
  DFFR_X1 DP_reg_pipe03_Q_reg_2_ ( .D(DP_sw2[2]), .CK(clk), .RN(n1160), .Q(
        DP_pipe03[2]) );
  DFFR_X1 DP_reg_sw2_Q_reg_1_ ( .D(n531), .CK(clk), .RN(n1160), .Q(DP_sw2[1]), 
        .QN(n285) );
  DFFR_X1 DP_reg_pipe03_Q_reg_1_ ( .D(DP_sw2[1]), .CK(clk), .RN(n1160), .Q(
        DP_pipe03[1]) );
  DFFR_X1 DP_reg_sw2_Q_reg_0_ ( .D(n529), .CK(clk), .RN(n1160), .Q(DP_sw2[0]), 
        .QN(n284) );
  DFFR_X1 DP_reg_pipe03_Q_reg_0_ ( .D(DP_sw2[0]), .CK(clk), .RN(n1161), .Q(
        DP_pipe03[0]) );
  DFFR_X1 CU_presentState_reg_0_ ( .D(CU_nextState_0_), .CK(clk), .RN(n1161), 
        .QN(n283) );
  DFFR_X1 reg_delay_0_Q_reg_0_ ( .D(delayed_controls_0__1_), .CK(clk), .RN(
        n1161), .Q(delayed_controls_1__1_) );
  DFFR_X1 reg_delay_0_Q_reg_1_ ( .D(n1026), .CK(clk), .RN(n1161), .Q(
        delayed_controls_1__0_) );
  DFFR_X1 reg_delay_1_Q_reg_0_ ( .D(delayed_controls_1__1_), .CK(clk), .RN(
        n1161), .Q(vOut) );
  DFFR_X1 reg_delay_1_Q_reg_1_ ( .D(delayed_controls_1__0_), .CK(clk), .RN(
        n1161), .Q(delayed_controls_2__0_), .QN(n1020) );
  DFFR_X1 DP_reg_out_Q_reg_11_ ( .D(n524), .CK(clk), .RN(n1161), .Q(dOut[11]), 
        .QN(n281) );
  DFFR_X1 DP_reg_out_Q_reg_10_ ( .D(n523), .CK(clk), .RN(n1161), .Q(dOut[10]), 
        .QN(n280) );
  DFFR_X1 DP_reg_out_Q_reg_9_ ( .D(n522), .CK(clk), .RN(n1161), .Q(dOut[9]), 
        .QN(n279) );
  DFFR_X1 DP_reg_out_Q_reg_8_ ( .D(n521), .CK(clk), .RN(n1161), .Q(dOut[8]), 
        .QN(n278) );
  DFFR_X1 DP_reg_out_Q_reg_7_ ( .D(n520), .CK(clk), .RN(n1161), .Q(dOut[7]), 
        .QN(n277) );
  DFFR_X1 DP_reg_out_Q_reg_6_ ( .D(n519), .CK(clk), .RN(n1161), .Q(dOut[6]), 
        .QN(n276) );
  DFFR_X1 DP_reg_out_Q_reg_5_ ( .D(n518), .CK(clk), .RN(n1162), .Q(dOut[5]), 
        .QN(n275) );
  DFFR_X1 DP_reg_out_Q_reg_4_ ( .D(n517), .CK(clk), .RN(n1162), .Q(dOut[4]), 
        .QN(n274) );
  DFFR_X1 DP_reg_out_Q_reg_3_ ( .D(n516), .CK(clk), .RN(n1162), .Q(dOut[3]), 
        .QN(n273) );
  DFFR_X1 DP_reg_out_Q_reg_2_ ( .D(n515), .CK(clk), .RN(n1162), .Q(dOut[2]), 
        .QN(n272) );
  DFFR_X1 DP_reg_out_Q_reg_1_ ( .D(n514), .CK(clk), .RN(n1162), .Q(dOut[1]), 
        .QN(n271) );
  DFFR_X1 DP_reg_out_Q_reg_0_ ( .D(n513), .CK(clk), .RN(n1162), .Q(dOut[0]), 
        .QN(n270) );
  XOR2_X1 U491 ( .A(n1091), .B(n1026), .Z(CU_nextState_0_) );
  XOR2_X1 U493 ( .A(n283), .B(delayed_controls_0__1_), .Z(n40) );
  iir_filter_DW01_add_3 add_1_root_sub_0_root_DP_sub_217 ( .A({DP_ret0[23], 
        DP_ret0[22], DP_ret0[21], DP_ret0[20], DP_ret0[19], DP_ret0[18], 
        DP_ret0[17], DP_ret0[16], DP_ret0[15], DP_ret0[14], DP_ret0[13], 
        DP_ret0[12], DP_ret0[11], DP_ret0[10], DP_ret0[9], DP_ret0[8], 
        DP_ret0[7], DP_ret0[6], DP_ret0[5], DP_ret0[4], DP_ret0[3], DP_ret0[2], 
        DP_ret0[1], DP_ret0[0]}), .B({DP_ret1[23], DP_ret1[22], DP_ret1[21], 
        DP_ret1[20], DP_ret1[19], DP_ret1[18], DP_ret1[17], DP_ret1[16], 
        DP_ret1[15], DP_ret1[14], DP_ret1[13], DP_ret1[12], DP_ret1[11], 
        DP_ret1[10], DP_ret1[9], DP_ret1[8], DP_ret1[7], DP_ret1[6], 
        DP_ret1[5], DP_ret1[4], DP_ret1[3], DP_ret1[2], DP_ret1[1], DP_ret1[0]}), .CI(1'b0), .SUM({DP_fb_23_, DP_fb_22_, DP_fb_21_, DP_fb_20_, DP_fb_19_, 
        DP_fb_18_, DP_fb_17_, DP_fb_16_, DP_fb_15_, DP_fb_14_, DP_fb_13_, 
        DP_fb_12_, DP_fb_11_, DP_fb_10_, DP_fb_9_, DP_fb_8_, DP_fb_7_, 
        DP_fb_6_, DP_fb_5_, DP_fb_4_, DP_fb_3_, DP_fb_2_, DP_fb_1_, DP_fb_0_})
         );
  iir_filter_DW01_sub_0 sub_0_root_sub_0_root_DP_sub_217 ( .A({DP_x[11], 
        DP_x[11], DP_x[10], DP_x[9], DP_x[8], DP_x[7], DP_x[6], DP_x[5], 
        DP_x[4], DP_x[3], DP_x[2], DP_x[1], DP_x[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({DP_fb_23_, DP_fb_22_, 
        DP_fb_21_, DP_fb_20_, DP_fb_19_, DP_fb_18_, DP_fb_17_, DP_fb_16_, 
        DP_fb_15_, DP_fb_14_, DP_fb_13_, DP_fb_12_, DP_fb_11_, DP_fb_10_, 
        DP_fb_9_, DP_fb_8_, DP_fb_7_, DP_fb_6_, DP_fb_5_, DP_fb_4_, DP_fb_3_, 
        DP_fb_2_, DP_fb_1_, DP_fb_0_}), .CI(1'b0), .DIFF({DP_w_23_, DP_w_22_, 
        DP_w_21_, DP_w_20_, DP_w_19_, DP_w_18_, DP_w_17_, DP_w_16_, DP_w_15_, 
        DP_w_14_, DP_w_13_, DP_w_12_, DP_w_11_, DP_w_10_, DP_w_9_, DP_w_8_, 
        DP_w_7_, DP_w_6_, DP_w_5_, DP_w_4_, DP_w_3_, DP_w_2_, DP_w_1_, DP_w_0_}) );
  iir_filter_DW01_add_2 add_2_root_add_0_root_DP_add_223 ( .A({DP_pipe11[23], 
        DP_pipe11[22], DP_pipe11[21], DP_pipe11[20], DP_pipe11[19], 
        DP_pipe11[18], DP_pipe11[17], DP_pipe11[16], DP_pipe11[15], 
        DP_pipe11[14], DP_pipe11[13], DP_pipe11[12], DP_pipe11[11], 
        DP_pipe11[10], DP_pipe11[9], DP_pipe11[8], DP_pipe11[7], DP_pipe11[6], 
        DP_pipe11[5], DP_pipe11[4], DP_pipe11[3], DP_pipe11[2], DP_pipe11[1], 
        DP_pipe11[0]}), .B({DP_pipe13[23], DP_pipe13[22], DP_pipe13[21], 
        DP_pipe13[20], DP_pipe13[19], DP_pipe13[18], DP_pipe13[17], 
        DP_pipe13[16], DP_pipe13[15], DP_pipe13[14], DP_pipe13[13], 
        DP_pipe13[12], DP_pipe13[11], DP_pipe13[10], DP_pipe13[9], 
        DP_pipe13[8], DP_pipe13[7], DP_pipe13[6], DP_pipe13[5], DP_pipe13[4], 
        DP_pipe13[3], DP_pipe13[2], DP_pipe13[1], DP_pipe13[0]}), .CI(1'b0), 
        .SUM({DP_ff_23_, DP_ff_22_, DP_ff_21_, DP_ff_20_, DP_ff_19_, DP_ff_18_, 
        DP_ff_17_, DP_ff_16_, DP_ff_15_, DP_ff_14_, DP_ff_13_, DP_ff_12_, 
        DP_ff_11_, DP_ff_10_, DP_ff_9_, DP_ff_8_, DP_ff_7_, DP_ff_6_, DP_ff_5_, 
        DP_ff_4_, DP_ff_3_, DP_ff_2_, DP_ff_1_, DP_ff_0_}) );
  iir_filter_DW01_add_1 add_1_root_add_0_root_DP_add_223 ( .A({DP_pipe10[23], 
        DP_pipe10[22], DP_pipe10[21], DP_pipe10[20], DP_pipe10[19], 
        DP_pipe10[18], DP_pipe10[17], DP_pipe10[16], DP_pipe10[15], 
        DP_pipe10[14], DP_pipe10[13], DP_pipe10[12], DP_pipe10[11], 
        DP_pipe10[10], DP_pipe10[9], DP_pipe10[8], DP_pipe10[7], DP_pipe10[6], 
        DP_pipe10[5], DP_pipe10[4], DP_pipe10[3], DP_pipe10[2], DP_pipe10[1], 
        DP_pipe10[0]}), .B({DP_pipe12[23], DP_pipe12[22], DP_pipe12[21], 
        DP_pipe12[20], DP_pipe12[19], DP_pipe12[18], DP_pipe12[17], 
        DP_pipe12[16], DP_pipe12[15], DP_pipe12[14], DP_pipe12[13], 
        DP_pipe12[12], DP_pipe12[11], DP_pipe12[10], DP_pipe12[9], 
        DP_pipe12[8], DP_pipe12[7], DP_pipe12[6], DP_pipe12[5], DP_pipe12[4], 
        DP_pipe12[3], DP_pipe12[2], DP_pipe12[1], DP_pipe12[0]}), .CI(1'b0), 
        .SUM({DP_ff_part_23_, DP_ff_part_22_, DP_ff_part_21_, DP_ff_part_20_, 
        DP_ff_part_19_, DP_ff_part_18_, DP_ff_part_17_, DP_ff_part_16_, 
        DP_ff_part_15_, DP_ff_part_14_, DP_ff_part_13_, DP_ff_part_12_, 
        DP_ff_part_11_, DP_ff_part_10_, DP_ff_part_9_, DP_ff_part_8_, 
        DP_ff_part_7_, DP_ff_part_6_, DP_ff_part_5_, DP_ff_part_4_, 
        DP_ff_part_3_, DP_ff_part_2_, DP_ff_part_1_, DP_ff_part_0_}) );
  iir_filter_DW01_add_0 add_0_root_add_0_root_DP_add_223 ( .A({DP_ff_23_, 
        DP_ff_22_, DP_ff_21_, DP_ff_20_, DP_ff_19_, DP_ff_18_, DP_ff_17_, 
        DP_ff_16_, DP_ff_15_, DP_ff_14_, DP_ff_13_, DP_ff_12_, DP_ff_11_, 
        DP_ff_10_, DP_ff_9_, DP_ff_8_, DP_ff_7_, DP_ff_6_, DP_ff_5_, DP_ff_4_, 
        DP_ff_3_, DP_ff_2_, DP_ff_1_, DP_ff_0_}), .B({DP_ff_part_23_, 
        DP_ff_part_22_, DP_ff_part_21_, DP_ff_part_20_, DP_ff_part_19_, 
        DP_ff_part_18_, DP_ff_part_17_, DP_ff_part_16_, DP_ff_part_15_, 
        DP_ff_part_14_, DP_ff_part_13_, DP_ff_part_12_, DP_ff_part_11_, 
        DP_ff_part_10_, DP_ff_part_9_, DP_ff_part_8_, DP_ff_part_7_, 
        DP_ff_part_6_, DP_ff_part_5_, DP_ff_part_4_, DP_ff_part_3_, 
        DP_ff_part_2_, DP_ff_part_1_, DP_ff_part_0_}), .CI(1'b0), .SUM({
        DP_y_23, DP_y_11_, DP_y_10_, DP_y_9_, DP_y_8_, DP_y_7_, DP_y_6_, 
        DP_y_5_, DP_y_4_, DP_y_3_, DP_y_2_, DP_y_1_, DP_y_0_, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  iir_filter_DW_mult_tc_5 DP_mult_204 ( .a({DP_coeffs_fb_int[0], 
        DP_coeffs_fb_int[1], DP_coeffs_fb_int[2], DP_coeffs_fb_int[3], 
        DP_coeffs_fb_int[4], DP_coeffs_fb_int[5], DP_coeffs_fb_int[6], 
        DP_coeffs_fb_int[7], DP_coeffs_fb_int[8], DP_coeffs_fb_int[9], 
        DP_coeffs_fb_int[10], DP_coeffs_fb_int[11], DP_coeffs_fb_int[12], 
        DP_coeffs_fb_int[13], DP_coeffs_fb_int[14], DP_coeffs_fb_int[15], 
        DP_coeffs_fb_int[16], DP_coeffs_fb_int[17], DP_coeffs_fb_int[18], 
        DP_coeffs_fb_int[19], DP_coeffs_fb_int[20], DP_coeffs_fb_int[21], 
        DP_coeffs_fb_int[22], DP_coeffs_fb_int[23]}), .b({DP_sw0_23_, 
        DP_sw0_22_, DP_sw0_21_, DP_sw0_20_, DP_sw0_19_, DP_sw0_18_, DP_sw0_17_, 
        DP_sw0_16_, DP_sw0_15_, DP_sw0_14_, DP_sw0_13_, DP_sw0_12_, DP_sw0_11_, 
        DP_sw0_10_, DP_sw0_9_, DP_sw0_8_, DP_sw0_7_, DP_sw0_6_, DP_sw0_5_, 
        DP_sw0_4_, DP_sw0_3_, DP_sw0_2_, DP_sw0_1_, DP_sw0_0_}), .product({
        DP_sw0_coeff_ret0[23], SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, DP_sw0_coeff_ret0[22], DP_sw0_coeff_ret0[21], 
        DP_sw0_coeff_ret0[20], DP_sw0_coeff_ret0[19], DP_sw0_coeff_ret0[18], 
        DP_sw0_coeff_ret0[17], DP_sw0_coeff_ret0[16], DP_sw0_coeff_ret0[15], 
        DP_sw0_coeff_ret0[14], DP_sw0_coeff_ret0[13], DP_sw0_coeff_ret0[12], 
        DP_sw0_coeff_ret0[11], DP_sw0_coeff_ret0[10], DP_sw0_coeff_ret0[9], 
        DP_sw0_coeff_ret0[8], DP_sw0_coeff_ret0[7], DP_sw0_coeff_ret0[6], 
        DP_sw0_coeff_ret0[5], DP_sw0_coeff_ret0[4], DP_sw0_coeff_ret0[3], 
        DP_sw0_coeff_ret0[2], DP_sw0_coeff_ret0[1], DP_sw0_coeff_ret0[0], 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34}) );
  iir_filter_DW_mult_tc_4 DP_mult_205 ( .a({DP_coeffs_fb_int[24], 
        DP_coeffs_fb_int[25], DP_coeffs_fb_int[26], DP_coeffs_fb_int[27], 
        DP_coeffs_fb_int[28], DP_coeffs_fb_int[29], DP_coeffs_fb_int[30], 
        DP_coeffs_fb_int[31], DP_coeffs_fb_int[32], DP_coeffs_fb_int[33], 
        DP_coeffs_fb_int[34], DP_coeffs_fb_int[35], DP_coeffs_fb_int[36], 
        DP_coeffs_fb_int[37], DP_coeffs_fb_int[38], DP_coeffs_fb_int[39], 
        DP_coeffs_fb_int[40], DP_coeffs_fb_int[41], DP_coeffs_fb_int[42], 
        DP_coeffs_fb_int[43], DP_coeffs_fb_int[44], DP_coeffs_fb_int[45], 
        DP_coeffs_fb_int[46], DP_coeffs_fb_int[47]}), .b({n1051, DP_sw1_22_, 
        DP_sw1_21_, DP_sw1_20_, DP_sw1_19_, DP_sw1_18_, DP_sw1_17_, DP_sw1_16_, 
        DP_sw1_15_, DP_sw1_14_, DP_sw1_13_, DP_sw1_12_, DP_sw1_11_, DP_sw1_10_, 
        DP_sw1_9_, DP_sw1_8_, DP_sw1_7_, DP_sw1_6_, DP_sw1_5_, DP_sw1_4_, 
        DP_sw1_3_, DP_sw1_2_, DP_sw1_1_, DP_sw1_0_}), .product({
        DP_sw1_coeff_ret1[23], SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, DP_sw1_coeff_ret1[22], DP_sw1_coeff_ret1[21], 
        DP_sw1_coeff_ret1[20], DP_sw1_coeff_ret1[19], DP_sw1_coeff_ret1[18], 
        DP_sw1_coeff_ret1[17], DP_sw1_coeff_ret1[16], DP_sw1_coeff_ret1[15], 
        DP_sw1_coeff_ret1[14], DP_sw1_coeff_ret1[13], DP_sw1_coeff_ret1[12], 
        DP_sw1_coeff_ret1[11], DP_sw1_coeff_ret1[10], DP_sw1_coeff_ret1[9], 
        DP_sw1_coeff_ret1[8], DP_sw1_coeff_ret1[7], DP_sw1_coeff_ret1[6], 
        DP_sw1_coeff_ret1[5], DP_sw1_coeff_ret1[4], DP_sw1_coeff_ret1[3], 
        DP_sw1_coeff_ret1[2], DP_sw1_coeff_ret1[1], DP_sw1_coeff_ret1[0], 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58}) );
  iir_filter_DW_mult_tc_3 DP_mult_206 ( .a({DP_coeffs_ff_int[0], 
        DP_coeffs_ff_int[1], DP_coeffs_ff_int[2], DP_coeffs_ff_int[3], 
        DP_coeffs_ff_int[4], DP_coeffs_ff_int[5], DP_coeffs_ff_int[6], 
        DP_coeffs_ff_int[7], DP_coeffs_ff_int[8], DP_coeffs_ff_int[9], 
        DP_coeffs_ff_int[10], DP_coeffs_ff_int[11], DP_coeffs_ff_int[12], 
        DP_coeffs_ff_int[13], DP_coeffs_ff_int[14], DP_coeffs_ff_int[15], 
        DP_coeffs_ff_int[16], DP_coeffs_ff_int[17], DP_coeffs_ff_int[18], 
        DP_coeffs_ff_int[19], DP_coeffs_ff_int[20], DP_coeffs_ff_int[21], 
        DP_coeffs_ff_int[22], DP_coeffs_ff_int[23]}), .b({DP_pipe00[23], 
        DP_pipe00[22], DP_pipe00[21], DP_pipe00[20], DP_pipe00[19], 
        DP_pipe00[18], DP_pipe00[17], DP_pipe00[16], DP_pipe00[15], 
        DP_pipe00[14], DP_pipe00[13], DP_pipe00[12], DP_pipe00[11], 
        DP_pipe00[10], DP_pipe00[9], DP_pipe00[8], DP_pipe00[7], DP_pipe00[6], 
        DP_pipe00[5], DP_pipe00[4], DP_pipe00[3], DP_pipe00[2], DP_pipe00[1], 
        DP_pipe00[0]}), .product({DP_pipe0_coeff_pipe00[23], 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        DP_pipe0_coeff_pipe00[22], DP_pipe0_coeff_pipe00[21], 
        DP_pipe0_coeff_pipe00[20], DP_pipe0_coeff_pipe00[19], 
        DP_pipe0_coeff_pipe00[18], DP_pipe0_coeff_pipe00[17], 
        DP_pipe0_coeff_pipe00[16], DP_pipe0_coeff_pipe00[15], 
        DP_pipe0_coeff_pipe00[14], DP_pipe0_coeff_pipe00[13], 
        DP_pipe0_coeff_pipe00[12], DP_pipe0_coeff_pipe00[11], 
        DP_pipe0_coeff_pipe00[10], DP_pipe0_coeff_pipe00[9], 
        DP_pipe0_coeff_pipe00[8], DP_pipe0_coeff_pipe00[7], 
        DP_pipe0_coeff_pipe00[6], DP_pipe0_coeff_pipe00[5], 
        DP_pipe0_coeff_pipe00[4], DP_pipe0_coeff_pipe00[3], 
        DP_pipe0_coeff_pipe00[2], DP_pipe0_coeff_pipe00[1], 
        DP_pipe0_coeff_pipe00[0], SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82}) );
  iir_filter_DW_mult_tc_2 DP_mult_207 ( .a({DP_coeffs_ff_int[24], 
        DP_coeffs_ff_int[25], DP_coeffs_ff_int[26], DP_coeffs_ff_int[27], 
        DP_coeffs_ff_int[28], DP_coeffs_ff_int[29], DP_coeffs_ff_int[30], 
        DP_coeffs_ff_int[31], DP_coeffs_ff_int[32], DP_coeffs_ff_int[33], 
        DP_coeffs_ff_int[34], DP_coeffs_ff_int[35], DP_coeffs_ff_int[36], 
        DP_coeffs_ff_int[37], DP_coeffs_ff_int[38], DP_coeffs_ff_int[39], 
        DP_coeffs_ff_int[40], DP_coeffs_ff_int[41], DP_coeffs_ff_int[42], 
        DP_coeffs_ff_int[43], DP_coeffs_ff_int[44], DP_coeffs_ff_int[45], 
        DP_coeffs_ff_int[46], DP_coeffs_ff_int[47]}), .b({DP_pipe01[23], 
        DP_pipe01[22], DP_pipe01[21], DP_pipe01[20], DP_pipe01[19], 
        DP_pipe01[18], DP_pipe01[17], DP_pipe01[16], DP_pipe01[15], 
        DP_pipe01[14], DP_pipe01[13], DP_pipe01[12], DP_pipe01[11], 
        DP_pipe01[10], DP_pipe01[9], DP_pipe01[8], DP_pipe01[7], DP_pipe01[6], 
        DP_pipe01[5], DP_pipe01[4], DP_pipe01[3], DP_pipe01[2], DP_pipe01[1], 
        DP_pipe01[0]}), .product({DP_pipe0_coeff_pipe01[23], 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        DP_pipe0_coeff_pipe01[22], DP_pipe0_coeff_pipe01[21], 
        DP_pipe0_coeff_pipe01[20], DP_pipe0_coeff_pipe01[19], 
        DP_pipe0_coeff_pipe01[18], DP_pipe0_coeff_pipe01[17], 
        DP_pipe0_coeff_pipe01[16], DP_pipe0_coeff_pipe01[15], 
        DP_pipe0_coeff_pipe01[14], DP_pipe0_coeff_pipe01[13], 
        DP_pipe0_coeff_pipe01[12], DP_pipe0_coeff_pipe01[11], 
        DP_pipe0_coeff_pipe01[10], DP_pipe0_coeff_pipe01[9], 
        DP_pipe0_coeff_pipe01[8], DP_pipe0_coeff_pipe01[7], 
        DP_pipe0_coeff_pipe01[6], DP_pipe0_coeff_pipe01[5], 
        DP_pipe0_coeff_pipe01[4], DP_pipe0_coeff_pipe01[3], 
        DP_pipe0_coeff_pipe01[2], DP_pipe0_coeff_pipe01[1], 
        DP_pipe0_coeff_pipe01[0], SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106}) );
  iir_filter_DW_mult_tc_1 DP_mult_208 ( .a({DP_coeffs_ff_int[48], 
        DP_coeffs_ff_int[49], DP_coeffs_ff_int[50], DP_coeffs_ff_int[51], 
        DP_coeffs_ff_int[52], DP_coeffs_ff_int[53], DP_coeffs_ff_int[54], 
        DP_coeffs_ff_int[55], DP_coeffs_ff_int[56], DP_coeffs_ff_int[57], 
        DP_coeffs_ff_int[58], DP_coeffs_ff_int[59], DP_coeffs_ff_int[60], 
        DP_coeffs_ff_int[61], DP_coeffs_ff_int[62], DP_coeffs_ff_int[63], 
        DP_coeffs_ff_int[64], DP_coeffs_ff_int[65], DP_coeffs_ff_int[66], 
        DP_coeffs_ff_int[67], DP_coeffs_ff_int[68], DP_coeffs_ff_int[69], 
        DP_coeffs_ff_int[70], DP_coeffs_ff_int[71]}), .b({DP_pipe02[23], 
        DP_pipe02[22], DP_pipe02[21], DP_pipe02[20], DP_pipe02[19], 
        DP_pipe02[18], DP_pipe02[17], DP_pipe02[16], DP_pipe02[15], 
        DP_pipe02[14], DP_pipe02[13], DP_pipe02[12], DP_pipe02[11], 
        DP_pipe02[10], DP_pipe02[9], DP_pipe02[8], DP_pipe02[7], DP_pipe02[6], 
        DP_pipe02[5], DP_pipe02[4], DP_pipe02[3], DP_pipe02[2], DP_pipe02[1], 
        DP_pipe02[0]}), .product({DP_pipe0_coeff_pipe02[23], 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        DP_pipe0_coeff_pipe02[22], DP_pipe0_coeff_pipe02[21], 
        DP_pipe0_coeff_pipe02[20], DP_pipe0_coeff_pipe02[19], 
        DP_pipe0_coeff_pipe02[18], DP_pipe0_coeff_pipe02[17], 
        DP_pipe0_coeff_pipe02[16], DP_pipe0_coeff_pipe02[15], 
        DP_pipe0_coeff_pipe02[14], DP_pipe0_coeff_pipe02[13], 
        DP_pipe0_coeff_pipe02[12], DP_pipe0_coeff_pipe02[11], 
        DP_pipe0_coeff_pipe02[10], DP_pipe0_coeff_pipe02[9], 
        DP_pipe0_coeff_pipe02[8], DP_pipe0_coeff_pipe02[7], 
        DP_pipe0_coeff_pipe02[6], DP_pipe0_coeff_pipe02[5], 
        DP_pipe0_coeff_pipe02[4], DP_pipe0_coeff_pipe02[3], 
        DP_pipe0_coeff_pipe02[2], DP_pipe0_coeff_pipe02[1], 
        DP_pipe0_coeff_pipe02[0], SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130}) );
  iir_filter_DW_mult_tc_0 DP_mult_209 ( .a({DP_coeffs_ff_int[72], 
        DP_coeffs_ff_int[73], DP_coeffs_ff_int[74], DP_coeffs_ff_int[75], 
        DP_coeffs_ff_int[76], DP_coeffs_ff_int[77], DP_coeffs_ff_int[78], 
        DP_coeffs_ff_int[79], DP_coeffs_ff_int[80], DP_coeffs_ff_int[81], 
        DP_coeffs_ff_int[82], DP_coeffs_ff_int[83], DP_coeffs_ff_int[84], 
        DP_coeffs_ff_int[85], DP_coeffs_ff_int[86], DP_coeffs_ff_int[87], 
        DP_coeffs_ff_int[88], DP_coeffs_ff_int[89], DP_coeffs_ff_int[90], 
        DP_coeffs_ff_int[91], DP_coeffs_ff_int[92], DP_coeffs_ff_int[93], 
        DP_coeffs_ff_int[94], DP_coeffs_ff_int[95]}), .b({DP_pipe03[23], 
        DP_pipe03[22], DP_pipe03[21], DP_pipe03[20], DP_pipe03[19], 
        DP_pipe03[18], DP_pipe03[17], DP_pipe03[16], DP_pipe03[15], 
        DP_pipe03[14], DP_pipe03[13], DP_pipe03[12], DP_pipe03[11], 
        DP_pipe03[10], DP_pipe03[9], DP_pipe03[8], DP_pipe03[7], DP_pipe03[6], 
        DP_pipe03[5], DP_pipe03[4], DP_pipe03[3], DP_pipe03[2], DP_pipe03[1], 
        DP_pipe03[0]}), .product({DP_pipe0_coeff_pipe03[23], 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        DP_pipe0_coeff_pipe03[22], DP_pipe0_coeff_pipe03[21], 
        DP_pipe0_coeff_pipe03[20], DP_pipe0_coeff_pipe03[19], 
        DP_pipe0_coeff_pipe03[18], DP_pipe0_coeff_pipe03[17], 
        DP_pipe0_coeff_pipe03[16], DP_pipe0_coeff_pipe03[15], 
        DP_pipe0_coeff_pipe03[14], DP_pipe0_coeff_pipe03[13], 
        DP_pipe0_coeff_pipe03[12], DP_pipe0_coeff_pipe03[11], 
        DP_pipe0_coeff_pipe03[10], DP_pipe0_coeff_pipe03[9], 
        DP_pipe0_coeff_pipe03[8], DP_pipe0_coeff_pipe03[7], 
        DP_pipe0_coeff_pipe03[6], DP_pipe0_coeff_pipe03[5], 
        DP_pipe0_coeff_pipe03[4], DP_pipe0_coeff_pipe03[3], 
        DP_pipe0_coeff_pipe03[2], DP_pipe0_coeff_pipe03[1], 
        DP_pipe0_coeff_pipe03[0], SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154}) );
  INV_X1 U494 ( .A(n1091), .ZN(n1114) );
  INV_X1 U495 ( .A(n1091), .ZN(n1115) );
  INV_X1 U496 ( .A(n1091), .ZN(n1116) );
  INV_X1 U497 ( .A(n1091), .ZN(n1118) );
  INV_X1 U498 ( .A(n1092), .ZN(n1119) );
  INV_X1 U499 ( .A(n1092), .ZN(n1120) );
  INV_X1 U500 ( .A(n1092), .ZN(n1121) );
  INV_X1 U501 ( .A(n1041), .ZN(n1025) );
  INV_X1 U502 ( .A(n1042), .ZN(n1026) );
  BUF_X1 U503 ( .A(n1093), .Z(n1091) );
  BUF_X1 U504 ( .A(n1093), .Z(n1092) );
  BUF_X1 U505 ( .A(n1105), .Z(n1054) );
  BUF_X1 U506 ( .A(n1105), .Z(n1055) );
  BUF_X1 U507 ( .A(n1105), .Z(n1056) );
  BUF_X1 U508 ( .A(n1104), .Z(n1057) );
  BUF_X1 U509 ( .A(n1104), .Z(n1058) );
  BUF_X1 U510 ( .A(n1104), .Z(n1059) );
  BUF_X1 U511 ( .A(n1103), .Z(n1060) );
  BUF_X1 U512 ( .A(n1103), .Z(n1061) );
  BUF_X1 U513 ( .A(n1103), .Z(n1062) );
  BUF_X1 U514 ( .A(n1102), .Z(n1063) );
  BUF_X1 U515 ( .A(n1102), .Z(n1064) );
  BUF_X1 U516 ( .A(n1102), .Z(n1065) );
  BUF_X1 U517 ( .A(n1101), .Z(n1066) );
  BUF_X1 U518 ( .A(n1101), .Z(n1067) );
  BUF_X1 U519 ( .A(n1101), .Z(n1068) );
  BUF_X1 U520 ( .A(n1100), .Z(n1069) );
  BUF_X1 U521 ( .A(n1100), .Z(n1070) );
  BUF_X1 U522 ( .A(n1100), .Z(n1071) );
  BUF_X1 U523 ( .A(n1099), .Z(n1072) );
  BUF_X1 U524 ( .A(n1099), .Z(n1073) );
  BUF_X1 U525 ( .A(n1099), .Z(n1074) );
  BUF_X1 U526 ( .A(n1098), .Z(n1075) );
  BUF_X1 U527 ( .A(n1098), .Z(n1076) );
  BUF_X1 U528 ( .A(n1098), .Z(n1077) );
  BUF_X1 U529 ( .A(n1097), .Z(n1078) );
  BUF_X1 U530 ( .A(n1097), .Z(n1079) );
  BUF_X1 U531 ( .A(n1097), .Z(n1080) );
  BUF_X1 U532 ( .A(n1096), .Z(n1081) );
  BUF_X1 U533 ( .A(n1096), .Z(n1082) );
  BUF_X1 U534 ( .A(n1096), .Z(n1083) );
  BUF_X1 U535 ( .A(n1095), .Z(n1084) );
  BUF_X1 U536 ( .A(n1095), .Z(n1085) );
  BUF_X1 U537 ( .A(n1095), .Z(n1086) );
  BUF_X1 U538 ( .A(n1094), .Z(n1087) );
  BUF_X1 U539 ( .A(n1094), .Z(n1088) );
  BUF_X1 U540 ( .A(n1094), .Z(n1089) );
  BUF_X1 U541 ( .A(n1106), .Z(n1052) );
  BUF_X1 U542 ( .A(n1106), .Z(n1053) );
  BUF_X1 U543 ( .A(n1093), .Z(n1090) );
  BUF_X1 U544 ( .A(n1043), .Z(n1041) );
  BUF_X1 U545 ( .A(n1050), .Z(n1028) );
  BUF_X1 U546 ( .A(n1049), .Z(n1029) );
  BUF_X1 U547 ( .A(n1050), .Z(n1027) );
  BUF_X1 U548 ( .A(n1049), .Z(n1030) );
  BUF_X1 U549 ( .A(n1048), .Z(n1031) );
  BUF_X1 U550 ( .A(n1044), .Z(n1040) );
  BUF_X1 U551 ( .A(n1044), .Z(n1039) );
  BUF_X1 U552 ( .A(n1045), .Z(n1038) );
  BUF_X1 U553 ( .A(n1046), .Z(n1036) );
  BUF_X1 U554 ( .A(n1046), .Z(n1035) );
  BUF_X1 U555 ( .A(n1047), .Z(n1034) );
  BUF_X1 U556 ( .A(n1048), .Z(n1032) );
  BUF_X1 U557 ( .A(n1047), .Z(n1033) );
  BUF_X1 U558 ( .A(n1045), .Z(n1037) );
  BUF_X1 U559 ( .A(n1043), .Z(n1042) );
  BUF_X1 U560 ( .A(n1107), .Z(n1105) );
  BUF_X1 U561 ( .A(n1107), .Z(n1104) );
  BUF_X1 U562 ( .A(n1108), .Z(n1103) );
  BUF_X1 U563 ( .A(n1108), .Z(n1102) );
  BUF_X1 U564 ( .A(n1108), .Z(n1101) );
  BUF_X1 U565 ( .A(n1109), .Z(n1100) );
  BUF_X1 U566 ( .A(n1109), .Z(n1099) );
  BUF_X1 U567 ( .A(n1109), .Z(n1098) );
  BUF_X1 U568 ( .A(n1110), .Z(n1097) );
  BUF_X1 U569 ( .A(n1110), .Z(n1096) );
  BUF_X1 U570 ( .A(n1110), .Z(n1095) );
  BUF_X1 U571 ( .A(n1111), .Z(n1093) );
  BUF_X1 U572 ( .A(n1111), .Z(n1094) );
  BUF_X1 U573 ( .A(n1107), .Z(n1106) );
  BUF_X1 U574 ( .A(n1021), .Z(n1043) );
  BUF_X1 U575 ( .A(n1021), .Z(n1044) );
  BUF_X1 U576 ( .A(n1022), .Z(n1046) );
  BUF_X1 U577 ( .A(n1022), .Z(n1048) );
  BUF_X1 U578 ( .A(n1022), .Z(n1047) );
  BUF_X1 U579 ( .A(n1021), .Z(n1045) );
  BUF_X1 U580 ( .A(n1023), .Z(n1050) );
  BUF_X1 U581 ( .A(n1023), .Z(n1049) );
  NOR2_X1 U582 ( .A1(DP_y_23), .A2(DP_y_11_), .ZN(n1174) );
  NAND2_X1 U583 ( .A1(DP_y_23), .A2(DP_y_23), .ZN(n1170) );
  BUF_X1 U584 ( .A(n1112), .Z(n1109) );
  BUF_X1 U585 ( .A(n1112), .Z(n1110) );
  BUF_X1 U586 ( .A(n1113), .Z(n1107) );
  BUF_X1 U587 ( .A(n1113), .Z(n1108) );
  BUF_X1 U588 ( .A(n1112), .Z(n1111) );
  BUF_X1 U589 ( .A(n40), .Z(n1022) );
  BUF_X1 U590 ( .A(n40), .Z(n1021) );
  BUF_X1 U591 ( .A(n40), .Z(n1023) );
  NAND2_X1 U592 ( .A1(delayed_controls_2__0_), .A2(DP_N2), .ZN(n26) );
  OR2_X1 U593 ( .A1(n1020), .A2(DP_N4), .ZN(n24) );
  OAI221_X1 U594 ( .B1(n24), .B2(n25), .C1(delayed_controls_2__0_), .C2(n270), 
        .A(n26), .ZN(n513) );
  INV_X1 U595 ( .A(DP_y_0_), .ZN(n25) );
  OAI221_X1 U596 ( .B1(n24), .B2(n27), .C1(delayed_controls_2__0_), .C2(n271), 
        .A(n26), .ZN(n514) );
  INV_X1 U597 ( .A(DP_y_1_), .ZN(n27) );
  OAI221_X1 U598 ( .B1(n24), .B2(n28), .C1(delayed_controls_2__0_), .C2(n272), 
        .A(n26), .ZN(n515) );
  INV_X1 U599 ( .A(DP_y_2_), .ZN(n28) );
  OAI221_X1 U600 ( .B1(n24), .B2(n29), .C1(delayed_controls_2__0_), .C2(n273), 
        .A(n26), .ZN(n516) );
  INV_X1 U601 ( .A(DP_y_3_), .ZN(n29) );
  OAI221_X1 U602 ( .B1(n24), .B2(n30), .C1(delayed_controls_2__0_), .C2(n274), 
        .A(n26), .ZN(n517) );
  INV_X1 U603 ( .A(DP_y_4_), .ZN(n30) );
  OAI221_X1 U604 ( .B1(n24), .B2(n31), .C1(delayed_controls_2__0_), .C2(n275), 
        .A(n26), .ZN(n518) );
  INV_X1 U605 ( .A(DP_y_5_), .ZN(n31) );
  OAI221_X1 U606 ( .B1(n24), .B2(n32), .C1(delayed_controls_2__0_), .C2(n276), 
        .A(n26), .ZN(n519) );
  INV_X1 U607 ( .A(DP_y_6_), .ZN(n32) );
  OAI221_X1 U608 ( .B1(n24), .B2(n33), .C1(delayed_controls_2__0_), .C2(n277), 
        .A(n26), .ZN(n520) );
  INV_X1 U609 ( .A(DP_y_7_), .ZN(n33) );
  OAI221_X1 U610 ( .B1(n24), .B2(n34), .C1(delayed_controls_2__0_), .C2(n278), 
        .A(n26), .ZN(n521) );
  INV_X1 U611 ( .A(DP_y_8_), .ZN(n34) );
  OAI221_X1 U612 ( .B1(n24), .B2(n35), .C1(delayed_controls_2__0_), .C2(n279), 
        .A(n26), .ZN(n522) );
  INV_X1 U613 ( .A(DP_y_9_), .ZN(n35) );
  OAI221_X1 U614 ( .B1(n24), .B2(n36), .C1(delayed_controls_2__0_), .C2(n280), 
        .A(n26), .ZN(n523) );
  INV_X1 U615 ( .A(DP_y_10_), .ZN(n36) );
  OAI21_X1 U616 ( .B1(delayed_controls_2__0_), .B2(n281), .A(n38), .ZN(n524)
         );
  OAI211_X1 U617 ( .C1(DP_N4), .C2(DP_y_23), .A(n39), .B(
        delayed_controls_2__0_), .ZN(n38) );
  INV_X1 U618 ( .A(DP_N2), .ZN(n39) );
  INV_X1 U619 ( .A(DP_y_23), .ZN(n1173) );
  INV_X1 U620 ( .A(n107), .ZN(n661) );
  AOI22_X1 U621 ( .A1(n1025), .A2(DP_w_18_), .B1(n1032), .B2(DP_sw0_18_), .ZN(
        n107) );
  INV_X1 U622 ( .A(n108), .ZN(n663) );
  AOI22_X1 U623 ( .A1(n1025), .A2(DP_w_19_), .B1(n1032), .B2(DP_sw0_19_), .ZN(
        n108) );
  INV_X1 U624 ( .A(n111), .ZN(n669) );
  AOI22_X1 U625 ( .A1(n1025), .A2(DP_w_22_), .B1(n1033), .B2(DP_sw0_22_), .ZN(
        n111) );
  INV_X1 U626 ( .A(n109), .ZN(n665) );
  AOI22_X1 U627 ( .A1(n1025), .A2(DP_w_20_), .B1(n1032), .B2(DP_sw0_20_), .ZN(
        n109) );
  INV_X1 U628 ( .A(n103), .ZN(n653) );
  AOI22_X1 U629 ( .A1(n1025), .A2(DP_w_14_), .B1(n1033), .B2(DP_sw0_14_), .ZN(
        n103) );
  INV_X1 U630 ( .A(n104), .ZN(n655) );
  AOI22_X1 U631 ( .A1(n1025), .A2(DP_w_15_), .B1(n1033), .B2(DP_sw0_15_), .ZN(
        n104) );
  INV_X1 U632 ( .A(n105), .ZN(n657) );
  AOI22_X1 U633 ( .A1(n1025), .A2(DP_w_16_), .B1(n1032), .B2(DP_sw0_16_), .ZN(
        n105) );
  INV_X1 U634 ( .A(n106), .ZN(n659) );
  AOI22_X1 U635 ( .A1(n1025), .A2(DP_w_17_), .B1(n1032), .B2(DP_sw0_17_), .ZN(
        n106) );
  INV_X1 U636 ( .A(n110), .ZN(n667) );
  AOI22_X1 U637 ( .A1(n1025), .A2(DP_w_21_), .B1(n1031), .B2(DP_sw0_21_), .ZN(
        n110) );
  INV_X1 U638 ( .A(n112), .ZN(n671) );
  AOI22_X1 U639 ( .A1(n1026), .A2(DP_w_23_), .B1(n1037), .B2(DP_sw0_23_), .ZN(
        n112) );
  INV_X1 U640 ( .A(n135), .ZN(n861) );
  AOI22_X1 U641 ( .A1(DP_coeffs_ff_int[93]), .A2(n1115), .B1(coeffs_ff[2]), 
        .B2(n1057), .ZN(n135) );
  INV_X1 U642 ( .A(n159), .ZN(n885) );
  AOI22_X1 U643 ( .A1(DP_coeffs_ff_int[69]), .A2(n1119), .B1(coeffs_ff[26]), 
        .B2(n1062), .ZN(n159) );
  INV_X1 U644 ( .A(n183), .ZN(n909) );
  AOI22_X1 U645 ( .A1(DP_coeffs_ff_int[45]), .A2(n1118), .B1(coeffs_ff[50]), 
        .B2(n1068), .ZN(n183) );
  INV_X1 U646 ( .A(n207), .ZN(n933) );
  AOI22_X1 U647 ( .A1(DP_coeffs_ff_int[21]), .A2(n1120), .B1(coeffs_ff[74]), 
        .B2(n1075), .ZN(n207) );
  INV_X1 U648 ( .A(n231), .ZN(n957) );
  AOI22_X1 U649 ( .A1(DP_coeffs_fb_int[45]), .A2(n1119), .B1(coeffs_fb[2]), 
        .B2(n1081), .ZN(n231) );
  INV_X1 U650 ( .A(n255), .ZN(n981) );
  AOI22_X1 U651 ( .A1(DP_coeffs_fb_int[21]), .A2(n1118), .B1(coeffs_fb[26]), 
        .B2(n1087), .ZN(n255) );
  INV_X1 U652 ( .A(n93), .ZN(n633) );
  AOI22_X1 U653 ( .A1(n1025), .A2(DP_w_4_), .B1(n1035), .B2(DP_sw0_4_), .ZN(
        n93) );
  INV_X1 U654 ( .A(n94), .ZN(n635) );
  AOI22_X1 U655 ( .A1(n1026), .A2(DP_w_5_), .B1(n1035), .B2(DP_sw0_5_), .ZN(
        n94) );
  INV_X1 U656 ( .A(n95), .ZN(n637) );
  AOI22_X1 U657 ( .A1(n1025), .A2(DP_w_6_), .B1(n1035), .B2(DP_sw0_6_), .ZN(
        n95) );
  INV_X1 U658 ( .A(n96), .ZN(n639) );
  AOI22_X1 U659 ( .A1(n1025), .A2(DP_w_7_), .B1(n1034), .B2(DP_sw0_7_), .ZN(
        n96) );
  INV_X1 U660 ( .A(n97), .ZN(n641) );
  AOI22_X1 U661 ( .A1(n1026), .A2(DP_w_8_), .B1(n1034), .B2(DP_sw0_8_), .ZN(
        n97) );
  INV_X1 U662 ( .A(n98), .ZN(n643) );
  AOI22_X1 U663 ( .A1(n1024), .A2(DP_w_9_), .B1(n1034), .B2(DP_sw0_9_), .ZN(
        n98) );
  INV_X1 U664 ( .A(n99), .ZN(n645) );
  AOI22_X1 U665 ( .A1(n1025), .A2(DP_w_10_), .B1(n1034), .B2(DP_sw0_10_), .ZN(
        n99) );
  INV_X1 U666 ( .A(n100), .ZN(n647) );
  AOI22_X1 U667 ( .A1(n1026), .A2(DP_w_11_), .B1(n1034), .B2(DP_sw0_11_), .ZN(
        n100) );
  INV_X1 U668 ( .A(n101), .ZN(n649) );
  AOI22_X1 U669 ( .A1(n1025), .A2(DP_w_12_), .B1(n1033), .B2(DP_sw0_12_), .ZN(
        n101) );
  INV_X1 U670 ( .A(n102), .ZN(n651) );
  AOI22_X1 U671 ( .A1(n1025), .A2(DP_w_13_), .B1(n1033), .B2(DP_sw0_13_), .ZN(
        n102) );
  BUF_X1 U672 ( .A(vIn), .Z(n1112) );
  INV_X1 U673 ( .A(n162), .ZN(n888) );
  AOI22_X1 U674 ( .A1(DP_coeffs_ff_int[24]), .A2(n1117), .B1(coeffs_ff[71]), 
        .B2(n1063), .ZN(n162) );
  INV_X1 U675 ( .A(n163), .ZN(n889) );
  AOI22_X1 U676 ( .A1(DP_coeffs_ff_int[25]), .A2(n1117), .B1(coeffs_ff[70]), 
        .B2(n1063), .ZN(n163) );
  INV_X1 U677 ( .A(n164), .ZN(n890) );
  AOI22_X1 U678 ( .A1(DP_coeffs_ff_int[26]), .A2(n1117), .B1(coeffs_ff[69]), 
        .B2(n1064), .ZN(n164) );
  INV_X1 U679 ( .A(n165), .ZN(n891) );
  AOI22_X1 U680 ( .A1(DP_coeffs_ff_int[27]), .A2(n1117), .B1(coeffs_ff[68]), 
        .B2(n1064), .ZN(n165) );
  INV_X1 U681 ( .A(n166), .ZN(n892) );
  AOI22_X1 U682 ( .A1(DP_coeffs_ff_int[28]), .A2(n1117), .B1(coeffs_ff[67]), 
        .B2(n1064), .ZN(n166) );
  INV_X1 U683 ( .A(n167), .ZN(n893) );
  AOI22_X1 U684 ( .A1(DP_coeffs_ff_int[29]), .A2(n1117), .B1(coeffs_ff[66]), 
        .B2(n1064), .ZN(n167) );
  INV_X1 U685 ( .A(n168), .ZN(n894) );
  AOI22_X1 U686 ( .A1(DP_coeffs_ff_int[30]), .A2(n1117), .B1(coeffs_ff[65]), 
        .B2(n1065), .ZN(n168) );
  INV_X1 U687 ( .A(n169), .ZN(n895) );
  AOI22_X1 U688 ( .A1(DP_coeffs_ff_int[31]), .A2(n1117), .B1(coeffs_ff[64]), 
        .B2(n1065), .ZN(n169) );
  INV_X1 U689 ( .A(n170), .ZN(n896) );
  AOI22_X1 U690 ( .A1(DP_coeffs_ff_int[32]), .A2(n1117), .B1(coeffs_ff[63]), 
        .B2(n1065), .ZN(n170) );
  INV_X1 U691 ( .A(n171), .ZN(n897) );
  AOI22_X1 U692 ( .A1(DP_coeffs_ff_int[33]), .A2(n1117), .B1(coeffs_ff[62]), 
        .B2(n1065), .ZN(n171) );
  INV_X1 U693 ( .A(n172), .ZN(n898) );
  AOI22_X1 U694 ( .A1(DP_coeffs_ff_int[34]), .A2(n1117), .B1(coeffs_ff[61]), 
        .B2(n1066), .ZN(n172) );
  INV_X1 U695 ( .A(n173), .ZN(n899) );
  AOI22_X1 U696 ( .A1(DP_coeffs_ff_int[35]), .A2(n1117), .B1(coeffs_ff[60]), 
        .B2(n1066), .ZN(n173) );
  BUF_X1 U697 ( .A(vIn), .Z(n1113) );
  INV_X1 U698 ( .A(n113), .ZN(n840) );
  AOI22_X1 U699 ( .A1(DP_coeffs_ff_int[72]), .A2(n1114), .B1(n1090), .B2(
        coeffs_ff[23]), .ZN(n113) );
  INV_X1 U700 ( .A(n115), .ZN(n841) );
  AOI22_X1 U701 ( .A1(DP_coeffs_ff_int[73]), .A2(n1114), .B1(coeffs_ff[22]), 
        .B2(n1052), .ZN(n115) );
  INV_X1 U702 ( .A(n116), .ZN(n842) );
  AOI22_X1 U703 ( .A1(DP_coeffs_ff_int[74]), .A2(n1114), .B1(coeffs_ff[21]), 
        .B2(n1052), .ZN(n116) );
  INV_X1 U704 ( .A(n117), .ZN(n843) );
  AOI22_X1 U705 ( .A1(DP_coeffs_ff_int[75]), .A2(n1114), .B1(coeffs_ff[20]), 
        .B2(n1052), .ZN(n117) );
  INV_X1 U706 ( .A(n118), .ZN(n844) );
  AOI22_X1 U707 ( .A1(DP_coeffs_ff_int[76]), .A2(n1114), .B1(coeffs_ff[19]), 
        .B2(n1052), .ZN(n118) );
  INV_X1 U708 ( .A(n119), .ZN(n845) );
  AOI22_X1 U709 ( .A1(DP_coeffs_ff_int[77]), .A2(n1114), .B1(coeffs_ff[18]), 
        .B2(n1053), .ZN(n119) );
  INV_X1 U710 ( .A(n120), .ZN(n846) );
  AOI22_X1 U711 ( .A1(DP_coeffs_ff_int[78]), .A2(n1114), .B1(coeffs_ff[17]), 
        .B2(n1053), .ZN(n120) );
  INV_X1 U712 ( .A(n121), .ZN(n847) );
  AOI22_X1 U713 ( .A1(DP_coeffs_ff_int[79]), .A2(n1114), .B1(coeffs_ff[16]), 
        .B2(n1053), .ZN(n121) );
  INV_X1 U714 ( .A(n122), .ZN(n848) );
  AOI22_X1 U715 ( .A1(DP_coeffs_ff_int[80]), .A2(n1114), .B1(coeffs_ff[15]), 
        .B2(n1053), .ZN(n122) );
  INV_X1 U716 ( .A(n123), .ZN(n849) );
  AOI22_X1 U717 ( .A1(DP_coeffs_ff_int[81]), .A2(n1114), .B1(coeffs_ff[14]), 
        .B2(n1054), .ZN(n123) );
  INV_X1 U718 ( .A(n124), .ZN(n850) );
  AOI22_X1 U719 ( .A1(DP_coeffs_ff_int[82]), .A2(n1114), .B1(coeffs_ff[13]), 
        .B2(n1054), .ZN(n124) );
  INV_X1 U720 ( .A(n125), .ZN(n851) );
  AOI22_X1 U721 ( .A1(DP_coeffs_ff_int[83]), .A2(n1114), .B1(coeffs_ff[12]), 
        .B2(n1054), .ZN(n125) );
  INV_X1 U722 ( .A(n126), .ZN(n852) );
  AOI22_X1 U723 ( .A1(DP_coeffs_ff_int[84]), .A2(n1115), .B1(coeffs_ff[11]), 
        .B2(n1054), .ZN(n126) );
  INV_X1 U724 ( .A(n127), .ZN(n853) );
  AOI22_X1 U725 ( .A1(DP_coeffs_ff_int[85]), .A2(n1115), .B1(coeffs_ff[10]), 
        .B2(n1055), .ZN(n127) );
  INV_X1 U726 ( .A(n128), .ZN(n854) );
  AOI22_X1 U727 ( .A1(DP_coeffs_ff_int[86]), .A2(n1115), .B1(coeffs_ff[9]), 
        .B2(n1055), .ZN(n128) );
  INV_X1 U728 ( .A(n129), .ZN(n855) );
  AOI22_X1 U729 ( .A1(DP_coeffs_ff_int[87]), .A2(n1115), .B1(coeffs_ff[8]), 
        .B2(n1055), .ZN(n129) );
  INV_X1 U730 ( .A(n130), .ZN(n856) );
  AOI22_X1 U731 ( .A1(DP_coeffs_ff_int[88]), .A2(n1115), .B1(coeffs_ff[7]), 
        .B2(n1055), .ZN(n130) );
  INV_X1 U732 ( .A(n131), .ZN(n857) );
  AOI22_X1 U733 ( .A1(DP_coeffs_ff_int[89]), .A2(n1115), .B1(coeffs_ff[6]), 
        .B2(n1056), .ZN(n131) );
  INV_X1 U734 ( .A(n132), .ZN(n858) );
  AOI22_X1 U735 ( .A1(DP_coeffs_ff_int[90]), .A2(n1115), .B1(coeffs_ff[5]), 
        .B2(n1056), .ZN(n132) );
  INV_X1 U736 ( .A(n133), .ZN(n859) );
  AOI22_X1 U737 ( .A1(DP_coeffs_ff_int[91]), .A2(n1115), .B1(coeffs_ff[4]), 
        .B2(n1056), .ZN(n133) );
  INV_X1 U738 ( .A(n134), .ZN(n860) );
  AOI22_X1 U739 ( .A1(DP_coeffs_ff_int[92]), .A2(n1115), .B1(coeffs_ff[3]), 
        .B2(n1056), .ZN(n134) );
  INV_X1 U740 ( .A(n136), .ZN(n862) );
  AOI22_X1 U741 ( .A1(DP_coeffs_ff_int[94]), .A2(n1115), .B1(coeffs_ff[1]), 
        .B2(n1057), .ZN(n136) );
  INV_X1 U742 ( .A(n137), .ZN(n863) );
  AOI22_X1 U743 ( .A1(DP_coeffs_ff_int[95]), .A2(n1115), .B1(coeffs_ff[0]), 
        .B2(n1057), .ZN(n137) );
  INV_X1 U744 ( .A(n138), .ZN(n864) );
  AOI22_X1 U745 ( .A1(DP_coeffs_ff_int[48]), .A2(n1116), .B1(coeffs_ff[47]), 
        .B2(n1057), .ZN(n138) );
  INV_X1 U746 ( .A(n139), .ZN(n865) );
  AOI22_X1 U747 ( .A1(DP_coeffs_ff_int[49]), .A2(n1116), .B1(coeffs_ff[46]), 
        .B2(n1058), .ZN(n139) );
  INV_X1 U748 ( .A(n140), .ZN(n866) );
  AOI22_X1 U749 ( .A1(DP_coeffs_ff_int[50]), .A2(n1116), .B1(coeffs_ff[45]), 
        .B2(n1058), .ZN(n140) );
  INV_X1 U750 ( .A(n141), .ZN(n867) );
  AOI22_X1 U751 ( .A1(DP_coeffs_ff_int[51]), .A2(n1116), .B1(coeffs_ff[44]), 
        .B2(n1058), .ZN(n141) );
  INV_X1 U752 ( .A(n142), .ZN(n868) );
  AOI22_X1 U753 ( .A1(DP_coeffs_ff_int[52]), .A2(n1116), .B1(coeffs_ff[43]), 
        .B2(n1058), .ZN(n142) );
  INV_X1 U754 ( .A(n143), .ZN(n869) );
  AOI22_X1 U755 ( .A1(DP_coeffs_ff_int[53]), .A2(n1116), .B1(coeffs_ff[42]), 
        .B2(n1071), .ZN(n143) );
  INV_X1 U756 ( .A(n144), .ZN(n870) );
  AOI22_X1 U757 ( .A1(DP_coeffs_ff_int[54]), .A2(n1116), .B1(coeffs_ff[41]), 
        .B2(n1059), .ZN(n144) );
  INV_X1 U758 ( .A(n145), .ZN(n871) );
  AOI22_X1 U759 ( .A1(DP_coeffs_ff_int[55]), .A2(n1116), .B1(coeffs_ff[40]), 
        .B2(n1059), .ZN(n145) );
  INV_X1 U760 ( .A(n146), .ZN(n872) );
  AOI22_X1 U761 ( .A1(DP_coeffs_ff_int[56]), .A2(n1116), .B1(coeffs_ff[39]), 
        .B2(n1059), .ZN(n146) );
  INV_X1 U762 ( .A(n147), .ZN(n873) );
  AOI22_X1 U763 ( .A1(DP_coeffs_ff_int[57]), .A2(n1116), .B1(coeffs_ff[38]), 
        .B2(n1059), .ZN(n147) );
  INV_X1 U764 ( .A(n148), .ZN(n874) );
  AOI22_X1 U765 ( .A1(DP_coeffs_ff_int[58]), .A2(n1116), .B1(coeffs_ff[37]), 
        .B2(n1060), .ZN(n148) );
  INV_X1 U766 ( .A(n149), .ZN(n875) );
  AOI22_X1 U767 ( .A1(DP_coeffs_ff_int[59]), .A2(n1116), .B1(coeffs_ff[36]), 
        .B2(n1060), .ZN(n149) );
  INV_X1 U768 ( .A(n150), .ZN(n876) );
  AOI22_X1 U769 ( .A1(DP_coeffs_ff_int[60]), .A2(n1118), .B1(coeffs_ff[35]), 
        .B2(n1060), .ZN(n150) );
  INV_X1 U770 ( .A(n151), .ZN(n877) );
  AOI22_X1 U771 ( .A1(DP_coeffs_ff_int[61]), .A2(n1115), .B1(coeffs_ff[34]), 
        .B2(n1060), .ZN(n151) );
  INV_X1 U772 ( .A(n152), .ZN(n878) );
  AOI22_X1 U773 ( .A1(DP_coeffs_ff_int[62]), .A2(n1117), .B1(coeffs_ff[33]), 
        .B2(n1061), .ZN(n152) );
  INV_X1 U774 ( .A(n153), .ZN(n879) );
  AOI22_X1 U775 ( .A1(DP_coeffs_ff_int[63]), .A2(n1120), .B1(coeffs_ff[32]), 
        .B2(n1061), .ZN(n153) );
  INV_X1 U776 ( .A(n154), .ZN(n880) );
  AOI22_X1 U777 ( .A1(DP_coeffs_ff_int[64]), .A2(n1116), .B1(coeffs_ff[31]), 
        .B2(n1061), .ZN(n154) );
  INV_X1 U778 ( .A(n155), .ZN(n881) );
  AOI22_X1 U779 ( .A1(DP_coeffs_ff_int[65]), .A2(n1114), .B1(coeffs_ff[30]), 
        .B2(n1061), .ZN(n155) );
  INV_X1 U780 ( .A(n156), .ZN(n882) );
  AOI22_X1 U781 ( .A1(DP_coeffs_ff_int[66]), .A2(n1114), .B1(coeffs_ff[29]), 
        .B2(n1062), .ZN(n156) );
  INV_X1 U782 ( .A(n157), .ZN(n883) );
  AOI22_X1 U783 ( .A1(DP_coeffs_ff_int[67]), .A2(n1120), .B1(coeffs_ff[28]), 
        .B2(n1062), .ZN(n157) );
  INV_X1 U784 ( .A(n158), .ZN(n884) );
  AOI22_X1 U785 ( .A1(DP_coeffs_ff_int[68]), .A2(n1117), .B1(coeffs_ff[27]), 
        .B2(n1062), .ZN(n158) );
  INV_X1 U786 ( .A(n160), .ZN(n886) );
  AOI22_X1 U787 ( .A1(DP_coeffs_ff_int[70]), .A2(n1115), .B1(coeffs_ff[25]), 
        .B2(n1063), .ZN(n160) );
  INV_X1 U788 ( .A(n161), .ZN(n887) );
  AOI22_X1 U789 ( .A1(DP_coeffs_ff_int[71]), .A2(n1117), .B1(coeffs_ff[24]), 
        .B2(n1063), .ZN(n161) );
  INV_X1 U790 ( .A(n174), .ZN(n900) );
  AOI22_X1 U791 ( .A1(DP_coeffs_ff_int[36]), .A2(n1118), .B1(coeffs_ff[59]), 
        .B2(n1066), .ZN(n174) );
  INV_X1 U792 ( .A(n175), .ZN(n901) );
  AOI22_X1 U793 ( .A1(DP_coeffs_ff_int[37]), .A2(n1118), .B1(coeffs_ff[58]), 
        .B2(n1066), .ZN(n175) );
  INV_X1 U794 ( .A(n176), .ZN(n902) );
  AOI22_X1 U795 ( .A1(DP_coeffs_ff_int[38]), .A2(n1118), .B1(coeffs_ff[57]), 
        .B2(n1067), .ZN(n176) );
  INV_X1 U796 ( .A(n177), .ZN(n903) );
  AOI22_X1 U797 ( .A1(DP_coeffs_ff_int[39]), .A2(n1118), .B1(coeffs_ff[56]), 
        .B2(n1067), .ZN(n177) );
  INV_X1 U798 ( .A(n178), .ZN(n904) );
  AOI22_X1 U799 ( .A1(DP_coeffs_ff_int[40]), .A2(n1118), .B1(coeffs_ff[55]), 
        .B2(n1067), .ZN(n178) );
  INV_X1 U800 ( .A(n179), .ZN(n905) );
  AOI22_X1 U801 ( .A1(DP_coeffs_ff_int[41]), .A2(n1118), .B1(coeffs_ff[54]), 
        .B2(n1067), .ZN(n179) );
  INV_X1 U802 ( .A(n180), .ZN(n906) );
  AOI22_X1 U803 ( .A1(DP_coeffs_ff_int[42]), .A2(n1118), .B1(coeffs_ff[53]), 
        .B2(n1068), .ZN(n180) );
  INV_X1 U804 ( .A(n181), .ZN(n907) );
  AOI22_X1 U805 ( .A1(DP_coeffs_ff_int[43]), .A2(n1118), .B1(coeffs_ff[52]), 
        .B2(n1068), .ZN(n181) );
  INV_X1 U806 ( .A(n182), .ZN(n908) );
  AOI22_X1 U807 ( .A1(DP_coeffs_ff_int[44]), .A2(n1118), .B1(coeffs_ff[51]), 
        .B2(n1068), .ZN(n182) );
  INV_X1 U808 ( .A(n184), .ZN(n910) );
  AOI22_X1 U809 ( .A1(DP_coeffs_ff_int[46]), .A2(n1118), .B1(coeffs_ff[49]), 
        .B2(n1069), .ZN(n184) );
  INV_X1 U810 ( .A(n185), .ZN(n911) );
  AOI22_X1 U811 ( .A1(DP_coeffs_ff_int[47]), .A2(n1118), .B1(coeffs_ff[48]), 
        .B2(n1069), .ZN(n185) );
  INV_X1 U812 ( .A(n258), .ZN(n984) );
  AOI22_X1 U813 ( .A1(DP_x[11]), .A2(n1118), .B1(dIn[11]), .B2(n1088), .ZN(
        n258) );
  INV_X1 U814 ( .A(n259), .ZN(n985) );
  AOI22_X1 U815 ( .A1(DP_x[10]), .A2(n1120), .B1(dIn[10]), .B2(n1087), .ZN(
        n259) );
  INV_X1 U816 ( .A(n260), .ZN(n986) );
  AOI22_X1 U817 ( .A1(DP_x[9]), .A2(n1119), .B1(dIn[9]), .B2(n1088), .ZN(n260)
         );
  INV_X1 U818 ( .A(n261), .ZN(n987) );
  AOI22_X1 U819 ( .A1(DP_x[8]), .A2(n1120), .B1(dIn[8]), .B2(n1088), .ZN(n261)
         );
  INV_X1 U820 ( .A(n262), .ZN(n988) );
  AOI22_X1 U821 ( .A1(DP_x[7]), .A2(n1115), .B1(dIn[7]), .B2(n1088), .ZN(n262)
         );
  INV_X1 U822 ( .A(n263), .ZN(n989) );
  AOI22_X1 U823 ( .A1(DP_x[6]), .A2(n1117), .B1(dIn[6]), .B2(n1089), .ZN(n263)
         );
  INV_X1 U824 ( .A(n264), .ZN(n990) );
  AOI22_X1 U825 ( .A1(DP_x[5]), .A2(n1117), .B1(dIn[5]), .B2(n1089), .ZN(n264)
         );
  INV_X1 U826 ( .A(n265), .ZN(n991) );
  AOI22_X1 U827 ( .A1(DP_x[4]), .A2(n1121), .B1(dIn[4]), .B2(n1089), .ZN(n265)
         );
  INV_X1 U828 ( .A(n266), .ZN(n992) );
  AOI22_X1 U829 ( .A1(DP_x[3]), .A2(n1116), .B1(dIn[3]), .B2(n1090), .ZN(n266)
         );
  INV_X1 U830 ( .A(n267), .ZN(n993) );
  AOI22_X1 U831 ( .A1(DP_x[2]), .A2(n1114), .B1(dIn[2]), .B2(n1090), .ZN(n267)
         );
  INV_X1 U832 ( .A(n268), .ZN(n994) );
  AOI22_X1 U833 ( .A1(DP_x[1]), .A2(n1121), .B1(dIn[1]), .B2(n1089), .ZN(n268)
         );
  INV_X1 U834 ( .A(n269), .ZN(n995) );
  AOI22_X1 U835 ( .A1(DP_x[0]), .A2(n1118), .B1(dIn[0]), .B2(n1090), .ZN(n269)
         );
  INV_X1 U836 ( .A(n186), .ZN(n912) );
  AOI22_X1 U837 ( .A1(DP_coeffs_ff_int[0]), .A2(n1119), .B1(coeffs_ff[95]), 
        .B2(n1069), .ZN(n186) );
  INV_X1 U838 ( .A(n187), .ZN(n913) );
  AOI22_X1 U839 ( .A1(DP_coeffs_ff_int[1]), .A2(n1119), .B1(coeffs_ff[94]), 
        .B2(n1069), .ZN(n187) );
  INV_X1 U840 ( .A(n188), .ZN(n914) );
  AOI22_X1 U841 ( .A1(DP_coeffs_ff_int[2]), .A2(n1119), .B1(coeffs_ff[93]), 
        .B2(n1070), .ZN(n188) );
  INV_X1 U842 ( .A(n189), .ZN(n915) );
  AOI22_X1 U843 ( .A1(DP_coeffs_ff_int[3]), .A2(n1119), .B1(coeffs_ff[92]), 
        .B2(n1070), .ZN(n189) );
  INV_X1 U844 ( .A(n190), .ZN(n916) );
  AOI22_X1 U845 ( .A1(DP_coeffs_ff_int[4]), .A2(n1119), .B1(coeffs_ff[91]), 
        .B2(n1070), .ZN(n190) );
  INV_X1 U846 ( .A(n191), .ZN(n917) );
  AOI22_X1 U847 ( .A1(DP_coeffs_ff_int[5]), .A2(n1119), .B1(coeffs_ff[90]), 
        .B2(n1070), .ZN(n191) );
  INV_X1 U848 ( .A(n192), .ZN(n918) );
  AOI22_X1 U849 ( .A1(DP_coeffs_ff_int[6]), .A2(n1119), .B1(coeffs_ff[89]), 
        .B2(n1071), .ZN(n192) );
  INV_X1 U850 ( .A(n193), .ZN(n919) );
  AOI22_X1 U851 ( .A1(DP_coeffs_ff_int[7]), .A2(n1119), .B1(coeffs_ff[88]), 
        .B2(n1071), .ZN(n193) );
  INV_X1 U852 ( .A(n194), .ZN(n920) );
  AOI22_X1 U853 ( .A1(DP_coeffs_ff_int[8]), .A2(n1119), .B1(coeffs_ff[87]), 
        .B2(n1071), .ZN(n194) );
  INV_X1 U854 ( .A(n195), .ZN(n921) );
  AOI22_X1 U855 ( .A1(DP_coeffs_ff_int[9]), .A2(n1119), .B1(coeffs_ff[86]), 
        .B2(n1072), .ZN(n195) );
  INV_X1 U856 ( .A(n196), .ZN(n922) );
  AOI22_X1 U857 ( .A1(DP_coeffs_ff_int[10]), .A2(n1119), .B1(coeffs_ff[85]), 
        .B2(n1072), .ZN(n196) );
  INV_X1 U858 ( .A(n197), .ZN(n923) );
  AOI22_X1 U859 ( .A1(DP_coeffs_ff_int[11]), .A2(n1119), .B1(coeffs_ff[84]), 
        .B2(n1072), .ZN(n197) );
  INV_X1 U860 ( .A(n198), .ZN(n924) );
  AOI22_X1 U861 ( .A1(DP_coeffs_ff_int[12]), .A2(n1120), .B1(coeffs_ff[83]), 
        .B2(n1072), .ZN(n198) );
  INV_X1 U862 ( .A(n199), .ZN(n925) );
  AOI22_X1 U863 ( .A1(DP_coeffs_ff_int[13]), .A2(n1120), .B1(coeffs_ff[82]), 
        .B2(n1073), .ZN(n199) );
  INV_X1 U864 ( .A(n200), .ZN(n926) );
  AOI22_X1 U865 ( .A1(DP_coeffs_ff_int[14]), .A2(n1120), .B1(coeffs_ff[81]), 
        .B2(n1073), .ZN(n200) );
  INV_X1 U866 ( .A(n201), .ZN(n927) );
  AOI22_X1 U867 ( .A1(DP_coeffs_ff_int[15]), .A2(n1120), .B1(coeffs_ff[80]), 
        .B2(n1073), .ZN(n201) );
  INV_X1 U868 ( .A(n202), .ZN(n928) );
  AOI22_X1 U869 ( .A1(DP_coeffs_ff_int[16]), .A2(n1120), .B1(coeffs_ff[79]), 
        .B2(n1073), .ZN(n202) );
  INV_X1 U870 ( .A(n203), .ZN(n929) );
  AOI22_X1 U871 ( .A1(DP_coeffs_ff_int[17]), .A2(n1120), .B1(coeffs_ff[78]), 
        .B2(n1074), .ZN(n203) );
  INV_X1 U872 ( .A(n204), .ZN(n930) );
  AOI22_X1 U873 ( .A1(DP_coeffs_ff_int[18]), .A2(n1120), .B1(coeffs_ff[77]), 
        .B2(n1074), .ZN(n204) );
  INV_X1 U874 ( .A(n205), .ZN(n931) );
  AOI22_X1 U875 ( .A1(DP_coeffs_ff_int[19]), .A2(n1120), .B1(coeffs_ff[76]), 
        .B2(n1074), .ZN(n205) );
  INV_X1 U876 ( .A(n206), .ZN(n932) );
  AOI22_X1 U877 ( .A1(DP_coeffs_ff_int[20]), .A2(n1120), .B1(coeffs_ff[75]), 
        .B2(n1074), .ZN(n206) );
  INV_X1 U878 ( .A(n208), .ZN(n934) );
  AOI22_X1 U879 ( .A1(DP_coeffs_ff_int[22]), .A2(n1120), .B1(coeffs_ff[73]), 
        .B2(n1075), .ZN(n208) );
  INV_X1 U880 ( .A(n209), .ZN(n935) );
  AOI22_X1 U881 ( .A1(DP_coeffs_ff_int[23]), .A2(n1120), .B1(coeffs_ff[72]), 
        .B2(n1075), .ZN(n209) );
  INV_X1 U882 ( .A(n210), .ZN(n936) );
  AOI22_X1 U883 ( .A1(DP_coeffs_fb_int[24]), .A2(n1121), .B1(coeffs_fb[23]), 
        .B2(n1075), .ZN(n210) );
  INV_X1 U884 ( .A(n211), .ZN(n937) );
  AOI22_X1 U885 ( .A1(DP_coeffs_fb_int[25]), .A2(n1121), .B1(coeffs_fb[22]), 
        .B2(n1076), .ZN(n211) );
  INV_X1 U886 ( .A(n212), .ZN(n938) );
  AOI22_X1 U887 ( .A1(DP_coeffs_fb_int[26]), .A2(n1121), .B1(coeffs_fb[21]), 
        .B2(n1076), .ZN(n212) );
  INV_X1 U888 ( .A(n213), .ZN(n939) );
  AOI22_X1 U889 ( .A1(DP_coeffs_fb_int[27]), .A2(n1121), .B1(coeffs_fb[20]), 
        .B2(n1076), .ZN(n213) );
  INV_X1 U890 ( .A(n214), .ZN(n940) );
  AOI22_X1 U891 ( .A1(DP_coeffs_fb_int[28]), .A2(n1121), .B1(coeffs_fb[19]), 
        .B2(n1076), .ZN(n214) );
  INV_X1 U892 ( .A(n215), .ZN(n941) );
  AOI22_X1 U893 ( .A1(DP_coeffs_fb_int[29]), .A2(n1121), .B1(coeffs_fb[18]), 
        .B2(n1077), .ZN(n215) );
  INV_X1 U894 ( .A(n216), .ZN(n942) );
  AOI22_X1 U895 ( .A1(DP_coeffs_fb_int[30]), .A2(n1121), .B1(coeffs_fb[17]), 
        .B2(n1077), .ZN(n216) );
  INV_X1 U896 ( .A(n217), .ZN(n943) );
  AOI22_X1 U897 ( .A1(DP_coeffs_fb_int[31]), .A2(n1121), .B1(coeffs_fb[16]), 
        .B2(n1077), .ZN(n217) );
  INV_X1 U898 ( .A(n218), .ZN(n944) );
  AOI22_X1 U899 ( .A1(DP_coeffs_fb_int[32]), .A2(n1121), .B1(coeffs_fb[15]), 
        .B2(n1077), .ZN(n218) );
  INV_X1 U900 ( .A(n219), .ZN(n945) );
  AOI22_X1 U901 ( .A1(DP_coeffs_fb_int[33]), .A2(n1121), .B1(coeffs_fb[14]), 
        .B2(n1078), .ZN(n219) );
  INV_X1 U902 ( .A(n220), .ZN(n946) );
  AOI22_X1 U903 ( .A1(DP_coeffs_fb_int[34]), .A2(n1121), .B1(coeffs_fb[13]), 
        .B2(n1078), .ZN(n220) );
  INV_X1 U904 ( .A(n221), .ZN(n947) );
  AOI22_X1 U905 ( .A1(DP_coeffs_fb_int[35]), .A2(n1121), .B1(coeffs_fb[12]), 
        .B2(n1078), .ZN(n221) );
  INV_X1 U906 ( .A(n222), .ZN(n948) );
  AOI22_X1 U907 ( .A1(DP_coeffs_fb_int[36]), .A2(n1116), .B1(coeffs_fb[11]), 
        .B2(n1078), .ZN(n222) );
  INV_X1 U908 ( .A(n223), .ZN(n949) );
  AOI22_X1 U909 ( .A1(DP_coeffs_fb_int[37]), .A2(n1119), .B1(coeffs_fb[10]), 
        .B2(n1079), .ZN(n223) );
  INV_X1 U910 ( .A(n224), .ZN(n950) );
  AOI22_X1 U911 ( .A1(DP_coeffs_fb_int[38]), .A2(n1118), .B1(coeffs_fb[9]), 
        .B2(n1079), .ZN(n224) );
  INV_X1 U912 ( .A(n225), .ZN(n951) );
  AOI22_X1 U913 ( .A1(DP_coeffs_fb_int[39]), .A2(n1114), .B1(coeffs_fb[8]), 
        .B2(n1079), .ZN(n225) );
  INV_X1 U914 ( .A(n226), .ZN(n952) );
  AOI22_X1 U915 ( .A1(DP_coeffs_fb_int[40]), .A2(n1115), .B1(coeffs_fb[7]), 
        .B2(n1079), .ZN(n226) );
  INV_X1 U916 ( .A(n227), .ZN(n953) );
  AOI22_X1 U917 ( .A1(DP_coeffs_fb_int[41]), .A2(n1117), .B1(coeffs_fb[6]), 
        .B2(n1080), .ZN(n227) );
  INV_X1 U918 ( .A(n228), .ZN(n954) );
  AOI22_X1 U919 ( .A1(DP_coeffs_fb_int[42]), .A2(n1121), .B1(coeffs_fb[5]), 
        .B2(n1080), .ZN(n228) );
  INV_X1 U920 ( .A(n229), .ZN(n955) );
  AOI22_X1 U921 ( .A1(DP_coeffs_fb_int[43]), .A2(n1118), .B1(coeffs_fb[4]), 
        .B2(n1080), .ZN(n229) );
  INV_X1 U922 ( .A(n230), .ZN(n956) );
  AOI22_X1 U923 ( .A1(DP_coeffs_fb_int[44]), .A2(n1116), .B1(coeffs_fb[3]), 
        .B2(n1080), .ZN(n230) );
  INV_X1 U924 ( .A(n232), .ZN(n958) );
  AOI22_X1 U925 ( .A1(DP_coeffs_fb_int[46]), .A2(n1120), .B1(coeffs_fb[1]), 
        .B2(n1081), .ZN(n232) );
  INV_X1 U926 ( .A(n233), .ZN(n959) );
  AOI22_X1 U927 ( .A1(DP_coeffs_fb_int[47]), .A2(n1119), .B1(coeffs_fb[0]), 
        .B2(n1081), .ZN(n233) );
  INV_X1 U928 ( .A(n234), .ZN(n960) );
  AOI22_X1 U929 ( .A1(DP_coeffs_fb_int[0]), .A2(n1115), .B1(coeffs_fb[47]), 
        .B2(n1081), .ZN(n234) );
  INV_X1 U930 ( .A(n235), .ZN(n961) );
  AOI22_X1 U931 ( .A1(DP_coeffs_fb_int[1]), .A2(n1115), .B1(coeffs_fb[46]), 
        .B2(n1082), .ZN(n235) );
  INV_X1 U932 ( .A(n236), .ZN(n962) );
  AOI22_X1 U933 ( .A1(DP_coeffs_fb_int[2]), .A2(n1118), .B1(coeffs_fb[45]), 
        .B2(n1082), .ZN(n236) );
  INV_X1 U934 ( .A(n237), .ZN(n963) );
  AOI22_X1 U935 ( .A1(DP_coeffs_fb_int[3]), .A2(n1117), .B1(coeffs_fb[44]), 
        .B2(n1082), .ZN(n237) );
  INV_X1 U936 ( .A(n238), .ZN(n964) );
  AOI22_X1 U937 ( .A1(DP_coeffs_fb_int[4]), .A2(n1121), .B1(coeffs_fb[43]), 
        .B2(n1082), .ZN(n238) );
  INV_X1 U938 ( .A(n239), .ZN(n965) );
  AOI22_X1 U939 ( .A1(DP_coeffs_fb_int[5]), .A2(n1114), .B1(coeffs_fb[42]), 
        .B2(n1083), .ZN(n239) );
  INV_X1 U940 ( .A(n240), .ZN(n966) );
  AOI22_X1 U941 ( .A1(DP_coeffs_fb_int[6]), .A2(n1119), .B1(coeffs_fb[41]), 
        .B2(n1083), .ZN(n240) );
  INV_X1 U942 ( .A(n241), .ZN(n967) );
  AOI22_X1 U943 ( .A1(DP_coeffs_fb_int[7]), .A2(n1116), .B1(coeffs_fb[40]), 
        .B2(n1083), .ZN(n241) );
  INV_X1 U944 ( .A(n242), .ZN(n968) );
  AOI22_X1 U945 ( .A1(DP_coeffs_fb_int[8]), .A2(n1120), .B1(coeffs_fb[39]), 
        .B2(n1084), .ZN(n242) );
  INV_X1 U946 ( .A(n243), .ZN(n969) );
  AOI22_X1 U947 ( .A1(DP_coeffs_fb_int[9]), .A2(n1116), .B1(coeffs_fb[38]), 
        .B2(n1084), .ZN(n243) );
  INV_X1 U948 ( .A(n244), .ZN(n970) );
  AOI22_X1 U949 ( .A1(DP_coeffs_fb_int[10]), .A2(n1121), .B1(coeffs_fb[37]), 
        .B2(n1083), .ZN(n244) );
  INV_X1 U950 ( .A(n245), .ZN(n971) );
  AOI22_X1 U951 ( .A1(DP_coeffs_fb_int[11]), .A2(n1114), .B1(coeffs_fb[36]), 
        .B2(n1084), .ZN(n245) );
  INV_X1 U952 ( .A(n246), .ZN(n972) );
  AOI22_X1 U953 ( .A1(DP_coeffs_fb_int[12]), .A2(n1119), .B1(coeffs_fb[35]), 
        .B2(n1085), .ZN(n246) );
  INV_X1 U954 ( .A(n247), .ZN(n973) );
  AOI22_X1 U955 ( .A1(DP_coeffs_fb_int[13]), .A2(n1116), .B1(coeffs_fb[34]), 
        .B2(n1084), .ZN(n247) );
  INV_X1 U956 ( .A(n248), .ZN(n974) );
  AOI22_X1 U957 ( .A1(DP_coeffs_fb_int[14]), .A2(n1115), .B1(coeffs_fb[33]), 
        .B2(n1085), .ZN(n248) );
  INV_X1 U958 ( .A(n249), .ZN(n975) );
  AOI22_X1 U959 ( .A1(DP_coeffs_fb_int[15]), .A2(n1114), .B1(coeffs_fb[32]), 
        .B2(n1085), .ZN(n249) );
  INV_X1 U960 ( .A(n250), .ZN(n976) );
  AOI22_X1 U961 ( .A1(DP_coeffs_fb_int[16]), .A2(n1120), .B1(coeffs_fb[31]), 
        .B2(n1085), .ZN(n250) );
  INV_X1 U962 ( .A(n251), .ZN(n977) );
  AOI22_X1 U963 ( .A1(DP_coeffs_fb_int[17]), .A2(n1121), .B1(coeffs_fb[30]), 
        .B2(n1086), .ZN(n251) );
  INV_X1 U964 ( .A(n252), .ZN(n978) );
  AOI22_X1 U965 ( .A1(DP_coeffs_fb_int[18]), .A2(n1117), .B1(coeffs_fb[29]), 
        .B2(n1086), .ZN(n252) );
  INV_X1 U966 ( .A(n253), .ZN(n979) );
  AOI22_X1 U967 ( .A1(DP_coeffs_fb_int[19]), .A2(n1120), .B1(coeffs_fb[28]), 
        .B2(n1086), .ZN(n253) );
  INV_X1 U968 ( .A(n254), .ZN(n980) );
  AOI22_X1 U969 ( .A1(DP_coeffs_fb_int[20]), .A2(n1121), .B1(coeffs_fb[27]), 
        .B2(n1087), .ZN(n254) );
  INV_X1 U970 ( .A(n256), .ZN(n982) );
  AOI22_X1 U971 ( .A1(DP_coeffs_fb_int[22]), .A2(n1119), .B1(coeffs_fb[25]), 
        .B2(n1086), .ZN(n256) );
  INV_X1 U972 ( .A(n257), .ZN(n983) );
  AOI22_X1 U973 ( .A1(DP_coeffs_fb_int[23]), .A2(n1121), .B1(coeffs_fb[24]), 
        .B2(n1087), .ZN(n257) );
  INV_X1 U974 ( .A(n87), .ZN(n621) );
  AOI22_X1 U975 ( .A1(n1026), .A2(DP_sw0_22_), .B1(n1036), .B2(DP_sw1_22_), 
        .ZN(n87) );
  OAI22_X1 U976 ( .A1(n1027), .A2(n1019), .B1(n1024), .B2(n284), .ZN(n529) );
  OAI22_X1 U977 ( .A1(n1027), .A2(n1017), .B1(n1024), .B2(n285), .ZN(n531) );
  OAI22_X1 U978 ( .A1(n1028), .A2(n1016), .B1(n1024), .B2(n286), .ZN(n533) );
  OAI22_X1 U979 ( .A1(n1027), .A2(n998), .B1(n1024), .B2(n287), .ZN(n535) );
  OAI22_X1 U980 ( .A1(n1028), .A2(n999), .B1(n1024), .B2(n288), .ZN(n537) );
  OAI22_X1 U981 ( .A1(n1028), .A2(n1000), .B1(n1024), .B2(n289), .ZN(n539) );
  OAI22_X1 U982 ( .A1(n1028), .A2(n1001), .B1(n1024), .B2(n290), .ZN(n541) );
  OAI22_X1 U983 ( .A1(n1028), .A2(n1002), .B1(n1024), .B2(n291), .ZN(n543) );
  OAI22_X1 U984 ( .A1(n1029), .A2(n1003), .B1(n1024), .B2(n292), .ZN(n545) );
  OAI22_X1 U985 ( .A1(n1029), .A2(n1004), .B1(n1024), .B2(n293), .ZN(n547) );
  OAI22_X1 U986 ( .A1(n1029), .A2(n1005), .B1(n1024), .B2(n294), .ZN(n549) );
  OAI22_X1 U987 ( .A1(n1029), .A2(n1006), .B1(n1024), .B2(n295), .ZN(n551) );
  OAI22_X1 U988 ( .A1(n1030), .A2(n1007), .B1(n1025), .B2(n296), .ZN(n553) );
  OAI22_X1 U989 ( .A1(n1027), .A2(n1008), .B1(n1024), .B2(n297), .ZN(n555) );
  OAI22_X1 U990 ( .A1(n1030), .A2(n1009), .B1(n1024), .B2(n298), .ZN(n557) );
  OAI22_X1 U991 ( .A1(n1029), .A2(n1010), .B1(n1026), .B2(n299), .ZN(n559) );
  OAI22_X1 U992 ( .A1(n1030), .A2(n1011), .B1(n1024), .B2(n300), .ZN(n561) );
  OAI22_X1 U993 ( .A1(n1031), .A2(n1012), .B1(n1025), .B2(n301), .ZN(n563) );
  OAI22_X1 U994 ( .A1(n1031), .A2(n1013), .B1(n1026), .B2(n302), .ZN(n565) );
  OAI22_X1 U995 ( .A1(n1030), .A2(n1014), .B1(n1024), .B2(n303), .ZN(n567) );
  OAI22_X1 U996 ( .A1(n1031), .A2(n997), .B1(n1024), .B2(n304), .ZN(n569) );
  OAI22_X1 U997 ( .A1(n1027), .A2(n1018), .B1(n1024), .B2(n305), .ZN(n571) );
  OAI22_X1 U998 ( .A1(n1031), .A2(n1015), .B1(n1024), .B2(n306), .ZN(n573) );
  OAI22_X1 U999 ( .A1(n1030), .A2(n996), .B1(n1025), .B2(n307), .ZN(n575) );
  INV_X1 U1000 ( .A(n92), .ZN(n631) );
  AOI22_X1 U1001 ( .A1(n1024), .A2(DP_w_3_), .B1(n1035), .B2(DP_sw0_3_), .ZN(
        n92) );
  INV_X1 U1002 ( .A(n85), .ZN(n617) );
  AOI22_X1 U1003 ( .A1(n1025), .A2(DP_sw0_20_), .B1(n1037), .B2(DP_sw1_20_), 
        .ZN(n85) );
  INV_X1 U1004 ( .A(n68), .ZN(n583) );
  AOI22_X1 U1005 ( .A1(n1026), .A2(DP_sw0_3_), .B1(n1040), .B2(DP_sw1_3_), 
        .ZN(n68) );
  INV_X1 U1006 ( .A(n69), .ZN(n585) );
  AOI22_X1 U1007 ( .A1(n1026), .A2(DP_sw0_4_), .B1(n1040), .B2(DP_sw1_4_), 
        .ZN(n69) );
  INV_X1 U1008 ( .A(n70), .ZN(n587) );
  AOI22_X1 U1009 ( .A1(n1026), .A2(DP_sw0_5_), .B1(n1040), .B2(DP_sw1_5_), 
        .ZN(n70) );
  INV_X1 U1010 ( .A(n71), .ZN(n589) );
  AOI22_X1 U1011 ( .A1(n1026), .A2(DP_sw0_6_), .B1(n1040), .B2(DP_sw1_6_), 
        .ZN(n71) );
  INV_X1 U1012 ( .A(n72), .ZN(n591) );
  AOI22_X1 U1013 ( .A1(n1026), .A2(DP_sw0_7_), .B1(n1039), .B2(DP_sw1_7_), 
        .ZN(n72) );
  INV_X1 U1014 ( .A(n73), .ZN(n593) );
  AOI22_X1 U1015 ( .A1(n1026), .A2(DP_sw0_8_), .B1(n1039), .B2(DP_sw1_8_), 
        .ZN(n73) );
  INV_X1 U1016 ( .A(n74), .ZN(n595) );
  AOI22_X1 U1017 ( .A1(n1026), .A2(DP_sw0_9_), .B1(n1039), .B2(DP_sw1_9_), 
        .ZN(n74) );
  INV_X1 U1018 ( .A(n75), .ZN(n597) );
  AOI22_X1 U1019 ( .A1(n1026), .A2(DP_sw0_10_), .B1(n1039), .B2(DP_sw1_10_), 
        .ZN(n75) );
  INV_X1 U1020 ( .A(n76), .ZN(n599) );
  AOI22_X1 U1021 ( .A1(n1025), .A2(DP_sw0_11_), .B1(n1039), .B2(DP_sw1_11_), 
        .ZN(n76) );
  INV_X1 U1022 ( .A(n77), .ZN(n601) );
  AOI22_X1 U1023 ( .A1(n1024), .A2(DP_sw0_12_), .B1(n1038), .B2(DP_sw1_12_), 
        .ZN(n77) );
  INV_X1 U1024 ( .A(n78), .ZN(n603) );
  AOI22_X1 U1025 ( .A1(n1025), .A2(DP_sw0_13_), .B1(n1038), .B2(DP_sw1_13_), 
        .ZN(n78) );
  INV_X1 U1026 ( .A(n79), .ZN(n605) );
  AOI22_X1 U1027 ( .A1(n1026), .A2(DP_sw0_14_), .B1(n1038), .B2(DP_sw1_14_), 
        .ZN(n79) );
  INV_X1 U1028 ( .A(n80), .ZN(n607) );
  AOI22_X1 U1029 ( .A1(n1024), .A2(DP_sw0_15_), .B1(n1038), .B2(DP_sw1_15_), 
        .ZN(n80) );
  INV_X1 U1030 ( .A(n81), .ZN(n609) );
  AOI22_X1 U1031 ( .A1(n1024), .A2(DP_sw0_16_), .B1(n1038), .B2(DP_sw1_16_), 
        .ZN(n81) );
  INV_X1 U1032 ( .A(n82), .ZN(n611) );
  AOI22_X1 U1033 ( .A1(n1025), .A2(DP_sw0_17_), .B1(n1037), .B2(DP_sw1_17_), 
        .ZN(n82) );
  INV_X1 U1034 ( .A(n83), .ZN(n613) );
  AOI22_X1 U1035 ( .A1(n1025), .A2(DP_sw0_18_), .B1(n1037), .B2(DP_sw1_18_), 
        .ZN(n83) );
  INV_X1 U1036 ( .A(n84), .ZN(n615) );
  AOI22_X1 U1037 ( .A1(n1026), .A2(DP_sw0_19_), .B1(n1037), .B2(DP_sw1_19_), 
        .ZN(n84) );
  INV_X1 U1038 ( .A(n91), .ZN(n629) );
  AOI22_X1 U1039 ( .A1(n1026), .A2(DP_w_2_), .B1(n1035), .B2(DP_sw0_2_), .ZN(
        n91) );
  INV_X1 U1040 ( .A(n67), .ZN(n581) );
  AOI22_X1 U1041 ( .A1(n1026), .A2(DP_sw0_2_), .B1(n1040), .B2(DP_sw1_2_), 
        .ZN(n67) );
  INV_X1 U1042 ( .A(n90), .ZN(n627) );
  AOI22_X1 U1043 ( .A1(n1024), .A2(DP_w_1_), .B1(n1036), .B2(DP_sw0_1_), .ZN(
        n90) );
  INV_X1 U1044 ( .A(n66), .ZN(n579) );
  AOI22_X1 U1045 ( .A1(n1026), .A2(DP_sw0_1_), .B1(n1041), .B2(DP_sw1_1_), 
        .ZN(n66) );
  INV_X1 U1046 ( .A(n86), .ZN(n619) );
  AOI22_X1 U1047 ( .A1(n1025), .A2(DP_sw0_21_), .B1(n1036), .B2(DP_sw1_21_), 
        .ZN(n86) );
  INV_X1 U1048 ( .A(n89), .ZN(n625) );
  AOI22_X1 U1049 ( .A1(n1025), .A2(DP_w_0_), .B1(n1036), .B2(DP_sw0_0_), .ZN(
        n89) );
  INV_X1 U1050 ( .A(n65), .ZN(n577) );
  AOI22_X1 U1051 ( .A1(n1026), .A2(DP_sw0_0_), .B1(n1041), .B2(DP_sw1_0_), 
        .ZN(n65) );
  INV_X1 U1052 ( .A(n88), .ZN(n623) );
  AOI22_X1 U1053 ( .A1(n1026), .A2(DP_sw0_23_), .B1(n1036), .B2(n1051), .ZN(
        n88) );
  BUF_X1 U1054 ( .A(rst_n), .Z(n1163) );
  BUF_X1 U1055 ( .A(rst_n), .Z(n1164) );
  BUF_X1 U1056 ( .A(rst_n), .Z(n1165) );
  BUF_X1 U1057 ( .A(rst_n), .Z(n1166) );
  BUF_X1 U1058 ( .A(rst_n), .Z(n1167) );
  BUF_X1 U1059 ( .A(rst_n), .Z(n1168) );
  BUF_X1 U1060 ( .A(rst_n), .Z(n1169) );
  NAND3_X1 U1061 ( .A1(DP_y_23), .A2(DP_y_11_), .A3(DP_y_23), .ZN(n1171) );
  INV_X1 U1062 ( .A(n1041), .ZN(n1024) );
  INV_X1 U1063 ( .A(n996), .ZN(n1051) );
  INV_X1 U1064 ( .A(n1092), .ZN(n1117) );
  CLKBUF_X1 U1065 ( .A(n1169), .Z(n1122) );
  CLKBUF_X1 U1066 ( .A(n1169), .Z(n1123) );
  CLKBUF_X1 U1067 ( .A(n1169), .Z(n1124) );
  CLKBUF_X1 U1068 ( .A(n1169), .Z(n1125) );
  CLKBUF_X1 U1069 ( .A(n1169), .Z(n1126) );
  CLKBUF_X1 U1070 ( .A(n1168), .Z(n1127) );
  CLKBUF_X1 U1071 ( .A(n1168), .Z(n1128) );
  CLKBUF_X1 U1072 ( .A(n1168), .Z(n1129) );
  CLKBUF_X1 U1073 ( .A(n1168), .Z(n1130) );
  CLKBUF_X1 U1074 ( .A(n1168), .Z(n1131) );
  CLKBUF_X1 U1075 ( .A(n1168), .Z(n1132) );
  CLKBUF_X1 U1076 ( .A(n1167), .Z(n1133) );
  CLKBUF_X1 U1077 ( .A(n1167), .Z(n1134) );
  CLKBUF_X1 U1078 ( .A(n1167), .Z(n1135) );
  CLKBUF_X1 U1079 ( .A(n1167), .Z(n1136) );
  CLKBUF_X1 U1080 ( .A(n1167), .Z(n1137) );
  CLKBUF_X1 U1081 ( .A(n1167), .Z(n1138) );
  CLKBUF_X1 U1082 ( .A(n1166), .Z(n1139) );
  CLKBUF_X1 U1083 ( .A(n1166), .Z(n1140) );
  CLKBUF_X1 U1084 ( .A(n1166), .Z(n1141) );
  CLKBUF_X1 U1085 ( .A(n1166), .Z(n1142) );
  CLKBUF_X1 U1086 ( .A(n1166), .Z(n1143) );
  CLKBUF_X1 U1087 ( .A(n1166), .Z(n1144) );
  CLKBUF_X1 U1088 ( .A(n1165), .Z(n1145) );
  CLKBUF_X1 U1089 ( .A(n1165), .Z(n1146) );
  CLKBUF_X1 U1090 ( .A(n1165), .Z(n1147) );
  CLKBUF_X1 U1091 ( .A(n1165), .Z(n1148) );
  CLKBUF_X1 U1092 ( .A(n1165), .Z(n1149) );
  CLKBUF_X1 U1093 ( .A(n1165), .Z(n1150) );
  CLKBUF_X1 U1094 ( .A(n1164), .Z(n1151) );
  CLKBUF_X1 U1095 ( .A(n1164), .Z(n1152) );
  CLKBUF_X1 U1096 ( .A(n1164), .Z(n1153) );
  CLKBUF_X1 U1097 ( .A(n1164), .Z(n1154) );
  CLKBUF_X1 U1098 ( .A(n1164), .Z(n1155) );
  CLKBUF_X1 U1099 ( .A(n1164), .Z(n1156) );
  CLKBUF_X1 U1100 ( .A(n1163), .Z(n1157) );
  CLKBUF_X1 U1101 ( .A(n1163), .Z(n1158) );
  CLKBUF_X1 U1102 ( .A(n1163), .Z(n1159) );
  CLKBUF_X1 U1103 ( .A(n1163), .Z(n1160) );
  CLKBUF_X1 U1104 ( .A(n1163), .Z(n1161) );
  CLKBUF_X1 U1105 ( .A(n1163), .Z(n1162) );
  NOR2_X1 U1106 ( .A1(n1171), .A2(n1170), .ZN(n1172) );
  OAI22_X1 U1107 ( .A1(n1172), .A2(n1173), .B1(DP_y_23), .B2(n1173), .ZN(DP_N4) );
  AND2_X1 U1108 ( .A1(n1174), .A2(n1173), .ZN(n1175) );
  OAI22_X1 U1109 ( .A1(DP_y_23), .A2(n1175), .B1(DP_y_23), .B2(n1173), .ZN(
        DP_N2) );
endmodule

