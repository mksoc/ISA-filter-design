
module iir_filter ( clk, rst_n, vIn, dIn, a, b, dOut, vOut );
  input [11:0] dIn;
  input [23:0] a;
  input [35:0] b;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   regs_clr_int, reg_sw0_en_int, DP_n35, DP_n34, DP_n33, DP_n32, DP_n31,
         DP_n30, DP_n29, DP_n28, DP_n27, DP_n26, DP_n25, DP_n24, DP_n23,
         DP_n22, DP_n21, DP_n20, DP_n19, DP_n18, DP_n17, DP_n16, DP_n15,
         DP_n14, DP_n13, DP_n12, DP_n11, DP_n10, DP_n9, DP_n8, DP_n7, DP_n6,
         DP_n5, DP_n4, DP_n3, DP_n2, DP_n1, DP_fb_0_, DP_fb_10_, DP_fb_11_,
         DP_fb_12_, DP_fb_1_, DP_fb_2_, DP_fb_3_, DP_fb_4_, DP_fb_5_, DP_fb_6_,
         DP_fb_7_, DP_fb_8_, DP_fb_9_, DP_ff_0_, DP_ff_10_, DP_ff_11_,
         DP_ff_12_, DP_ff_1_, DP_ff_2_, DP_ff_3_, DP_ff_4_, DP_ff_5_, DP_ff_6_,
         DP_ff_7_, DP_ff_8_, DP_ff_9_, DP_y_0_, DP_y_1_, DP_y_2_, DP_y_3_,
         DP_y_4_, DP_y_5_, DP_y_6_, DP_y_7_, DP_y_8_, DP_y_9_, DP_y_10_,
         DP_y_11_, DP_w_b0_0_, DP_w_b0_1_, DP_w_b0_2_, DP_w_b0_3_, DP_w_b0_4_,
         DP_w_b0_5_, DP_w_b0_6_, DP_w_b0_7_, DP_w_b0_8_, DP_w_b0_9_,
         DP_w_b0_10_, DP_w_b0_11_, DP_sw1_b2_0_, DP_sw1_b2_1_, DP_sw1_b2_2_,
         DP_sw1_b2_3_, DP_sw1_b2_4_, DP_sw1_b2_5_, DP_sw1_b2_6_, DP_sw1_b2_7_,
         DP_sw1_b2_8_, DP_sw1_b2_9_, DP_sw1_b2_10_, DP_sw1_b2_11_,
         DP_sw0_b1_0_, DP_sw0_b1_1_, DP_sw0_b1_2_, DP_sw0_b1_3_, DP_sw0_b1_4_,
         DP_sw0_b1_5_, DP_sw0_b1_6_, DP_sw0_b1_7_, DP_sw0_b1_8_, DP_sw0_b1_9_,
         DP_sw0_b1_10_, DP_sw0_b1_11_, DP_sw1_a2_0_, DP_sw1_a2_1_,
         DP_sw1_a2_2_, DP_sw1_a2_3_, DP_sw1_a2_4_, DP_sw1_a2_5_, DP_sw1_a2_6_,
         DP_sw1_a2_7_, DP_sw1_a2_8_, DP_sw1_a2_9_, DP_sw1_a2_10_,
         DP_sw1_a2_11_, DP_sw0_a1_0_, DP_sw0_a1_1_, DP_sw0_a1_2_, DP_sw0_a1_3_,
         DP_sw0_a1_4_, DP_sw0_a1_5_, DP_sw0_a1_6_, DP_sw0_a1_7_, DP_sw0_a1_8_,
         DP_sw0_a1_9_, DP_sw0_a1_10_, DP_sw0_a1_11_, DP_y_out_0_, DP_y_out_1_,
         DP_y_out_2_, DP_y_out_3_, DP_y_out_4_, DP_y_out_5_, DP_y_out_6_,
         DP_y_out_7_, DP_y_out_8_, DP_y_out_9_, DP_y_out_10_, DP_y_out_11_,
         DP_sw1_0_, DP_sw1_1_, DP_sw1_2_, DP_sw1_3_, DP_sw1_4_, DP_sw1_5_,
         DP_sw1_6_, DP_sw1_7_, DP_sw1_8_, DP_sw1_9_, DP_sw1_10_, DP_sw1_11_,
         DP_sw1_12_, DP_sw0_0_, DP_sw0_1_, DP_sw0_2_, DP_sw0_3_, DP_sw0_4_,
         DP_sw0_5_, DP_sw0_6_, DP_sw0_7_, DP_sw0_8_, DP_sw0_9_, DP_sw0_10_,
         DP_sw0_11_, DP_sw0_12_, DP_w_0_, DP_w_1_, DP_w_2_, DP_w_3_, DP_w_4_,
         DP_w_5_, DP_w_6_, DP_w_7_, DP_w_8_, DP_w_9_, DP_w_10_, DP_w_11_,
         DP_w_12_, DP_x_0_, DP_x_1_, DP_x_2_, DP_x_3_, DP_x_4_, DP_x_5_,
         DP_x_6_, DP_x_7_, DP_x_8_, DP_x_9_, DP_x_10_, DP_x_11_, DP_reg_in_n39,
         DP_reg_in_n38, DP_reg_in_n37, DP_reg_in_n36, DP_reg_in_n35,
         DP_reg_in_n34, DP_reg_in_n33, DP_reg_in_n32, DP_reg_in_n31,
         DP_reg_in_n30, DP_reg_in_n29, DP_reg_in_n28, DP_reg_in_n27,
         DP_reg_in_n26, DP_reg_in_n25, DP_reg_in_n24, DP_reg_in_n23,
         DP_reg_in_n22, DP_reg_in_n21, DP_reg_in_n20, DP_reg_in_n19,
         DP_reg_in_n18, DP_reg_in_n17, DP_reg_in_n16, DP_reg_in_n15,
         DP_reg_in_n14, DP_reg_in_n13, DP_reg_in_n12, DP_reg_in_n11,
         DP_reg_in_n10, DP_reg_in_n9, DP_reg_in_n8, DP_reg_in_n7, DP_reg_in_n6,
         DP_reg_in_n5, DP_reg_in_n4, DP_reg_in_n3, DP_reg_in_n2, DP_reg_in_n1,
         DP_reg_a_i_1_n76, DP_reg_a_i_1_n75, DP_reg_a_i_1_n74,
         DP_reg_a_i_1_n73, DP_reg_a_i_1_n72, DP_reg_a_i_1_n71,
         DP_reg_a_i_1_n70, DP_reg_a_i_1_n69, DP_reg_a_i_1_n68,
         DP_reg_a_i_1_n67, DP_reg_a_i_1_n66, DP_reg_a_i_1_n65,
         DP_reg_a_i_1_n64, DP_reg_a_i_1_n63, DP_reg_a_i_1_n62,
         DP_reg_a_i_1_n61, DP_reg_a_i_1_n60, DP_reg_a_i_1_n59,
         DP_reg_a_i_1_n58, DP_reg_a_i_1_n57, DP_reg_a_i_1_n56,
         DP_reg_a_i_1_n55, DP_reg_a_i_1_n54, DP_reg_a_i_1_n53,
         DP_reg_a_i_1_n52, DP_reg_a_i_1_n51, DP_reg_a_i_1_n50,
         DP_reg_a_i_1_n49, DP_reg_a_i_1_n48, DP_reg_a_i_1_n47,
         DP_reg_a_i_1_n46, DP_reg_a_i_1_n45, DP_reg_a_i_1_n44,
         DP_reg_a_i_1_n43, DP_reg_a_i_1_n42, DP_reg_a_i_1_n41,
         DP_reg_a_i_1_n40, DP_reg_a_i_1_n39, DP_reg_a_i_1_n38,
         DP_reg_a_i_2_n92, DP_reg_a_i_2_n91, DP_reg_a_i_2_n90,
         DP_reg_a_i_2_n89, DP_reg_a_i_2_n88, DP_reg_a_i_2_n87,
         DP_reg_a_i_2_n86, DP_reg_a_i_2_n85, DP_reg_a_i_2_n84,
         DP_reg_a_i_2_n83, DP_reg_a_i_2_n82, DP_reg_a_i_2_n81,
         DP_reg_a_i_2_n80, DP_reg_a_i_2_n79, DP_reg_a_i_2_n78,
         DP_reg_a_i_2_n77, DP_reg_a_i_2_n76, DP_reg_a_i_2_n75,
         DP_reg_a_i_2_n74, DP_reg_a_i_2_n73, DP_reg_a_i_2_n72,
         DP_reg_a_i_2_n71, DP_reg_a_i_2_n70, DP_reg_a_i_2_n69,
         DP_reg_a_i_2_n68, DP_reg_a_i_2_n67, DP_reg_a_i_2_n66,
         DP_reg_a_i_2_n65, DP_reg_a_i_2_n64, DP_reg_a_i_2_n63,
         DP_reg_a_i_2_n62, DP_reg_a_i_2_n61, DP_reg_a_i_2_n60,
         DP_reg_a_i_2_n59, DP_reg_a_i_2_n58, DP_reg_a_i_2_n57,
         DP_reg_a_i_2_n56, DP_reg_a_i_2_n55, DP_reg_a_i_2_n54,
         DP_reg_b_i_0_n76, DP_reg_b_i_0_n75, DP_reg_b_i_0_n74,
         DP_reg_b_i_0_n73, DP_reg_b_i_0_n72, DP_reg_b_i_0_n71,
         DP_reg_b_i_0_n70, DP_reg_b_i_0_n69, DP_reg_b_i_0_n68,
         DP_reg_b_i_0_n67, DP_reg_b_i_0_n66, DP_reg_b_i_0_n65,
         DP_reg_b_i_0_n64, DP_reg_b_i_0_n63, DP_reg_b_i_0_n62,
         DP_reg_b_i_0_n61, DP_reg_b_i_0_n60, DP_reg_b_i_0_n59,
         DP_reg_b_i_0_n58, DP_reg_b_i_0_n57, DP_reg_b_i_0_n56,
         DP_reg_b_i_0_n55, DP_reg_b_i_0_n54, DP_reg_b_i_0_n53,
         DP_reg_b_i_0_n52, DP_reg_b_i_0_n51, DP_reg_b_i_0_n50,
         DP_reg_b_i_0_n49, DP_reg_b_i_0_n48, DP_reg_b_i_0_n47,
         DP_reg_b_i_0_n46, DP_reg_b_i_0_n45, DP_reg_b_i_0_n44,
         DP_reg_b_i_0_n43, DP_reg_b_i_0_n42, DP_reg_b_i_0_n41,
         DP_reg_b_i_0_n40, DP_reg_b_i_0_n39, DP_reg_b_i_0_n38,
         DP_reg_b_i_1_n76, DP_reg_b_i_1_n75, DP_reg_b_i_1_n74,
         DP_reg_b_i_1_n73, DP_reg_b_i_1_n72, DP_reg_b_i_1_n71,
         DP_reg_b_i_1_n70, DP_reg_b_i_1_n69, DP_reg_b_i_1_n68,
         DP_reg_b_i_1_n67, DP_reg_b_i_1_n66, DP_reg_b_i_1_n65,
         DP_reg_b_i_1_n64, DP_reg_b_i_1_n63, DP_reg_b_i_1_n62,
         DP_reg_b_i_1_n61, DP_reg_b_i_1_n60, DP_reg_b_i_1_n59,
         DP_reg_b_i_1_n58, DP_reg_b_i_1_n57, DP_reg_b_i_1_n56,
         DP_reg_b_i_1_n55, DP_reg_b_i_1_n54, DP_reg_b_i_1_n53,
         DP_reg_b_i_1_n52, DP_reg_b_i_1_n51, DP_reg_b_i_1_n50,
         DP_reg_b_i_1_n49, DP_reg_b_i_1_n48, DP_reg_b_i_1_n47,
         DP_reg_b_i_1_n46, DP_reg_b_i_1_n45, DP_reg_b_i_1_n44,
         DP_reg_b_i_1_n43, DP_reg_b_i_1_n42, DP_reg_b_i_1_n41,
         DP_reg_b_i_1_n40, DP_reg_b_i_1_n39, DP_reg_b_i_1_n38,
         DP_reg_b_i_2_n76, DP_reg_b_i_2_n75, DP_reg_b_i_2_n74,
         DP_reg_b_i_2_n73, DP_reg_b_i_2_n72, DP_reg_b_i_2_n71,
         DP_reg_b_i_2_n70, DP_reg_b_i_2_n69, DP_reg_b_i_2_n68,
         DP_reg_b_i_2_n67, DP_reg_b_i_2_n66, DP_reg_b_i_2_n65,
         DP_reg_b_i_2_n64, DP_reg_b_i_2_n63, DP_reg_b_i_2_n62,
         DP_reg_b_i_2_n61, DP_reg_b_i_2_n60, DP_reg_b_i_2_n59,
         DP_reg_b_i_2_n58, DP_reg_b_i_2_n57, DP_reg_b_i_2_n56,
         DP_reg_b_i_2_n55, DP_reg_b_i_2_n54, DP_reg_b_i_2_n53,
         DP_reg_b_i_2_n52, DP_reg_b_i_2_n51, DP_reg_b_i_2_n50,
         DP_reg_b_i_2_n49, DP_reg_b_i_2_n48, DP_reg_b_i_2_n47,
         DP_reg_b_i_2_n46, DP_reg_b_i_2_n45, DP_reg_b_i_2_n44,
         DP_reg_b_i_2_n43, DP_reg_b_i_2_n42, DP_reg_b_i_2_n41,
         DP_reg_b_i_2_n40, DP_reg_b_i_2_n39, DP_reg_b_i_2_n38, DP_reg_sw0_n47,
         DP_reg_sw0_n46, DP_reg_sw0_n40, DP_reg_sw0_n39, DP_reg_sw0_n38,
         DP_reg_sw0_n37, DP_reg_sw0_n36, DP_reg_sw0_n35, DP_reg_sw0_n34,
         DP_reg_sw0_n33, DP_reg_sw0_n32, DP_reg_sw0_n31, DP_reg_sw0_n30,
         DP_reg_sw0_n29, DP_reg_sw0_n28, DP_reg_sw0_n27, DP_reg_sw0_n26,
         DP_reg_sw0_n25, DP_reg_sw0_n24, DP_reg_sw0_n23, DP_reg_sw0_n22,
         DP_reg_sw0_n21, DP_reg_sw0_n20, DP_reg_sw0_n19, DP_reg_sw0_n18,
         DP_reg_sw0_n17, DP_reg_sw0_n16, DP_reg_sw0_n15, DP_reg_sw0_n14,
         DP_reg_sw0_n13, DP_reg_sw0_n12, DP_reg_sw0_n11, DP_reg_sw0_n10,
         DP_reg_sw0_n9, DP_reg_sw0_n8, DP_reg_sw0_n7, DP_reg_sw0_n6,
         DP_reg_sw0_n5, DP_reg_sw0_n4, DP_reg_sw0_n3, DP_reg_sw0_n2,
         DP_reg_sw0_n1, DP_reg_sw1_n92, DP_reg_sw1_n91, DP_reg_sw1_n90,
         DP_reg_sw1_n89, DP_reg_sw1_n88, DP_reg_sw1_n87, DP_reg_sw1_n86,
         DP_reg_sw1_n85, DP_reg_sw1_n84, DP_reg_sw1_n83, DP_reg_sw1_n82,
         DP_reg_sw1_n81, DP_reg_sw1_n80, DP_reg_sw1_n79, DP_reg_sw1_n78,
         DP_reg_sw1_n77, DP_reg_sw1_n76, DP_reg_sw1_n75, DP_reg_sw1_n74,
         DP_reg_sw1_n73, DP_reg_sw1_n72, DP_reg_sw1_n71, DP_reg_sw1_n70,
         DP_reg_sw1_n69, DP_reg_sw1_n68, DP_reg_sw1_n67, DP_reg_sw1_n66,
         DP_reg_sw1_n65, DP_reg_sw1_n64, DP_reg_sw1_n63, DP_reg_sw1_n62,
         DP_reg_sw1_n61, DP_reg_sw1_n60, DP_reg_sw1_n59, DP_reg_sw1_n58,
         DP_reg_sw1_n57, DP_reg_sw1_n56, DP_reg_sw1_n55, DP_reg_sw1_n54,
         DP_reg_sw1_n53, DP_reg_sw1_n52, DP_reg_sw1_n48, DP_reg_sw1_n47,
         DP_reg_sw1_n46, DP_reg_sw1_n45, DP_reg_sw1_n41, DP_reg_out_n44,
         DP_reg_out_n43, DP_reg_out_n42, DP_reg_out_n41, DP_reg_out_n40,
         DP_reg_out_n39, DP_reg_out_n38, DP_reg_out_n37, DP_reg_out_n36,
         DP_reg_out_n35, DP_reg_out_n24, DP_reg_out_n23, DP_reg_out_n22,
         DP_reg_out_n9, DP_add_1_root_add_0_root_add_107_carry_1_,
         DP_add_1_root_add_0_root_add_107_carry_2_,
         DP_add_1_root_add_0_root_add_107_carry_3_,
         DP_add_1_root_add_0_root_add_107_carry_4_,
         DP_add_1_root_add_0_root_add_107_carry_5_,
         DP_add_1_root_add_0_root_add_107_carry_6_,
         DP_add_1_root_add_0_root_add_107_carry_7_,
         DP_add_1_root_add_0_root_add_107_carry_8_,
         DP_add_1_root_add_0_root_add_107_carry_9_,
         DP_add_1_root_add_0_root_add_107_carry_10_,
         DP_add_1_root_add_0_root_add_107_carry_11_,
         DP_add_1_root_add_0_root_add_107_carry_12_,
         DP_add_0_root_add_0_root_add_107_n82,
         DP_add_0_root_add_0_root_add_107_n81,
         DP_add_0_root_add_0_root_add_107_n80,
         DP_add_0_root_add_0_root_add_107_n79,
         DP_add_0_root_add_0_root_add_107_n78,
         DP_add_0_root_add_0_root_add_107_n77,
         DP_add_0_root_add_0_root_add_107_n76,
         DP_add_0_root_add_0_root_add_107_n75,
         DP_add_0_root_add_0_root_add_107_n74,
         DP_add_0_root_add_0_root_add_107_n73,
         DP_add_0_root_add_0_root_add_107_n72,
         DP_add_0_root_add_0_root_add_107_n71,
         DP_add_0_root_add_0_root_add_107_n70,
         DP_add_0_root_add_0_root_add_107_n69,
         DP_add_0_root_add_0_root_add_107_n68,
         DP_add_0_root_add_0_root_add_107_n67,
         DP_add_0_root_add_0_root_add_107_n66,
         DP_add_0_root_add_0_root_add_107_n65,
         DP_add_0_root_add_0_root_add_107_n64,
         DP_add_0_root_add_0_root_add_107_n63,
         DP_add_0_root_add_0_root_add_107_n62,
         DP_add_0_root_add_0_root_add_107_n61,
         DP_add_0_root_add_0_root_add_107_n60,
         DP_add_0_root_add_0_root_add_107_n59,
         DP_add_0_root_add_0_root_add_107_n58,
         DP_add_0_root_add_0_root_add_107_n57,
         DP_add_0_root_add_0_root_add_107_n56,
         DP_add_0_root_add_0_root_add_107_n55,
         DP_add_0_root_add_0_root_add_107_n54,
         DP_add_0_root_add_0_root_add_107_n53,
         DP_add_0_root_add_0_root_add_107_n52,
         DP_add_0_root_add_0_root_add_107_n51,
         DP_add_0_root_add_0_root_add_107_n50,
         DP_add_0_root_add_0_root_add_107_n49,
         DP_add_0_root_add_0_root_add_107_n48,
         DP_add_0_root_add_0_root_add_107_n47,
         DP_add_0_root_add_0_root_add_107_n46,
         DP_add_0_root_add_0_root_add_107_n45,
         DP_add_0_root_add_0_root_add_107_n44,
         DP_add_0_root_add_0_root_add_107_n43,
         DP_add_0_root_add_0_root_add_107_n42,
         DP_add_0_root_add_0_root_add_107_n41,
         DP_add_0_root_add_0_root_add_107_n40,
         DP_add_0_root_add_0_root_add_107_n39,
         DP_add_0_root_add_0_root_add_107_n38,
         DP_add_0_root_add_0_root_add_107_n37,
         DP_add_0_root_add_0_root_add_107_n36,
         DP_add_0_root_add_0_root_add_107_n35,
         DP_add_0_root_add_0_root_add_107_n34,
         DP_add_0_root_add_0_root_add_107_n33,
         DP_add_0_root_add_0_root_add_107_n32,
         DP_add_0_root_add_0_root_add_107_n31,
         DP_add_0_root_add_0_root_add_107_n30,
         DP_add_0_root_add_0_root_add_107_n29,
         DP_add_0_root_add_0_root_add_107_n28,
         DP_add_0_root_add_0_root_add_107_n27,
         DP_add_0_root_add_0_root_add_107_n26,
         DP_add_0_root_add_0_root_add_107_n25,
         DP_add_0_root_add_0_root_add_107_n24,
         DP_add_0_root_add_0_root_add_107_n23,
         DP_add_0_root_add_0_root_add_107_n22,
         DP_add_0_root_add_0_root_add_107_n21,
         DP_add_0_root_add_0_root_add_107_n20,
         DP_add_0_root_add_0_root_add_107_n19,
         DP_add_0_root_add_0_root_add_107_n18,
         DP_add_0_root_add_0_root_add_107_n17,
         DP_add_0_root_add_0_root_add_107_n16,
         DP_add_0_root_add_0_root_add_107_n15,
         DP_add_0_root_add_0_root_add_107_n14,
         DP_add_0_root_add_0_root_add_107_n13,
         DP_add_0_root_add_0_root_add_107_n12,
         DP_add_0_root_add_0_root_add_107_n11,
         DP_add_0_root_add_0_root_add_107_n10,
         DP_add_0_root_add_0_root_add_107_n9,
         DP_add_0_root_add_0_root_add_107_n8,
         DP_add_0_root_add_0_root_add_107_n7,
         DP_add_0_root_add_0_root_add_107_n6,
         DP_add_0_root_add_0_root_add_107_n5,
         DP_add_0_root_add_0_root_add_107_n4,
         DP_add_0_root_add_0_root_add_107_n3,
         DP_add_0_root_add_0_root_add_107_n2,
         DP_add_0_root_add_0_root_add_107_n1,
         DP_add_0_root_add_0_root_add_107_carry_1_,
         DP_add_0_root_add_0_root_add_107_carry_2_,
         DP_add_0_root_add_0_root_add_107_carry_3_,
         DP_add_0_root_add_0_root_add_107_carry_4_,
         DP_add_0_root_add_0_root_add_107_carry_6_,
         DP_add_0_root_add_0_root_add_107_carry_9_,
         DP_add_0_root_add_0_root_add_107_carry_12_,
         DP_sub_0_root_sub_0_root_sub_104_n82,
         DP_sub_0_root_sub_0_root_sub_104_n81,
         DP_sub_0_root_sub_0_root_sub_104_n80,
         DP_sub_0_root_sub_0_root_sub_104_n79,
         DP_sub_0_root_sub_0_root_sub_104_n78,
         DP_sub_0_root_sub_0_root_sub_104_n77,
         DP_sub_0_root_sub_0_root_sub_104_n76,
         DP_sub_0_root_sub_0_root_sub_104_n75,
         DP_sub_0_root_sub_0_root_sub_104_n74,
         DP_sub_0_root_sub_0_root_sub_104_n73,
         DP_sub_0_root_sub_0_root_sub_104_n72,
         DP_sub_0_root_sub_0_root_sub_104_n71,
         DP_sub_0_root_sub_0_root_sub_104_n70,
         DP_sub_0_root_sub_0_root_sub_104_n69,
         DP_sub_0_root_sub_0_root_sub_104_n68,
         DP_sub_0_root_sub_0_root_sub_104_n67,
         DP_sub_0_root_sub_0_root_sub_104_n66,
         DP_sub_0_root_sub_0_root_sub_104_n65,
         DP_sub_0_root_sub_0_root_sub_104_n64,
         DP_sub_0_root_sub_0_root_sub_104_n63,
         DP_sub_0_root_sub_0_root_sub_104_n62,
         DP_sub_0_root_sub_0_root_sub_104_n61,
         DP_sub_0_root_sub_0_root_sub_104_n60,
         DP_sub_0_root_sub_0_root_sub_104_n59,
         DP_sub_0_root_sub_0_root_sub_104_n58,
         DP_sub_0_root_sub_0_root_sub_104_n57,
         DP_sub_0_root_sub_0_root_sub_104_n56,
         DP_sub_0_root_sub_0_root_sub_104_n55,
         DP_sub_0_root_sub_0_root_sub_104_n54,
         DP_sub_0_root_sub_0_root_sub_104_n53,
         DP_sub_0_root_sub_0_root_sub_104_n52,
         DP_sub_0_root_sub_0_root_sub_104_n51,
         DP_sub_0_root_sub_0_root_sub_104_n50,
         DP_sub_0_root_sub_0_root_sub_104_n49,
         DP_sub_0_root_sub_0_root_sub_104_n48,
         DP_sub_0_root_sub_0_root_sub_104_n47,
         DP_sub_0_root_sub_0_root_sub_104_n46,
         DP_sub_0_root_sub_0_root_sub_104_n45,
         DP_sub_0_root_sub_0_root_sub_104_n44,
         DP_sub_0_root_sub_0_root_sub_104_n43,
         DP_sub_0_root_sub_0_root_sub_104_n42,
         DP_sub_0_root_sub_0_root_sub_104_n41,
         DP_sub_0_root_sub_0_root_sub_104_n40,
         DP_sub_0_root_sub_0_root_sub_104_n39,
         DP_sub_0_root_sub_0_root_sub_104_n38,
         DP_sub_0_root_sub_0_root_sub_104_n37,
         DP_sub_0_root_sub_0_root_sub_104_n36,
         DP_sub_0_root_sub_0_root_sub_104_n35,
         DP_sub_0_root_sub_0_root_sub_104_n34,
         DP_sub_0_root_sub_0_root_sub_104_n33,
         DP_sub_0_root_sub_0_root_sub_104_n32,
         DP_sub_0_root_sub_0_root_sub_104_n31,
         DP_sub_0_root_sub_0_root_sub_104_n30,
         DP_sub_0_root_sub_0_root_sub_104_n29,
         DP_sub_0_root_sub_0_root_sub_104_n28,
         DP_sub_0_root_sub_0_root_sub_104_n27,
         DP_sub_0_root_sub_0_root_sub_104_n26,
         DP_sub_0_root_sub_0_root_sub_104_n25,
         DP_sub_0_root_sub_0_root_sub_104_n24,
         DP_sub_0_root_sub_0_root_sub_104_n23,
         DP_sub_0_root_sub_0_root_sub_104_n22,
         DP_sub_0_root_sub_0_root_sub_104_n21,
         DP_sub_0_root_sub_0_root_sub_104_n20,
         DP_sub_0_root_sub_0_root_sub_104_n19,
         DP_sub_0_root_sub_0_root_sub_104_n18,
         DP_sub_0_root_sub_0_root_sub_104_n17,
         DP_sub_0_root_sub_0_root_sub_104_n16,
         DP_sub_0_root_sub_0_root_sub_104_n15,
         DP_sub_0_root_sub_0_root_sub_104_n14,
         DP_sub_0_root_sub_0_root_sub_104_n13,
         DP_sub_0_root_sub_0_root_sub_104_n12,
         DP_sub_0_root_sub_0_root_sub_104_n11,
         DP_sub_0_root_sub_0_root_sub_104_n10,
         DP_sub_0_root_sub_0_root_sub_104_n9,
         DP_sub_0_root_sub_0_root_sub_104_n8,
         DP_sub_0_root_sub_0_root_sub_104_n7,
         DP_sub_0_root_sub_0_root_sub_104_n6,
         DP_sub_0_root_sub_0_root_sub_104_n5,
         DP_sub_0_root_sub_0_root_sub_104_n4,
         DP_sub_0_root_sub_0_root_sub_104_n3,
         DP_sub_0_root_sub_0_root_sub_104_n2,
         DP_sub_0_root_sub_0_root_sub_104_n1,
         DP_sub_0_root_sub_0_root_sub_104_B_not_0_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_1_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_2_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_3_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_4_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_5_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_6_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_7_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_8_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_9_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_10_,
         DP_sub_0_root_sub_0_root_sub_104_B_not_12_,
         DP_sub_0_root_sub_0_root_sub_104_carry_2_,
         DP_sub_0_root_sub_0_root_sub_104_carry_3_,
         DP_sub_0_root_sub_0_root_sub_104_carry_4_,
         DP_sub_0_root_sub_0_root_sub_104_carry_5_,
         DP_sub_0_root_sub_0_root_sub_104_carry_6_,
         DP_sub_0_root_sub_0_root_sub_104_carry_7_,
         DP_sub_0_root_sub_0_root_sub_104_carry_8_,
         DP_sub_0_root_sub_0_root_sub_104_carry_9_,
         DP_sub_0_root_sub_0_root_sub_104_carry_10_,
         DP_sub_0_root_sub_0_root_sub_104_carry_12_, DP_mult_99_n660,
         DP_mult_99_n659, DP_mult_99_n658, DP_mult_99_n657, DP_mult_99_n656,
         DP_mult_99_n655, DP_mult_99_n654, DP_mult_99_n653, DP_mult_99_n652,
         DP_mult_99_n651, DP_mult_99_n650, DP_mult_99_n649, DP_mult_99_n648,
         DP_mult_99_n647, DP_mult_99_n646, DP_mult_99_n645, DP_mult_99_n644,
         DP_mult_99_n643, DP_mult_99_n642, DP_mult_99_n641, DP_mult_99_n640,
         DP_mult_99_n639, DP_mult_99_n638, DP_mult_99_n637, DP_mult_99_n636,
         DP_mult_99_n635, DP_mult_99_n634, DP_mult_99_n633, DP_mult_99_n632,
         DP_mult_99_n631, DP_mult_99_n630, DP_mult_99_n629, DP_mult_99_n628,
         DP_mult_99_n627, DP_mult_99_n626, DP_mult_99_n625, DP_mult_99_n624,
         DP_mult_99_n623, DP_mult_99_n622, DP_mult_99_n621, DP_mult_99_n620,
         DP_mult_99_n619, DP_mult_99_n618, DP_mult_99_n617, DP_mult_99_n616,
         DP_mult_99_n615, DP_mult_99_n614, DP_mult_99_n613, DP_mult_99_n612,
         DP_mult_99_n611, DP_mult_99_n610, DP_mult_99_n609, DP_mult_99_n608,
         DP_mult_99_n607, DP_mult_99_n606, DP_mult_99_n605, DP_mult_99_n604,
         DP_mult_99_n603, DP_mult_99_n602, DP_mult_99_n601, DP_mult_99_n600,
         DP_mult_99_n599, DP_mult_99_n598, DP_mult_99_n597, DP_mult_99_n596,
         DP_mult_99_n595, DP_mult_99_n594, DP_mult_99_n593, DP_mult_99_n592,
         DP_mult_99_n591, DP_mult_99_n590, DP_mult_99_n589, DP_mult_99_n588,
         DP_mult_99_n587, DP_mult_99_n586, DP_mult_99_n585, DP_mult_99_n584,
         DP_mult_99_n583, DP_mult_99_n582, DP_mult_99_n581, DP_mult_99_n580,
         DP_mult_99_n579, DP_mult_99_n578, DP_mult_99_n577, DP_mult_99_n576,
         DP_mult_99_n575, DP_mult_99_n574, DP_mult_99_n573, DP_mult_99_n572,
         DP_mult_99_n571, DP_mult_99_n570, DP_mult_99_n569, DP_mult_99_n568,
         DP_mult_99_n567, DP_mult_99_n566, DP_mult_99_n565, DP_mult_99_n564,
         DP_mult_99_n563, DP_mult_99_n562, DP_mult_99_n561, DP_mult_99_n560,
         DP_mult_99_n559, DP_mult_99_n558, DP_mult_99_n557, DP_mult_99_n556,
         DP_mult_99_n555, DP_mult_99_n554, DP_mult_99_n553, DP_mult_99_n552,
         DP_mult_99_n551, DP_mult_99_n550, DP_mult_99_n549, DP_mult_99_n548,
         DP_mult_99_n547, DP_mult_99_n546, DP_mult_99_n545, DP_mult_99_n544,
         DP_mult_99_n543, DP_mult_99_n542, DP_mult_99_n541, DP_mult_99_n540,
         DP_mult_99_n539, DP_mult_99_n538, DP_mult_99_n537, DP_mult_99_n536,
         DP_mult_99_n535, DP_mult_99_n534, DP_mult_99_n533, DP_mult_99_n532,
         DP_mult_99_n531, DP_mult_99_n530, DP_mult_99_n529, DP_mult_99_n528,
         DP_mult_99_n527, DP_mult_99_n526, DP_mult_99_n525, DP_mult_99_n524,
         DP_mult_99_n523, DP_mult_99_n522, DP_mult_99_n521, DP_mult_99_n520,
         DP_mult_99_n519, DP_mult_99_n337, DP_mult_99_n336, DP_mult_99_n335,
         DP_mult_99_n334, DP_mult_99_n333, DP_mult_99_n332, DP_mult_99_n331,
         DP_mult_99_n330, DP_mult_99_n329, DP_mult_99_n328, DP_mult_99_n327,
         DP_mult_99_n325, DP_mult_99_n324, DP_mult_99_n323, DP_mult_99_n322,
         DP_mult_99_n321, DP_mult_99_n320, DP_mult_99_n319, DP_mult_99_n318,
         DP_mult_99_n317, DP_mult_99_n316, DP_mult_99_n315, DP_mult_99_n314,
         DP_mult_99_n313, DP_mult_99_n312, DP_mult_99_n311, DP_mult_99_n310,
         DP_mult_99_n309, DP_mult_99_n308, DP_mult_99_n307, DP_mult_99_n306,
         DP_mult_99_n305, DP_mult_99_n303, DP_mult_99_n302, DP_mult_99_n301,
         DP_mult_99_n300, DP_mult_99_n299, DP_mult_99_n298, DP_mult_99_n297,
         DP_mult_99_n296, DP_mult_99_n295, DP_mult_99_n294, DP_mult_99_n293,
         DP_mult_99_n292, DP_mult_99_n291, DP_mult_99_n290, DP_mult_99_n289,
         DP_mult_99_n288, DP_mult_99_n287, DP_mult_99_n286, DP_mult_99_n285,
         DP_mult_99_n284, DP_mult_99_n283, DP_mult_99_n281, DP_mult_99_n280,
         DP_mult_99_n279, DP_mult_99_n278, DP_mult_99_n277, DP_mult_99_n276,
         DP_mult_99_n275, DP_mult_99_n274, DP_mult_99_n273, DP_mult_99_n272,
         DP_mult_99_n271, DP_mult_99_n270, DP_mult_99_n269, DP_mult_99_n268,
         DP_mult_99_n267, DP_mult_99_n266, DP_mult_99_n265, DP_mult_99_n264,
         DP_mult_99_n263, DP_mult_99_n259, DP_mult_99_n258, DP_mult_99_n257,
         DP_mult_99_n256, DP_mult_99_n255, DP_mult_99_n254, DP_mult_99_n253,
         DP_mult_99_n252, DP_mult_99_n251, DP_mult_99_n250, DP_mult_99_n249,
         DP_mult_99_n248, DP_mult_99_n247, DP_mult_99_n246, DP_mult_99_n245,
         DP_mult_99_n244, DP_mult_99_n243, DP_mult_99_n242, DP_mult_99_n241,
         DP_mult_99_n240, DP_mult_99_n239, DP_mult_99_n238, DP_mult_99_n237,
         DP_mult_99_n236, DP_mult_99_n235, DP_mult_99_n234, DP_mult_99_n233,
         DP_mult_99_n232, DP_mult_99_n231, DP_mult_99_n230, DP_mult_99_n229,
         DP_mult_99_n228, DP_mult_99_n227, DP_mult_99_n226, DP_mult_99_n225,
         DP_mult_99_n224, DP_mult_99_n223, DP_mult_99_n222, DP_mult_99_n221,
         DP_mult_99_n220, DP_mult_99_n219, DP_mult_99_n218, DP_mult_99_n217,
         DP_mult_99_n216, DP_mult_99_n215, DP_mult_99_n214, DP_mult_99_n213,
         DP_mult_99_n212, DP_mult_99_n211, DP_mult_99_n210, DP_mult_99_n209,
         DP_mult_99_n208, DP_mult_99_n207, DP_mult_99_n206, DP_mult_99_n205,
         DP_mult_99_n204, DP_mult_99_n203, DP_mult_99_n202, DP_mult_99_n201,
         DP_mult_99_n200, DP_mult_99_n199, DP_mult_99_n198, DP_mult_99_n197,
         DP_mult_99_n196, DP_mult_99_n195, DP_mult_99_n194, DP_mult_99_n193,
         DP_mult_99_n192, DP_mult_99_n191, DP_mult_99_n190, DP_mult_99_n189,
         DP_mult_99_n188, DP_mult_99_n187, DP_mult_99_n186, DP_mult_99_n185,
         DP_mult_99_n184, DP_mult_99_n183, DP_mult_99_n182, DP_mult_99_n181,
         DP_mult_99_n180, DP_mult_99_n179, DP_mult_99_n178, DP_mult_99_n177,
         DP_mult_99_n176, DP_mult_99_n175, DP_mult_99_n174, DP_mult_99_n173,
         DP_mult_99_n172, DP_mult_99_n171, DP_mult_99_n170, DP_mult_99_n169,
         DP_mult_99_n168, DP_mult_99_n167, DP_mult_99_n166, DP_mult_99_n165,
         DP_mult_99_n164, DP_mult_99_n163, DP_mult_99_n162, DP_mult_99_n161,
         DP_mult_99_n160, DP_mult_99_n159, DP_mult_99_n158, DP_mult_99_n157,
         DP_mult_99_n156, DP_mult_99_n155, DP_mult_99_n154, DP_mult_99_n153,
         DP_mult_99_n152, DP_mult_99_n151, DP_mult_99_n150, DP_mult_99_n149,
         DP_mult_99_n148, DP_mult_99_n147, DP_mult_99_n146, DP_mult_99_n145,
         DP_mult_99_n144, DP_mult_99_n143, DP_mult_99_n142, DP_mult_99_n141,
         DP_mult_99_n140, DP_mult_99_n139, DP_mult_99_n138, DP_mult_99_n126,
         DP_mult_99_n125, DP_mult_99_n124, DP_mult_99_n123, DP_mult_99_n122,
         DP_mult_99_n121, DP_mult_99_n120, DP_mult_99_n119, DP_mult_99_n118,
         DP_mult_99_n117, DP_mult_99_n116, DP_mult_99_n115, DP_mult_98_n661,
         DP_mult_98_n660, DP_mult_98_n659, DP_mult_98_n658, DP_mult_98_n657,
         DP_mult_98_n656, DP_mult_98_n655, DP_mult_98_n654, DP_mult_98_n653,
         DP_mult_98_n652, DP_mult_98_n651, DP_mult_98_n650, DP_mult_98_n649,
         DP_mult_98_n648, DP_mult_98_n647, DP_mult_98_n646, DP_mult_98_n645,
         DP_mult_98_n644, DP_mult_98_n643, DP_mult_98_n642, DP_mult_98_n641,
         DP_mult_98_n640, DP_mult_98_n639, DP_mult_98_n638, DP_mult_98_n637,
         DP_mult_98_n636, DP_mult_98_n635, DP_mult_98_n634, DP_mult_98_n633,
         DP_mult_98_n632, DP_mult_98_n631, DP_mult_98_n630, DP_mult_98_n629,
         DP_mult_98_n628, DP_mult_98_n627, DP_mult_98_n626, DP_mult_98_n625,
         DP_mult_98_n624, DP_mult_98_n623, DP_mult_98_n622, DP_mult_98_n621,
         DP_mult_98_n620, DP_mult_98_n619, DP_mult_98_n618, DP_mult_98_n617,
         DP_mult_98_n616, DP_mult_98_n615, DP_mult_98_n614, DP_mult_98_n613,
         DP_mult_98_n612, DP_mult_98_n611, DP_mult_98_n610, DP_mult_98_n609,
         DP_mult_98_n608, DP_mult_98_n607, DP_mult_98_n606, DP_mult_98_n605,
         DP_mult_98_n604, DP_mult_98_n603, DP_mult_98_n602, DP_mult_98_n601,
         DP_mult_98_n600, DP_mult_98_n599, DP_mult_98_n598, DP_mult_98_n597,
         DP_mult_98_n596, DP_mult_98_n595, DP_mult_98_n594, DP_mult_98_n593,
         DP_mult_98_n592, DP_mult_98_n591, DP_mult_98_n590, DP_mult_98_n589,
         DP_mult_98_n588, DP_mult_98_n587, DP_mult_98_n586, DP_mult_98_n585,
         DP_mult_98_n584, DP_mult_98_n583, DP_mult_98_n582, DP_mult_98_n581,
         DP_mult_98_n580, DP_mult_98_n579, DP_mult_98_n578, DP_mult_98_n577,
         DP_mult_98_n576, DP_mult_98_n575, DP_mult_98_n574, DP_mult_98_n573,
         DP_mult_98_n572, DP_mult_98_n571, DP_mult_98_n570, DP_mult_98_n569,
         DP_mult_98_n568, DP_mult_98_n567, DP_mult_98_n566, DP_mult_98_n565,
         DP_mult_98_n564, DP_mult_98_n563, DP_mult_98_n562, DP_mult_98_n561,
         DP_mult_98_n560, DP_mult_98_n559, DP_mult_98_n558, DP_mult_98_n557,
         DP_mult_98_n556, DP_mult_98_n555, DP_mult_98_n554, DP_mult_98_n553,
         DP_mult_98_n552, DP_mult_98_n551, DP_mult_98_n550, DP_mult_98_n549,
         DP_mult_98_n548, DP_mult_98_n547, DP_mult_98_n546, DP_mult_98_n545,
         DP_mult_98_n544, DP_mult_98_n543, DP_mult_98_n542, DP_mult_98_n541,
         DP_mult_98_n540, DP_mult_98_n539, DP_mult_98_n538, DP_mult_98_n537,
         DP_mult_98_n536, DP_mult_98_n535, DP_mult_98_n534, DP_mult_98_n533,
         DP_mult_98_n532, DP_mult_98_n531, DP_mult_98_n530, DP_mult_98_n529,
         DP_mult_98_n528, DP_mult_98_n527, DP_mult_98_n526, DP_mult_98_n525,
         DP_mult_98_n524, DP_mult_98_n523, DP_mult_98_n522, DP_mult_98_n521,
         DP_mult_98_n520, DP_mult_98_n519, DP_mult_98_n337, DP_mult_98_n336,
         DP_mult_98_n335, DP_mult_98_n334, DP_mult_98_n333, DP_mult_98_n332,
         DP_mult_98_n331, DP_mult_98_n330, DP_mult_98_n329, DP_mult_98_n328,
         DP_mult_98_n327, DP_mult_98_n325, DP_mult_98_n324, DP_mult_98_n323,
         DP_mult_98_n322, DP_mult_98_n321, DP_mult_98_n320, DP_mult_98_n319,
         DP_mult_98_n318, DP_mult_98_n317, DP_mult_98_n316, DP_mult_98_n315,
         DP_mult_98_n314, DP_mult_98_n313, DP_mult_98_n312, DP_mult_98_n311,
         DP_mult_98_n310, DP_mult_98_n309, DP_mult_98_n308, DP_mult_98_n307,
         DP_mult_98_n306, DP_mult_98_n305, DP_mult_98_n303, DP_mult_98_n302,
         DP_mult_98_n301, DP_mult_98_n300, DP_mult_98_n299, DP_mult_98_n298,
         DP_mult_98_n297, DP_mult_98_n296, DP_mult_98_n295, DP_mult_98_n294,
         DP_mult_98_n293, DP_mult_98_n292, DP_mult_98_n291, DP_mult_98_n290,
         DP_mult_98_n289, DP_mult_98_n288, DP_mult_98_n287, DP_mult_98_n286,
         DP_mult_98_n285, DP_mult_98_n284, DP_mult_98_n283, DP_mult_98_n281,
         DP_mult_98_n280, DP_mult_98_n279, DP_mult_98_n278, DP_mult_98_n277,
         DP_mult_98_n276, DP_mult_98_n275, DP_mult_98_n274, DP_mult_98_n273,
         DP_mult_98_n272, DP_mult_98_n271, DP_mult_98_n270, DP_mult_98_n269,
         DP_mult_98_n268, DP_mult_98_n267, DP_mult_98_n266, DP_mult_98_n265,
         DP_mult_98_n264, DP_mult_98_n263, DP_mult_98_n259, DP_mult_98_n258,
         DP_mult_98_n257, DP_mult_98_n256, DP_mult_98_n255, DP_mult_98_n254,
         DP_mult_98_n253, DP_mult_98_n252, DP_mult_98_n251, DP_mult_98_n250,
         DP_mult_98_n249, DP_mult_98_n248, DP_mult_98_n247, DP_mult_98_n246,
         DP_mult_98_n245, DP_mult_98_n244, DP_mult_98_n243, DP_mult_98_n242,
         DP_mult_98_n241, DP_mult_98_n240, DP_mult_98_n239, DP_mult_98_n238,
         DP_mult_98_n237, DP_mult_98_n236, DP_mult_98_n235, DP_mult_98_n234,
         DP_mult_98_n233, DP_mult_98_n232, DP_mult_98_n231, DP_mult_98_n230,
         DP_mult_98_n229, DP_mult_98_n228, DP_mult_98_n227, DP_mult_98_n226,
         DP_mult_98_n225, DP_mult_98_n224, DP_mult_98_n223, DP_mult_98_n222,
         DP_mult_98_n221, DP_mult_98_n220, DP_mult_98_n219, DP_mult_98_n218,
         DP_mult_98_n217, DP_mult_98_n216, DP_mult_98_n215, DP_mult_98_n214,
         DP_mult_98_n213, DP_mult_98_n212, DP_mult_98_n211, DP_mult_98_n210,
         DP_mult_98_n209, DP_mult_98_n208, DP_mult_98_n207, DP_mult_98_n206,
         DP_mult_98_n205, DP_mult_98_n204, DP_mult_98_n203, DP_mult_98_n202,
         DP_mult_98_n201, DP_mult_98_n200, DP_mult_98_n199, DP_mult_98_n198,
         DP_mult_98_n197, DP_mult_98_n196, DP_mult_98_n195, DP_mult_98_n194,
         DP_mult_98_n193, DP_mult_98_n192, DP_mult_98_n191, DP_mult_98_n190,
         DP_mult_98_n189, DP_mult_98_n188, DP_mult_98_n187, DP_mult_98_n186,
         DP_mult_98_n185, DP_mult_98_n184, DP_mult_98_n183, DP_mult_98_n182,
         DP_mult_98_n181, DP_mult_98_n180, DP_mult_98_n179, DP_mult_98_n178,
         DP_mult_98_n177, DP_mult_98_n176, DP_mult_98_n175, DP_mult_98_n174,
         DP_mult_98_n173, DP_mult_98_n172, DP_mult_98_n171, DP_mult_98_n170,
         DP_mult_98_n169, DP_mult_98_n168, DP_mult_98_n167, DP_mult_98_n166,
         DP_mult_98_n165, DP_mult_98_n164, DP_mult_98_n163, DP_mult_98_n162,
         DP_mult_98_n161, DP_mult_98_n160, DP_mult_98_n159, DP_mult_98_n158,
         DP_mult_98_n157, DP_mult_98_n156, DP_mult_98_n155, DP_mult_98_n154,
         DP_mult_98_n153, DP_mult_98_n152, DP_mult_98_n151, DP_mult_98_n150,
         DP_mult_98_n149, DP_mult_98_n148, DP_mult_98_n147, DP_mult_98_n146,
         DP_mult_98_n145, DP_mult_98_n144, DP_mult_98_n143, DP_mult_98_n142,
         DP_mult_98_n141, DP_mult_98_n140, DP_mult_98_n139, DP_mult_98_n138,
         DP_mult_98_n126, DP_mult_98_n125, DP_mult_98_n124, DP_mult_98_n123,
         DP_mult_98_n122, DP_mult_98_n121, DP_mult_98_n120, DP_mult_98_n119,
         DP_mult_98_n118, DP_mult_98_n117, DP_mult_98_n116, DP_mult_98_n115,
         DP_mult_97_n769, DP_mult_97_n768, DP_mult_97_n767, DP_mult_97_n766,
         DP_mult_97_n765, DP_mult_97_n764, DP_mult_97_n763, DP_mult_97_n762,
         DP_mult_97_n761, DP_mult_97_n760, DP_mult_97_n759, DP_mult_97_n758,
         DP_mult_97_n757, DP_mult_97_n756, DP_mult_97_n755, DP_mult_97_n754,
         DP_mult_97_n753, DP_mult_97_n752, DP_mult_97_n751, DP_mult_97_n750,
         DP_mult_97_n749, DP_mult_97_n748, DP_mult_97_n747, DP_mult_97_n746,
         DP_mult_97_n745, DP_mult_97_n744, DP_mult_97_n743, DP_mult_97_n742,
         DP_mult_97_n741, DP_mult_97_n740, DP_mult_97_n739, DP_mult_97_n738,
         DP_mult_97_n737, DP_mult_97_n736, DP_mult_97_n735, DP_mult_97_n734,
         DP_mult_97_n733, DP_mult_97_n732, DP_mult_97_n731, DP_mult_97_n730,
         DP_mult_97_n729, DP_mult_97_n728, DP_mult_97_n727, DP_mult_97_n726,
         DP_mult_97_n725, DP_mult_97_n724, DP_mult_97_n723, DP_mult_97_n722,
         DP_mult_97_n721, DP_mult_97_n720, DP_mult_97_n719, DP_mult_97_n718,
         DP_mult_97_n717, DP_mult_97_n716, DP_mult_97_n715, DP_mult_97_n714,
         DP_mult_97_n713, DP_mult_97_n712, DP_mult_97_n711, DP_mult_97_n710,
         DP_mult_97_n709, DP_mult_97_n708, DP_mult_97_n707, DP_mult_97_n706,
         DP_mult_97_n705, DP_mult_97_n704, DP_mult_97_n703, DP_mult_97_n702,
         DP_mult_97_n701, DP_mult_97_n700, DP_mult_97_n699, DP_mult_97_n698,
         DP_mult_97_n697, DP_mult_97_n696, DP_mult_97_n695, DP_mult_97_n694,
         DP_mult_97_n693, DP_mult_97_n692, DP_mult_97_n691, DP_mult_97_n690,
         DP_mult_97_n689, DP_mult_97_n688, DP_mult_97_n687, DP_mult_97_n686,
         DP_mult_97_n685, DP_mult_97_n684, DP_mult_97_n683, DP_mult_97_n682,
         DP_mult_97_n681, DP_mult_97_n680, DP_mult_97_n679, DP_mult_97_n678,
         DP_mult_97_n677, DP_mult_97_n676, DP_mult_97_n675, DP_mult_97_n674,
         DP_mult_97_n673, DP_mult_97_n672, DP_mult_97_n671, DP_mult_97_n670,
         DP_mult_97_n669, DP_mult_97_n668, DP_mult_97_n667, DP_mult_97_n666,
         DP_mult_97_n665, DP_mult_97_n664, DP_mult_97_n663, DP_mult_97_n662,
         DP_mult_97_n661, DP_mult_97_n620, DP_mult_97_n619, DP_mult_97_n618,
         DP_mult_97_n617, DP_mult_97_n616, DP_mult_97_n615, DP_mult_97_n614,
         DP_mult_97_n613, DP_mult_97_n612, DP_mult_97_n611, DP_mult_97_n610,
         DP_mult_97_n609, DP_mult_97_n608, DP_mult_97_n607, DP_mult_97_n606,
         DP_mult_97_n605, DP_mult_97_n604, DP_mult_97_n603, DP_mult_97_n602,
         DP_mult_97_n601, DP_mult_97_n600, DP_mult_97_n599, DP_mult_97_n597,
         DP_mult_97_n596, DP_mult_97_n595, DP_mult_97_n594, DP_mult_97_n593,
         DP_mult_97_n592, DP_mult_97_n591, DP_mult_97_n590, DP_mult_97_n589,
         DP_mult_97_n587, DP_mult_97_n585, DP_mult_97_n584, DP_mult_97_n583,
         DP_mult_97_n582, DP_mult_97_n581, DP_mult_97_n580, DP_mult_97_n579,
         DP_mult_97_n576, DP_mult_97_n575, DP_mult_97_n574, DP_mult_97_n572,
         DP_mult_97_n571, DP_mult_97_n568, DP_mult_97_n567, DP_mult_97_n566,
         DP_mult_97_n565, DP_mult_97_n564, DP_mult_97_n563, DP_mult_97_n562,
         DP_mult_97_n561, DP_mult_97_n560, DP_mult_97_n559, DP_mult_97_n558,
         DP_mult_97_n557, DP_mult_97_n555, DP_mult_97_n554, DP_mult_97_n553,
         DP_mult_97_n552, DP_mult_97_n551, DP_mult_97_n550, DP_mult_97_n549,
         DP_mult_97_n548, DP_mult_97_n547, DP_mult_97_n546, DP_mult_97_n545,
         DP_mult_97_n544, DP_mult_97_n543, DP_mult_97_n542, DP_mult_97_n541,
         DP_mult_97_n540, DP_mult_97_n539, DP_mult_97_n538, DP_mult_97_n537,
         DP_mult_97_n536, DP_mult_97_n535, DP_mult_97_n534, DP_mult_97_n533,
         DP_mult_97_n532, DP_mult_97_n531, DP_mult_97_n530, DP_mult_97_n529,
         DP_mult_97_n528, DP_mult_97_n527, DP_mult_97_n526, DP_mult_97_n525,
         DP_mult_97_n524, DP_mult_97_n523, DP_mult_97_n522, DP_mult_97_n521,
         DP_mult_97_n520, DP_mult_97_n519, DP_mult_97_n518, DP_mult_97_n517,
         DP_mult_97_n516, DP_mult_97_n515, DP_mult_97_n514, DP_mult_97_n513,
         DP_mult_97_n512, DP_mult_97_n511, DP_mult_97_n510, DP_mult_97_n509,
         DP_mult_97_n508, DP_mult_97_n507, DP_mult_97_n506, DP_mult_97_n505,
         DP_mult_97_n504, DP_mult_97_n503, DP_mult_97_n502, DP_mult_97_n501,
         DP_mult_97_n500, DP_mult_97_n499, DP_mult_97_n498, DP_mult_97_n497,
         DP_mult_97_n496, DP_mult_97_n495, DP_mult_97_n494, DP_mult_97_n493,
         DP_mult_97_n492, DP_mult_97_n491, DP_mult_97_n490, DP_mult_97_n489,
         DP_mult_97_n488, DP_mult_97_n487, DP_mult_97_n486, DP_mult_97_n485,
         DP_mult_97_n484, DP_mult_97_n483, DP_mult_97_n482, DP_mult_97_n481,
         DP_mult_97_n480, DP_mult_97_n479, DP_mult_97_n478, DP_mult_97_n477,
         DP_mult_97_n476, DP_mult_97_n475, DP_mult_97_n474, DP_mult_97_n473,
         DP_mult_97_n472, DP_mult_97_n471, DP_mult_97_n470, DP_mult_97_n469,
         DP_mult_97_n467, DP_mult_97_n466, DP_mult_97_n465, DP_mult_97_n464,
         DP_mult_97_n463, DP_mult_97_n462, DP_mult_97_n461, DP_mult_97_n460,
         DP_mult_97_n459, DP_mult_97_n458, DP_mult_97_n457, DP_mult_97_n456,
         DP_mult_97_n454, DP_mult_97_n453, DP_mult_97_n452, DP_mult_97_n451,
         DP_mult_97_n450, DP_mult_97_n449, DP_mult_97_n448, DP_mult_97_n447,
         DP_mult_97_n446, DP_mult_97_n445, DP_mult_97_n444, DP_mult_97_n443,
         DP_mult_97_n441, DP_mult_97_n440, DP_mult_97_n439, DP_mult_97_n438,
         DP_mult_97_n437, DP_mult_97_n436, DP_mult_97_n435, DP_mult_97_n434,
         DP_mult_97_n433, DP_mult_97_n432, DP_mult_97_n431, DP_mult_97_n430,
         DP_mult_97_n428, DP_mult_97_n427, DP_mult_97_n426, DP_mult_97_n425,
         DP_mult_97_n423, DP_mult_97_n422, DP_mult_97_n421, DP_mult_97_n420,
         DP_mult_97_n419, DP_mult_97_n418, DP_mult_97_n417, DP_mult_97_n415,
         DP_mult_97_n414, DP_mult_97_n413, DP_mult_97_n412, DP_mult_97_n411,
         DP_mult_97_n410, DP_mult_97_n409, DP_mult_97_n408, DP_mult_97_n407,
         DP_mult_97_n406, DP_mult_97_n405, DP_mult_97_n404, DP_mult_97_n403,
         DP_mult_97_n402, DP_mult_97_n401, DP_mult_97_n400, DP_mult_97_n399,
         DP_mult_97_n398, DP_mult_97_n397, DP_mult_97_n396, DP_mult_97_n395,
         DP_mult_97_n394, DP_mult_97_n393, DP_mult_97_n392, DP_mult_97_n391,
         DP_mult_97_n390, DP_mult_97_n389, DP_mult_97_n388, DP_mult_97_n387,
         DP_mult_97_n386, DP_mult_97_n385, DP_mult_97_n384, DP_mult_97_n383,
         DP_mult_97_n382, DP_mult_97_n381, DP_mult_97_n380, DP_mult_97_n379,
         DP_mult_97_n378, DP_mult_97_n377, DP_mult_97_n376, DP_mult_97_n375,
         DP_mult_97_n374, DP_mult_97_n373, DP_mult_97_n372, DP_mult_97_n371,
         DP_mult_97_n370, DP_mult_97_n369, DP_mult_97_n368, DP_mult_97_n367,
         DP_mult_97_n366, DP_mult_97_n365, DP_mult_97_n364, DP_mult_97_n363,
         DP_mult_97_n362, DP_mult_97_n361, DP_mult_97_n360, DP_mult_97_n359,
         DP_mult_97_n358, DP_mult_97_n357, DP_mult_97_n356, DP_mult_97_n355,
         DP_mult_97_n354, DP_mult_97_n353, DP_mult_97_n352, DP_mult_97_n351,
         DP_mult_97_n350, DP_mult_97_n349, DP_mult_97_n348, DP_mult_97_n347,
         DP_mult_97_n346, DP_mult_97_n345, DP_mult_97_n344, DP_mult_97_n343,
         DP_mult_97_n342, DP_mult_97_n341, DP_mult_97_n340, DP_mult_97_n339,
         DP_mult_97_n338, DP_mult_97_n337, DP_mult_97_n336, DP_mult_97_n335,
         DP_mult_97_n334, DP_mult_97_n333, DP_mult_97_n332, DP_mult_97_n331,
         DP_mult_97_n330, DP_mult_97_n329, DP_mult_97_n328, DP_mult_97_n327,
         DP_mult_97_n326, DP_mult_97_n325, DP_mult_97_n324, DP_mult_97_n323,
         DP_mult_97_n322, DP_mult_97_n321, DP_mult_97_n320, DP_mult_97_n319,
         DP_mult_97_n318, DP_mult_97_n317, DP_mult_97_n316, DP_mult_97_n315,
         DP_mult_97_n314, DP_mult_97_n313, DP_mult_97_n312, DP_mult_97_n311,
         DP_mult_97_n310, DP_mult_97_n309, DP_mult_97_n308, DP_mult_97_n307,
         DP_mult_97_n306, DP_mult_97_n305, DP_mult_97_n304, DP_mult_97_n303,
         DP_mult_97_n302, DP_mult_97_n301, DP_mult_97_n300, DP_mult_97_n299,
         DP_mult_97_n298, DP_mult_97_n297, DP_mult_97_n296, DP_mult_97_n295,
         DP_mult_97_n294, DP_mult_97_n293, DP_mult_97_n292, DP_mult_97_n291,
         DP_mult_97_n290, DP_mult_97_n289, DP_mult_97_n288, DP_mult_97_n287,
         DP_mult_97_n286, DP_mult_97_n285, DP_mult_97_n284, DP_mult_97_n283,
         DP_mult_97_n282, DP_mult_97_n281, DP_mult_97_n280, DP_mult_97_n279,
         DP_mult_97_n278, DP_mult_97_n275, DP_mult_97_n273, DP_mult_97_n260,
         DP_mult_97_n259, DP_mult_97_n258, DP_mult_97_n257, DP_mult_97_n256,
         DP_mult_97_n255, DP_mult_97_n254, DP_mult_97_n253, DP_mult_97_n252,
         DP_mult_97_n251, DP_mult_97_n250, DP_mult_97_n249, DP_mult_97_n248,
         DP_mult_97_n247, DP_mult_97_n242, DP_mult_97_n233, DP_mult_97_n232,
         DP_mult_97_n230, DP_mult_97_n229, DP_mult_97_n228, DP_mult_97_n227,
         DP_mult_97_n226, DP_mult_97_n225, DP_mult_97_n224, DP_mult_97_n223,
         DP_mult_97_n222, DP_mult_97_n221, DP_mult_97_n220, DP_mult_97_n219,
         DP_mult_97_n218, DP_mult_97_n216, DP_mult_97_n215, DP_mult_97_n214,
         DP_mult_97_n213, DP_mult_97_n212, DP_mult_97_n211, DP_mult_97_n210,
         DP_mult_97_n209, DP_mult_97_n208, DP_mult_97_n207, DP_mult_97_n206,
         DP_mult_97_n205, DP_mult_97_n203, DP_mult_97_n202, DP_mult_97_n201,
         DP_mult_97_n200, DP_mult_97_n199, DP_mult_97_n198, DP_mult_97_n197,
         DP_mult_97_n196, DP_mult_97_n195, DP_mult_97_n194, DP_mult_97_n193,
         DP_mult_97_n192, DP_mult_97_n191, DP_mult_97_n190, DP_mult_97_n185,
         DP_mult_97_n184, DP_mult_97_n183, DP_mult_97_n181, DP_mult_97_n179,
         DP_mult_97_n178, DP_mult_97_n177, DP_mult_97_n176, DP_mult_97_n175,
         DP_mult_97_n174, DP_mult_97_n172, DP_mult_97_n170, DP_mult_97_n169,
         DP_mult_97_n168, DP_mult_97_n167, DP_mult_97_n166, DP_mult_97_n165,
         DP_mult_97_n163, DP_mult_97_n159, DP_mult_97_n158, DP_mult_97_n157,
         DP_mult_97_n156, DP_mult_97_n155, DP_mult_97_n154, DP_mult_97_n152,
         DP_mult_97_n150, DP_mult_97_n149, DP_mult_97_n148, DP_mult_97_n147,
         DP_mult_97_n146, DP_mult_97_n145, DP_mult_97_n143, DP_mult_97_n141,
         DP_mult_97_n139, DP_mult_97_n137, DP_mult_97_n136, DP_mult_97_n135,
         DP_mult_97_n134, DP_mult_97_n133, DP_mult_97_n132, DP_mult_97_n131,
         DP_mult_97_n130, DP_mult_97_n129, DP_mult_97_n128, DP_mult_97_n127,
         DP_mult_97_n126, DP_mult_97_n124, DP_mult_97_n120, DP_mult_97_n119,
         DP_mult_97_n118, DP_mult_97_n105, DP_mult_97_n104, DP_mult_97_n103,
         DP_mult_97_n98, DP_mult_97_n89, DP_mult_97_n88, DP_mult_97_n87,
         DP_mult_97_n82, DP_mult_97_n77, DP_mult_97_n73, DP_mult_97_n69,
         DP_mult_97_n64, DP_mult_97_n48, DP_mult_97_n47, DP_mult_97_n40,
         DP_mult_97_n35, DP_mult_97_n30, DP_mult_97_n26, DP_mult_97_n24,
         DP_mult_97_n14, DP_mult_97_n10, DP_mult_97_n9, DP_mult_97_n8,
         DP_mult_96_n687, DP_mult_96_n686, DP_mult_96_n685, DP_mult_96_n684,
         DP_mult_96_n683, DP_mult_96_n682, DP_mult_96_n681, DP_mult_96_n680,
         DP_mult_96_n679, DP_mult_96_n678, DP_mult_96_n677, DP_mult_96_n676,
         DP_mult_96_n675, DP_mult_96_n674, DP_mult_96_n673, DP_mult_96_n672,
         DP_mult_96_n671, DP_mult_96_n670, DP_mult_96_n669, DP_mult_96_n668,
         DP_mult_96_n667, DP_mult_96_n666, DP_mult_96_n665, DP_mult_96_n664,
         DP_mult_96_n663, DP_mult_96_n662, DP_mult_96_n661, DP_mult_96_n620,
         DP_mult_96_n619, DP_mult_96_n618, DP_mult_96_n617, DP_mult_96_n616,
         DP_mult_96_n615, DP_mult_96_n614, DP_mult_96_n613, DP_mult_96_n612,
         DP_mult_96_n611, DP_mult_96_n610, DP_mult_96_n609, DP_mult_96_n608,
         DP_mult_96_n607, DP_mult_96_n606, DP_mult_96_n605, DP_mult_96_n604,
         DP_mult_96_n603, DP_mult_96_n602, DP_mult_96_n601, DP_mult_96_n600,
         DP_mult_96_n599, DP_mult_96_n598, DP_mult_96_n597, DP_mult_96_n596,
         DP_mult_96_n595, DP_mult_96_n594, DP_mult_96_n593, DP_mult_96_n592,
         DP_mult_96_n591, DP_mult_96_n590, DP_mult_96_n589, DP_mult_96_n588,
         DP_mult_96_n587, DP_mult_96_n586, DP_mult_96_n585, DP_mult_96_n584,
         DP_mult_96_n583, DP_mult_96_n582, DP_mult_96_n581, DP_mult_96_n580,
         DP_mult_96_n579, DP_mult_96_n577, DP_mult_96_n576, DP_mult_96_n575,
         DP_mult_96_n574, DP_mult_96_n573, DP_mult_96_n572, DP_mult_96_n571,
         DP_mult_96_n570, DP_mult_96_n569, DP_mult_96_n568, DP_mult_96_n567,
         DP_mult_96_n566, DP_mult_96_n565, DP_mult_96_n564, DP_mult_96_n563,
         DP_mult_96_n562, DP_mult_96_n561, DP_mult_96_n560, DP_mult_96_n559,
         DP_mult_96_n558, DP_mult_96_n557, DP_mult_96_n556, DP_mult_96_n555,
         DP_mult_96_n554, DP_mult_96_n553, DP_mult_96_n552, DP_mult_96_n551,
         DP_mult_96_n550, DP_mult_96_n549, DP_mult_96_n548, DP_mult_96_n547,
         DP_mult_96_n546, DP_mult_96_n545, DP_mult_96_n544, DP_mult_96_n543,
         DP_mult_96_n542, DP_mult_96_n541, DP_mult_96_n540, DP_mult_96_n539,
         DP_mult_96_n538, DP_mult_96_n537, DP_mult_96_n536, DP_mult_96_n535,
         DP_mult_96_n534, DP_mult_96_n533, DP_mult_96_n532, DP_mult_96_n531,
         DP_mult_96_n530, DP_mult_96_n529, DP_mult_96_n528, DP_mult_96_n527,
         DP_mult_96_n526, DP_mult_96_n525, DP_mult_96_n524, DP_mult_96_n523,
         DP_mult_96_n522, DP_mult_96_n521, DP_mult_96_n520, DP_mult_96_n519,
         DP_mult_96_n518, DP_mult_96_n517, DP_mult_96_n516, DP_mult_96_n515,
         DP_mult_96_n514, DP_mult_96_n513, DP_mult_96_n512, DP_mult_96_n511,
         DP_mult_96_n510, DP_mult_96_n509, DP_mult_96_n508, DP_mult_96_n507,
         DP_mult_96_n506, DP_mult_96_n505, DP_mult_96_n504, DP_mult_96_n503,
         DP_mult_96_n502, DP_mult_96_n501, DP_mult_96_n500, DP_mult_96_n499,
         DP_mult_96_n498, DP_mult_96_n497, DP_mult_96_n496, DP_mult_96_n495,
         DP_mult_96_n494, DP_mult_96_n493, DP_mult_96_n492, DP_mult_96_n491,
         DP_mult_96_n490, DP_mult_96_n489, DP_mult_96_n488, DP_mult_96_n487,
         DP_mult_96_n486, DP_mult_96_n485, DP_mult_96_n484, DP_mult_96_n483,
         DP_mult_96_n482, DP_mult_96_n481, DP_mult_96_n480, DP_mult_96_n479,
         DP_mult_96_n478, DP_mult_96_n477, DP_mult_96_n476, DP_mult_96_n475,
         DP_mult_96_n474, DP_mult_96_n473, DP_mult_96_n472, DP_mult_96_n471,
         DP_mult_96_n470, DP_mult_96_n469, DP_mult_96_n467, DP_mult_96_n466,
         DP_mult_96_n465, DP_mult_96_n464, DP_mult_96_n463, DP_mult_96_n462,
         DP_mult_96_n461, DP_mult_96_n460, DP_mult_96_n459, DP_mult_96_n458,
         DP_mult_96_n457, DP_mult_96_n456, DP_mult_96_n454, DP_mult_96_n453,
         DP_mult_96_n452, DP_mult_96_n451, DP_mult_96_n450, DP_mult_96_n449,
         DP_mult_96_n448, DP_mult_96_n447, DP_mult_96_n446, DP_mult_96_n445,
         DP_mult_96_n444, DP_mult_96_n443, DP_mult_96_n441, DP_mult_96_n440,
         DP_mult_96_n439, DP_mult_96_n438, DP_mult_96_n437, DP_mult_96_n436,
         DP_mult_96_n435, DP_mult_96_n434, DP_mult_96_n433, DP_mult_96_n432,
         DP_mult_96_n431, DP_mult_96_n430, DP_mult_96_n428, DP_mult_96_n427,
         DP_mult_96_n426, DP_mult_96_n425, DP_mult_96_n424, DP_mult_96_n423,
         DP_mult_96_n422, DP_mult_96_n421, DP_mult_96_n420, DP_mult_96_n419,
         DP_mult_96_n418, DP_mult_96_n417, DP_mult_96_n415, DP_mult_96_n414,
         DP_mult_96_n413, DP_mult_96_n412, DP_mult_96_n411, DP_mult_96_n410,
         DP_mult_96_n409, DP_mult_96_n408, DP_mult_96_n407, DP_mult_96_n406,
         DP_mult_96_n405, DP_mult_96_n404, DP_mult_96_n403, DP_mult_96_n402,
         DP_mult_96_n401, DP_mult_96_n400, DP_mult_96_n399, DP_mult_96_n398,
         DP_mult_96_n397, DP_mult_96_n396, DP_mult_96_n395, DP_mult_96_n394,
         DP_mult_96_n393, DP_mult_96_n392, DP_mult_96_n391, DP_mult_96_n390,
         DP_mult_96_n389, DP_mult_96_n388, DP_mult_96_n387, DP_mult_96_n386,
         DP_mult_96_n385, DP_mult_96_n384, DP_mult_96_n383, DP_mult_96_n382,
         DP_mult_96_n381, DP_mult_96_n380, DP_mult_96_n379, DP_mult_96_n378,
         DP_mult_96_n377, DP_mult_96_n376, DP_mult_96_n375, DP_mult_96_n374,
         DP_mult_96_n373, DP_mult_96_n372, DP_mult_96_n371, DP_mult_96_n370,
         DP_mult_96_n369, DP_mult_96_n368, DP_mult_96_n367, DP_mult_96_n366,
         DP_mult_96_n365, DP_mult_96_n364, DP_mult_96_n363, DP_mult_96_n362,
         DP_mult_96_n361, DP_mult_96_n360, DP_mult_96_n359, DP_mult_96_n358,
         DP_mult_96_n357, DP_mult_96_n356, DP_mult_96_n355, DP_mult_96_n354,
         DP_mult_96_n353, DP_mult_96_n352, DP_mult_96_n351, DP_mult_96_n350,
         DP_mult_96_n349, DP_mult_96_n348, DP_mult_96_n347, DP_mult_96_n346,
         DP_mult_96_n345, DP_mult_96_n344, DP_mult_96_n343, DP_mult_96_n342,
         DP_mult_96_n341, DP_mult_96_n340, DP_mult_96_n339, DP_mult_96_n338,
         DP_mult_96_n337, DP_mult_96_n336, DP_mult_96_n335, DP_mult_96_n334,
         DP_mult_96_n333, DP_mult_96_n332, DP_mult_96_n331, DP_mult_96_n330,
         DP_mult_96_n329, DP_mult_96_n328, DP_mult_96_n327, DP_mult_96_n326,
         DP_mult_96_n325, DP_mult_96_n324, DP_mult_96_n323, DP_mult_96_n322,
         DP_mult_96_n321, DP_mult_96_n320, DP_mult_96_n319, DP_mult_96_n318,
         DP_mult_96_n317, DP_mult_96_n316, DP_mult_96_n315, DP_mult_96_n314,
         DP_mult_96_n313, DP_mult_96_n312, DP_mult_96_n311, DP_mult_96_n310,
         DP_mult_96_n309, DP_mult_96_n308, DP_mult_96_n307, DP_mult_96_n306,
         DP_mult_96_n305, DP_mult_96_n304, DP_mult_96_n303, DP_mult_96_n302,
         DP_mult_96_n301, DP_mult_96_n300, DP_mult_96_n299, DP_mult_96_n298,
         DP_mult_96_n297, DP_mult_96_n296, DP_mult_96_n295, DP_mult_96_n294,
         DP_mult_96_n293, DP_mult_96_n292, DP_mult_96_n291, DP_mult_96_n290,
         DP_mult_96_n289, DP_mult_96_n288, DP_mult_96_n287, DP_mult_96_n286,
         DP_mult_96_n285, DP_mult_96_n284, DP_mult_96_n283, DP_mult_96_n282,
         DP_mult_96_n281, DP_mult_96_n280, DP_mult_96_n279, DP_mult_96_n278,
         DP_mult_96_n277, DP_mult_96_n275, DP_mult_96_n273, DP_mult_96_n269,
         DP_mult_96_n260, DP_mult_96_n259, DP_mult_96_n258, DP_mult_96_n257,
         DP_mult_96_n256, DP_mult_96_n255, DP_mult_96_n254, DP_mult_96_n253,
         DP_mult_96_n252, DP_mult_96_n251, DP_mult_96_n250, DP_mult_96_n249,
         DP_mult_96_n248, DP_mult_96_n247, DP_mult_96_n242, DP_mult_96_n233,
         DP_mult_96_n232, DP_mult_96_n231, DP_mult_96_n230, DP_mult_96_n229,
         DP_mult_96_n228, DP_mult_96_n227, DP_mult_96_n226, DP_mult_96_n225,
         DP_mult_96_n224, DP_mult_96_n223, DP_mult_96_n222, DP_mult_96_n221,
         DP_mult_96_n220, DP_mult_96_n219, DP_mult_96_n218, DP_mult_96_n217,
         DP_mult_96_n216, DP_mult_96_n215, DP_mult_96_n214, DP_mult_96_n213,
         DP_mult_96_n212, DP_mult_96_n211, DP_mult_96_n210, DP_mult_96_n209,
         DP_mult_96_n208, DP_mult_96_n207, DP_mult_96_n206, DP_mult_96_n205,
         DP_mult_96_n204, DP_mult_96_n203, DP_mult_96_n202, DP_mult_96_n201,
         DP_mult_96_n200, DP_mult_96_n199, DP_mult_96_n198, DP_mult_96_n197,
         DP_mult_96_n196, DP_mult_96_n195, DP_mult_96_n194, DP_mult_96_n193,
         DP_mult_96_n192, DP_mult_96_n191, DP_mult_96_n189, DP_mult_96_n186,
         DP_mult_96_n185, DP_mult_96_n184, DP_mult_96_n183, DP_mult_96_n181,
         DP_mult_96_n179, DP_mult_96_n178, DP_mult_96_n177, DP_mult_96_n176,
         DP_mult_96_n175, DP_mult_96_n174, DP_mult_96_n172, DP_mult_96_n170,
         DP_mult_96_n169, DP_mult_96_n168, DP_mult_96_n167, DP_mult_96_n166,
         DP_mult_96_n165, DP_mult_96_n164, DP_mult_96_n163, DP_mult_96_n161,
         DP_mult_96_n160, DP_mult_96_n159, DP_mult_96_n158, DP_mult_96_n157,
         DP_mult_96_n156, DP_mult_96_n155, DP_mult_96_n154, DP_mult_96_n152,
         DP_mult_96_n150, DP_mult_96_n149, DP_mult_96_n148, DP_mult_96_n147,
         DP_mult_96_n146, DP_mult_96_n145, DP_mult_96_n143, DP_mult_96_n141,
         DP_mult_96_n139, DP_mult_96_n137, DP_mult_96_n136, DP_mult_96_n135,
         DP_mult_96_n134, DP_mult_96_n133, DP_mult_96_n132, DP_mult_96_n131,
         DP_mult_96_n130, DP_mult_96_n129, DP_mult_96_n128, DP_mult_96_n127,
         DP_mult_96_n126, DP_mult_96_n124, DP_mult_96_n122, DP_mult_96_n121,
         DP_mult_96_n120, DP_mult_96_n119, DP_mult_96_n118, DP_mult_96_n117,
         DP_mult_96_n116, DP_mult_96_n115, DP_mult_96_n114, DP_mult_96_n113,
         DP_mult_96_n111, DP_mult_96_n109, DP_mult_96_n105, DP_mult_96_n104,
         DP_mult_96_n103, DP_mult_96_n93, DP_mult_96_n89, DP_mult_96_n87,
         DP_mult_96_n77, DP_mult_96_n73, DP_mult_96_n69, DP_mult_96_n57,
         DP_mult_96_n48, DP_mult_96_n40, DP_mult_96_n30, DP_mult_96_n26,
         DP_mult_96_n24, DP_mult_96_n14, DP_mult_96_n10, DP_mult_96_n8,
         DP_sub_1_root_sub_0_root_sub_104_n157,
         DP_sub_1_root_sub_0_root_sub_104_n156,
         DP_sub_1_root_sub_0_root_sub_104_n155,
         DP_sub_1_root_sub_0_root_sub_104_n154,
         DP_sub_1_root_sub_0_root_sub_104_n153,
         DP_sub_1_root_sub_0_root_sub_104_n152,
         DP_sub_1_root_sub_0_root_sub_104_n151,
         DP_sub_1_root_sub_0_root_sub_104_n150,
         DP_sub_1_root_sub_0_root_sub_104_n149,
         DP_sub_1_root_sub_0_root_sub_104_n148,
         DP_sub_1_root_sub_0_root_sub_104_n147,
         DP_sub_1_root_sub_0_root_sub_104_n146,
         DP_sub_1_root_sub_0_root_sub_104_n145,
         DP_sub_1_root_sub_0_root_sub_104_n101,
         DP_sub_1_root_sub_0_root_sub_104_n96,
         DP_sub_1_root_sub_0_root_sub_104_n95,
         DP_sub_1_root_sub_0_root_sub_104_n94,
         DP_sub_1_root_sub_0_root_sub_104_n93,
         DP_sub_1_root_sub_0_root_sub_104_n92,
         DP_sub_1_root_sub_0_root_sub_104_n91,
         DP_sub_1_root_sub_0_root_sub_104_n90,
         DP_sub_1_root_sub_0_root_sub_104_n88,
         DP_sub_1_root_sub_0_root_sub_104_n87,
         DP_sub_1_root_sub_0_root_sub_104_n85,
         DP_sub_1_root_sub_0_root_sub_104_n83,
         DP_sub_1_root_sub_0_root_sub_104_n81,
         DP_sub_1_root_sub_0_root_sub_104_n79,
         DP_sub_1_root_sub_0_root_sub_104_n78,
         DP_sub_1_root_sub_0_root_sub_104_n77,
         DP_sub_1_root_sub_0_root_sub_104_n75,
         DP_sub_1_root_sub_0_root_sub_104_n74,
         DP_sub_1_root_sub_0_root_sub_104_n73,
         DP_sub_1_root_sub_0_root_sub_104_n72,
         DP_sub_1_root_sub_0_root_sub_104_n71,
         DP_sub_1_root_sub_0_root_sub_104_n70,
         DP_sub_1_root_sub_0_root_sub_104_n69,
         DP_sub_1_root_sub_0_root_sub_104_n68,
         DP_sub_1_root_sub_0_root_sub_104_n67,
         DP_sub_1_root_sub_0_root_sub_104_n66,
         DP_sub_1_root_sub_0_root_sub_104_n65,
         DP_sub_1_root_sub_0_root_sub_104_n64,
         DP_sub_1_root_sub_0_root_sub_104_n63,
         DP_sub_1_root_sub_0_root_sub_104_n62,
         DP_sub_1_root_sub_0_root_sub_104_n61,
         DP_sub_1_root_sub_0_root_sub_104_n60,
         DP_sub_1_root_sub_0_root_sub_104_n59,
         DP_sub_1_root_sub_0_root_sub_104_n58,
         DP_sub_1_root_sub_0_root_sub_104_n57,
         DP_sub_1_root_sub_0_root_sub_104_n56,
         DP_sub_1_root_sub_0_root_sub_104_n55,
         DP_sub_1_root_sub_0_root_sub_104_n54,
         DP_sub_1_root_sub_0_root_sub_104_n51,
         DP_sub_1_root_sub_0_root_sub_104_n50,
         DP_sub_1_root_sub_0_root_sub_104_n49,
         DP_sub_1_root_sub_0_root_sub_104_n48,
         DP_sub_1_root_sub_0_root_sub_104_n46,
         DP_sub_1_root_sub_0_root_sub_104_n45,
         DP_sub_1_root_sub_0_root_sub_104_n44,
         DP_sub_1_root_sub_0_root_sub_104_n43,
         DP_sub_1_root_sub_0_root_sub_104_n42,
         DP_sub_1_root_sub_0_root_sub_104_n41,
         DP_sub_1_root_sub_0_root_sub_104_n40,
         DP_sub_1_root_sub_0_root_sub_104_n39,
         DP_sub_1_root_sub_0_root_sub_104_n38,
         DP_sub_1_root_sub_0_root_sub_104_n37,
         DP_sub_1_root_sub_0_root_sub_104_n36,
         DP_sub_1_root_sub_0_root_sub_104_n35,
         DP_sub_1_root_sub_0_root_sub_104_n34,
         DP_sub_1_root_sub_0_root_sub_104_n33,
         DP_sub_1_root_sub_0_root_sub_104_n32,
         DP_sub_1_root_sub_0_root_sub_104_n31,
         DP_sub_1_root_sub_0_root_sub_104_n30,
         DP_sub_1_root_sub_0_root_sub_104_n29,
         DP_sub_1_root_sub_0_root_sub_104_n28,
         DP_sub_1_root_sub_0_root_sub_104_n27,
         DP_sub_1_root_sub_0_root_sub_104_n26,
         DP_sub_1_root_sub_0_root_sub_104_n24,
         DP_sub_1_root_sub_0_root_sub_104_n22,
         DP_sub_1_root_sub_0_root_sub_104_n21,
         DP_sub_1_root_sub_0_root_sub_104_n20,
         DP_sub_1_root_sub_0_root_sub_104_n19,
         DP_sub_1_root_sub_0_root_sub_104_n18,
         DP_sub_1_root_sub_0_root_sub_104_n17,
         DP_sub_1_root_sub_0_root_sub_104_n16,
         DP_sub_1_root_sub_0_root_sub_104_n15,
         DP_sub_1_root_sub_0_root_sub_104_n14,
         DP_sub_1_root_sub_0_root_sub_104_n11,
         DP_sub_1_root_sub_0_root_sub_104_n10,
         DP_sub_1_root_sub_0_root_sub_104_n7,
         DP_sub_1_root_sub_0_root_sub_104_n6,
         DP_sub_1_root_sub_0_root_sub_104_n5,
         DP_sub_1_root_sub_0_root_sub_104_n4,
         DP_sub_1_root_sub_0_root_sub_104_n3,
         DP_sub_1_root_sub_0_root_sub_104_n1, DP_mult_105_n763,
         DP_mult_105_n762, DP_mult_105_n761, DP_mult_105_n760,
         DP_mult_105_n759, DP_mult_105_n758, DP_mult_105_n757,
         DP_mult_105_n756, DP_mult_105_n755, DP_mult_105_n754,
         DP_mult_105_n753, DP_mult_105_n752, DP_mult_105_n751,
         DP_mult_105_n750, DP_mult_105_n749, DP_mult_105_n748,
         DP_mult_105_n747, DP_mult_105_n746, DP_mult_105_n745,
         DP_mult_105_n744, DP_mult_105_n743, DP_mult_105_n742,
         DP_mult_105_n741, DP_mult_105_n740, DP_mult_105_n739,
         DP_mult_105_n738, DP_mult_105_n737, DP_mult_105_n736,
         DP_mult_105_n735, DP_mult_105_n734, DP_mult_105_n733,
         DP_mult_105_n732, DP_mult_105_n731, DP_mult_105_n730,
         DP_mult_105_n729, DP_mult_105_n728, DP_mult_105_n727,
         DP_mult_105_n726, DP_mult_105_n725, DP_mult_105_n724,
         DP_mult_105_n723, DP_mult_105_n722, DP_mult_105_n721,
         DP_mult_105_n720, DP_mult_105_n719, DP_mult_105_n718,
         DP_mult_105_n717, DP_mult_105_n716, DP_mult_105_n715,
         DP_mult_105_n714, DP_mult_105_n713, DP_mult_105_n712,
         DP_mult_105_n711, DP_mult_105_n710, DP_mult_105_n709,
         DP_mult_105_n708, DP_mult_105_n707, DP_mult_105_n706,
         DP_mult_105_n705, DP_mult_105_n704, DP_mult_105_n703,
         DP_mult_105_n702, DP_mult_105_n701, DP_mult_105_n700,
         DP_mult_105_n699, DP_mult_105_n698, DP_mult_105_n697,
         DP_mult_105_n696, DP_mult_105_n695, DP_mult_105_n694,
         DP_mult_105_n693, DP_mult_105_n692, DP_mult_105_n691,
         DP_mult_105_n690, DP_mult_105_n689, DP_mult_105_n688,
         DP_mult_105_n687, DP_mult_105_n686, DP_mult_105_n685,
         DP_mult_105_n684, DP_mult_105_n683, DP_mult_105_n682,
         DP_mult_105_n681, DP_mult_105_n680, DP_mult_105_n679,
         DP_mult_105_n678, DP_mult_105_n677, DP_mult_105_n676,
         DP_mult_105_n675, DP_mult_105_n674, DP_mult_105_n673,
         DP_mult_105_n672, DP_mult_105_n671, DP_mult_105_n670,
         DP_mult_105_n669, DP_mult_105_n668, DP_mult_105_n667,
         DP_mult_105_n666, DP_mult_105_n665, DP_mult_105_n664,
         DP_mult_105_n663, DP_mult_105_n662, DP_mult_105_n661,
         DP_mult_105_n620, DP_mult_105_n619, DP_mult_105_n618,
         DP_mult_105_n617, DP_mult_105_n616, DP_mult_105_n615,
         DP_mult_105_n614, DP_mult_105_n613, DP_mult_105_n612,
         DP_mult_105_n611, DP_mult_105_n610, DP_mult_105_n609,
         DP_mult_105_n608, DP_mult_105_n607, DP_mult_105_n606,
         DP_mult_105_n605, DP_mult_105_n604, DP_mult_105_n603,
         DP_mult_105_n602, DP_mult_105_n601, DP_mult_105_n600,
         DP_mult_105_n599, DP_mult_105_n598, DP_mult_105_n597,
         DP_mult_105_n596, DP_mult_105_n595, DP_mult_105_n594,
         DP_mult_105_n593, DP_mult_105_n592, DP_mult_105_n591,
         DP_mult_105_n590, DP_mult_105_n589, DP_mult_105_n588,
         DP_mult_105_n587, DP_mult_105_n586, DP_mult_105_n585,
         DP_mult_105_n584, DP_mult_105_n583, DP_mult_105_n582,
         DP_mult_105_n581, DP_mult_105_n580, DP_mult_105_n579,
         DP_mult_105_n577, DP_mult_105_n576, DP_mult_105_n575,
         DP_mult_105_n574, DP_mult_105_n573, DP_mult_105_n572,
         DP_mult_105_n570, DP_mult_105_n569, DP_mult_105_n566,
         DP_mult_105_n565, DP_mult_105_n564, DP_mult_105_n563,
         DP_mult_105_n562, DP_mult_105_n561, DP_mult_105_n560,
         DP_mult_105_n559, DP_mult_105_n558, DP_mult_105_n557,
         DP_mult_105_n556, DP_mult_105_n555, DP_mult_105_n554,
         DP_mult_105_n553, DP_mult_105_n552, DP_mult_105_n551,
         DP_mult_105_n550, DP_mult_105_n549, DP_mult_105_n548,
         DP_mult_105_n547, DP_mult_105_n546, DP_mult_105_n545,
         DP_mult_105_n544, DP_mult_105_n543, DP_mult_105_n542,
         DP_mult_105_n541, DP_mult_105_n540, DP_mult_105_n539,
         DP_mult_105_n538, DP_mult_105_n537, DP_mult_105_n536,
         DP_mult_105_n535, DP_mult_105_n534, DP_mult_105_n533,
         DP_mult_105_n532, DP_mult_105_n531, DP_mult_105_n530,
         DP_mult_105_n529, DP_mult_105_n528, DP_mult_105_n527,
         DP_mult_105_n526, DP_mult_105_n525, DP_mult_105_n524,
         DP_mult_105_n523, DP_mult_105_n522, DP_mult_105_n521,
         DP_mult_105_n520, DP_mult_105_n519, DP_mult_105_n518,
         DP_mult_105_n517, DP_mult_105_n516, DP_mult_105_n515,
         DP_mult_105_n514, DP_mult_105_n513, DP_mult_105_n512,
         DP_mult_105_n511, DP_mult_105_n510, DP_mult_105_n509,
         DP_mult_105_n508, DP_mult_105_n507, DP_mult_105_n506,
         DP_mult_105_n505, DP_mult_105_n504, DP_mult_105_n503,
         DP_mult_105_n502, DP_mult_105_n501, DP_mult_105_n500,
         DP_mult_105_n499, DP_mult_105_n498, DP_mult_105_n497,
         DP_mult_105_n496, DP_mult_105_n495, DP_mult_105_n494,
         DP_mult_105_n493, DP_mult_105_n492, DP_mult_105_n491,
         DP_mult_105_n490, DP_mult_105_n489, DP_mult_105_n488,
         DP_mult_105_n487, DP_mult_105_n486, DP_mult_105_n485,
         DP_mult_105_n484, DP_mult_105_n483, DP_mult_105_n482,
         DP_mult_105_n481, DP_mult_105_n480, DP_mult_105_n479,
         DP_mult_105_n478, DP_mult_105_n477, DP_mult_105_n476,
         DP_mult_105_n475, DP_mult_105_n474, DP_mult_105_n473,
         DP_mult_105_n472, DP_mult_105_n471, DP_mult_105_n469,
         DP_mult_105_n467, DP_mult_105_n466, DP_mult_105_n465,
         DP_mult_105_n464, DP_mult_105_n463, DP_mult_105_n462,
         DP_mult_105_n461, DP_mult_105_n460, DP_mult_105_n459,
         DP_mult_105_n458, DP_mult_105_n457, DP_mult_105_n456,
         DP_mult_105_n454, DP_mult_105_n453, DP_mult_105_n452,
         DP_mult_105_n451, DP_mult_105_n450, DP_mult_105_n449,
         DP_mult_105_n448, DP_mult_105_n447, DP_mult_105_n446,
         DP_mult_105_n445, DP_mult_105_n444, DP_mult_105_n443,
         DP_mult_105_n441, DP_mult_105_n440, DP_mult_105_n439,
         DP_mult_105_n438, DP_mult_105_n437, DP_mult_105_n436,
         DP_mult_105_n435, DP_mult_105_n434, DP_mult_105_n433,
         DP_mult_105_n432, DP_mult_105_n431, DP_mult_105_n430,
         DP_mult_105_n428, DP_mult_105_n427, DP_mult_105_n426,
         DP_mult_105_n425, DP_mult_105_n424, DP_mult_105_n423,
         DP_mult_105_n422, DP_mult_105_n421, DP_mult_105_n420,
         DP_mult_105_n419, DP_mult_105_n418, DP_mult_105_n417,
         DP_mult_105_n415, DP_mult_105_n414, DP_mult_105_n413,
         DP_mult_105_n412, DP_mult_105_n411, DP_mult_105_n410,
         DP_mult_105_n409, DP_mult_105_n408, DP_mult_105_n407,
         DP_mult_105_n406, DP_mult_105_n405, DP_mult_105_n404,
         DP_mult_105_n403, DP_mult_105_n402, DP_mult_105_n401,
         DP_mult_105_n400, DP_mult_105_n399, DP_mult_105_n398,
         DP_mult_105_n397, DP_mult_105_n396, DP_mult_105_n395,
         DP_mult_105_n394, DP_mult_105_n393, DP_mult_105_n392,
         DP_mult_105_n391, DP_mult_105_n390, DP_mult_105_n389,
         DP_mult_105_n388, DP_mult_105_n387, DP_mult_105_n386,
         DP_mult_105_n385, DP_mult_105_n384, DP_mult_105_n383,
         DP_mult_105_n382, DP_mult_105_n381, DP_mult_105_n380,
         DP_mult_105_n379, DP_mult_105_n378, DP_mult_105_n377,
         DP_mult_105_n376, DP_mult_105_n375, DP_mult_105_n374,
         DP_mult_105_n373, DP_mult_105_n372, DP_mult_105_n371,
         DP_mult_105_n370, DP_mult_105_n369, DP_mult_105_n368,
         DP_mult_105_n367, DP_mult_105_n366, DP_mult_105_n365,
         DP_mult_105_n364, DP_mult_105_n363, DP_mult_105_n362,
         DP_mult_105_n361, DP_mult_105_n360, DP_mult_105_n359,
         DP_mult_105_n358, DP_mult_105_n357, DP_mult_105_n356,
         DP_mult_105_n355, DP_mult_105_n354, DP_mult_105_n353,
         DP_mult_105_n352, DP_mult_105_n351, DP_mult_105_n350,
         DP_mult_105_n349, DP_mult_105_n348, DP_mult_105_n347,
         DP_mult_105_n346, DP_mult_105_n345, DP_mult_105_n344,
         DP_mult_105_n343, DP_mult_105_n342, DP_mult_105_n341,
         DP_mult_105_n340, DP_mult_105_n339, DP_mult_105_n338,
         DP_mult_105_n337, DP_mult_105_n336, DP_mult_105_n335,
         DP_mult_105_n334, DP_mult_105_n333, DP_mult_105_n332,
         DP_mult_105_n331, DP_mult_105_n330, DP_mult_105_n329,
         DP_mult_105_n328, DP_mult_105_n327, DP_mult_105_n326,
         DP_mult_105_n325, DP_mult_105_n324, DP_mult_105_n323,
         DP_mult_105_n322, DP_mult_105_n321, DP_mult_105_n320,
         DP_mult_105_n319, DP_mult_105_n318, DP_mult_105_n317,
         DP_mult_105_n316, DP_mult_105_n315, DP_mult_105_n314,
         DP_mult_105_n313, DP_mult_105_n312, DP_mult_105_n311,
         DP_mult_105_n310, DP_mult_105_n309, DP_mult_105_n308,
         DP_mult_105_n307, DP_mult_105_n306, DP_mult_105_n305,
         DP_mult_105_n304, DP_mult_105_n303, DP_mult_105_n302,
         DP_mult_105_n301, DP_mult_105_n300, DP_mult_105_n299,
         DP_mult_105_n298, DP_mult_105_n297, DP_mult_105_n296,
         DP_mult_105_n295, DP_mult_105_n294, DP_mult_105_n293,
         DP_mult_105_n292, DP_mult_105_n291, DP_mult_105_n290,
         DP_mult_105_n289, DP_mult_105_n288, DP_mult_105_n287,
         DP_mult_105_n286, DP_mult_105_n285, DP_mult_105_n284,
         DP_mult_105_n283, DP_mult_105_n282, DP_mult_105_n281,
         DP_mult_105_n280, DP_mult_105_n279, DP_mult_105_n278,
         DP_mult_105_n273, DP_mult_105_n260, DP_mult_105_n259,
         DP_mult_105_n258, DP_mult_105_n257, DP_mult_105_n256,
         DP_mult_105_n255, DP_mult_105_n254, DP_mult_105_n253,
         DP_mult_105_n252, DP_mult_105_n251, DP_mult_105_n250,
         DP_mult_105_n249, DP_mult_105_n248, DP_mult_105_n247,
         DP_mult_105_n242, DP_mult_105_n233, DP_mult_105_n232,
         DP_mult_105_n231, DP_mult_105_n230, DP_mult_105_n229,
         DP_mult_105_n228, DP_mult_105_n227, DP_mult_105_n226,
         DP_mult_105_n225, DP_mult_105_n224, DP_mult_105_n223,
         DP_mult_105_n222, DP_mult_105_n221, DP_mult_105_n220,
         DP_mult_105_n219, DP_mult_105_n218, DP_mult_105_n216,
         DP_mult_105_n215, DP_mult_105_n214, DP_mult_105_n213,
         DP_mult_105_n212, DP_mult_105_n211, DP_mult_105_n209,
         DP_mult_105_n208, DP_mult_105_n207, DP_mult_105_n206,
         DP_mult_105_n203, DP_mult_105_n202, DP_mult_105_n201,
         DP_mult_105_n200, DP_mult_105_n199, DP_mult_105_n198,
         DP_mult_105_n197, DP_mult_105_n196, DP_mult_105_n195,
         DP_mult_105_n194, DP_mult_105_n193, DP_mult_105_n192,
         DP_mult_105_n191, DP_mult_105_n190, DP_mult_105_n185,
         DP_mult_105_n184, DP_mult_105_n183, DP_mult_105_n181,
         DP_mult_105_n179, DP_mult_105_n178, DP_mult_105_n177,
         DP_mult_105_n176, DP_mult_105_n175, DP_mult_105_n174,
         DP_mult_105_n172, DP_mult_105_n170, DP_mult_105_n169,
         DP_mult_105_n168, DP_mult_105_n167, DP_mult_105_n166,
         DP_mult_105_n165, DP_mult_105_n163, DP_mult_105_n161,
         DP_mult_105_n160, DP_mult_105_n159, DP_mult_105_n158,
         DP_mult_105_n157, DP_mult_105_n156, DP_mult_105_n155,
         DP_mult_105_n154, DP_mult_105_n152, DP_mult_105_n150,
         DP_mult_105_n149, DP_mult_105_n148, DP_mult_105_n147,
         DP_mult_105_n146, DP_mult_105_n145, DP_mult_105_n143,
         DP_mult_105_n141, DP_mult_105_n139, DP_mult_105_n137,
         DP_mult_105_n136, DP_mult_105_n135, DP_mult_105_n134,
         DP_mult_105_n133, DP_mult_105_n132, DP_mult_105_n131,
         DP_mult_105_n130, DP_mult_105_n129, DP_mult_105_n128,
         DP_mult_105_n127, DP_mult_105_n126, DP_mult_105_n123,
         DP_mult_105_n119, DP_mult_105_n118, DP_mult_105_n117,
         DP_mult_105_n116, DP_mult_105_n115, DP_mult_105_n114,
         DP_mult_105_n111, DP_mult_105_n109, DP_mult_105_n105,
         DP_mult_105_n103, DP_mult_105_n93, DP_mult_105_n87, DP_mult_105_n77,
         DP_mult_105_n73, DP_mult_105_n69, DP_mult_105_n57, DP_mult_105_n48,
         DP_mult_105_n40, DP_mult_105_n35, DP_mult_105_n30, DP_mult_105_n26,
         DP_mult_105_n24, DP_mult_105_n14, DP_mult_105_n10, DP_mult_105_n8,
         CU_n1, CU_n12, CU_n11, CU_n10, CU_n9, CU_n8, CU_n6, CU_n5, CU_n4,
         CU_n3, CU_N20, CU_presentState_0_, CU_presentState_1_,
         CU_presentState_2_;
  wire   [35:0] DP_b_int;
  wire   [23:0] DP_a_int;
  wire   [0:1] CU_nextState;

  OAI21_X1 DP_U48 ( .B1(DP_n20), .B2(DP_n35), .A(DP_n19), .ZN(DP_y_out_10_) );
  INV_X1 DP_U47 ( .A(DP_y_10_), .ZN(DP_n35) );
  OAI21_X1 DP_U46 ( .B1(DP_n20), .B2(DP_n33), .A(DP_n18), .ZN(DP_y_out_9_) );
  INV_X1 DP_U45 ( .A(DP_y_9_), .ZN(DP_n33) );
  OAI21_X1 DP_U44 ( .B1(DP_n17), .B2(DP_n32), .A(DP_n19), .ZN(DP_y_out_8_) );
  INV_X1 DP_U43 ( .A(DP_y_8_), .ZN(DP_n32) );
  OAI21_X1 DP_U42 ( .B1(DP_n17), .B2(DP_n31), .A(DP_n18), .ZN(DP_y_out_7_) );
  INV_X1 DP_U41 ( .A(DP_y_7_), .ZN(DP_n31) );
  OAI21_X1 DP_U40 ( .B1(DP_n17), .B2(DP_n30), .A(DP_n34), .ZN(DP_y_out_6_) );
  INV_X1 DP_U39 ( .A(DP_y_6_), .ZN(DP_n30) );
  OAI21_X1 DP_U38 ( .B1(DP_n17), .B2(DP_n29), .A(DP_n4), .ZN(DP_y_out_5_) );
  INV_X1 DP_U37 ( .A(DP_y_5_), .ZN(DP_n29) );
  OAI21_X1 DP_U36 ( .B1(DP_n20), .B2(DP_n28), .A(DP_n34), .ZN(DP_y_out_4_) );
  INV_X1 DP_U35 ( .A(DP_y_4_), .ZN(DP_n28) );
  OAI21_X1 DP_U34 ( .B1(DP_n20), .B2(DP_n27), .A(DP_n4), .ZN(DP_y_out_3_) );
  INV_X1 DP_U33 ( .A(DP_y_3_), .ZN(DP_n27) );
  OAI21_X1 DP_U32 ( .B1(DP_n17), .B2(DP_n26), .A(DP_n34), .ZN(DP_y_out_2_) );
  INV_X1 DP_U31 ( .A(DP_y_2_), .ZN(DP_n26) );
  OAI21_X1 DP_U30 ( .B1(DP_n20), .B2(DP_n25), .A(DP_n4), .ZN(DP_y_out_1_) );
  INV_X1 DP_U29 ( .A(DP_y_1_), .ZN(DP_n25) );
  NAND2_X1 DP_U28 ( .A1(DP_n19), .A2(DP_n23), .ZN(DP_y_out_0_) );
  INV_X1 DP_U27 ( .A(DP_y_out_11_), .ZN(DP_n22) );
  NAND2_X1 DP_U26 ( .A1(DP_n24), .A2(DP_y_0_), .ZN(DP_n23) );
  INV_X1 DP_U25 ( .A(DP_y_11_), .ZN(DP_n21) );
  NAND2_X1 DP_U24 ( .A1(DP_n21), .A2(DP_y_out_11_), .ZN(DP_n24) );
  INV_X1 DP_U23 ( .A(DP_n24), .ZN(DP_n20) );
  NAND2_X1 DP_U22 ( .A1(DP_n22), .A2(DP_y_11_), .ZN(DP_n34) );
  NAND2_X1 DP_U21 ( .A1(DP_n22), .A2(DP_y_11_), .ZN(DP_n18) );
  NAND2_X1 DP_U20 ( .A1(DP_n22), .A2(DP_y_11_), .ZN(DP_n19) );
  INV_X1 DP_U19 ( .A(DP_n24), .ZN(DP_n17) );
  CLKBUF_X1 DP_U18 ( .A(DP_sw1_3_), .Z(DP_n16) );
  INV_X1 DP_U17 ( .A(DP_n22), .ZN(DP_n15) );
  CLKBUF_X1 DP_U16 ( .A(DP_sw1_2_), .Z(DP_n14) );
  CLKBUF_X1 DP_U15 ( .A(DP_w_10_), .Z(DP_n13) );
  CLKBUF_X1 DP_U14 ( .A(DP_w_12_), .Z(DP_n12) );
  CLKBUF_X1 DP_U13 ( .A(DP_w_11_), .Z(DP_n11) );
  CLKBUF_X1 DP_U12 ( .A(DP_sw1_6_), .Z(DP_n10) );
  CLKBUF_X1 DP_U11 ( .A(DP_w_9_), .Z(DP_n9) );
  CLKBUF_X1 DP_U10 ( .A(DP_sw1_7_), .Z(DP_n8) );
  CLKBUF_X1 DP_U9 ( .A(DP_sw1_10_), .Z(DP_n7) );
  CLKBUF_X1 DP_U8 ( .A(DP_sw1_11_), .Z(DP_n6) );
  CLKBUF_X1 DP_U7 ( .A(DP_sw1_4_), .Z(DP_n5) );
  NAND2_X1 DP_U6 ( .A1(DP_n22), .A2(DP_y_11_), .ZN(DP_n4) );
  INV_X2 DP_U5 ( .A(DP_n2), .ZN(DP_n3) );
  INV_X1 DP_U4 ( .A(DP_sw1_0_), .ZN(DP_n2) );
  CLKBUF_X1 DP_U3 ( .A(DP_sw0_1_), .Z(DP_n1) );
  NAND2_X1 DP_reg_in_U28 ( .A1(dIn[10]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n11) );
  OAI21_X1 DP_reg_in_U27 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n23), .A(
        DP_reg_in_n11), .ZN(DP_reg_in_n35) );
  NAND2_X1 DP_reg_in_U26 ( .A1(dIn[9]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n10)
         );
  OAI21_X1 DP_reg_in_U25 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n22), .A(
        DP_reg_in_n10), .ZN(DP_reg_in_n34) );
  NAND2_X1 DP_reg_in_U24 ( .A1(dIn[8]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n9)
         );
  OAI21_X1 DP_reg_in_U23 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n21), .A(
        DP_reg_in_n9), .ZN(DP_reg_in_n33) );
  NAND2_X1 DP_reg_in_U22 ( .A1(dIn[7]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n8)
         );
  OAI21_X1 DP_reg_in_U21 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n20), .A(
        DP_reg_in_n8), .ZN(DP_reg_in_n32) );
  NAND2_X1 DP_reg_in_U20 ( .A1(dIn[6]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n7)
         );
  OAI21_X1 DP_reg_in_U19 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n19), .A(
        DP_reg_in_n7), .ZN(DP_reg_in_n31) );
  NAND2_X1 DP_reg_in_U18 ( .A1(dIn[5]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n6)
         );
  OAI21_X1 DP_reg_in_U17 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n18), .A(
        DP_reg_in_n6), .ZN(DP_reg_in_n30) );
  NAND2_X1 DP_reg_in_U16 ( .A1(dIn[4]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n5)
         );
  OAI21_X1 DP_reg_in_U15 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n17), .A(
        DP_reg_in_n5), .ZN(DP_reg_in_n29) );
  NAND2_X1 DP_reg_in_U14 ( .A1(dIn[3]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n4)
         );
  OAI21_X1 DP_reg_in_U13 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n16), .A(
        DP_reg_in_n4), .ZN(DP_reg_in_n28) );
  NAND2_X1 DP_reg_in_U12 ( .A1(dIn[2]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n3)
         );
  OAI21_X1 DP_reg_in_U11 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n15), .A(
        DP_reg_in_n3), .ZN(DP_reg_in_n27) );
  NAND2_X1 DP_reg_in_U10 ( .A1(dIn[1]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n2)
         );
  OAI21_X1 DP_reg_in_U9 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n14), .A(
        DP_reg_in_n2), .ZN(DP_reg_in_n26) );
  NAND2_X1 DP_reg_in_U8 ( .A1(DP_reg_in_n39), .A2(dIn[0]), .ZN(DP_reg_in_n1)
         );
  OAI21_X1 DP_reg_in_U7 ( .B1(DP_reg_in_n39), .B2(DP_reg_in_n13), .A(
        DP_reg_in_n1), .ZN(DP_reg_in_n25) );
  NAND2_X1 DP_reg_in_U6 ( .A1(dIn[11]), .A2(DP_reg_in_n38), .ZN(DP_reg_in_n12)
         );
  OAI21_X1 DP_reg_in_U5 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n24), .A(
        DP_reg_in_n12), .ZN(DP_reg_in_n37) );
  INV_X1 DP_reg_in_U4 ( .A(regs_clr_int), .ZN(DP_reg_in_n36) );
  BUF_X1 DP_reg_in_U3 ( .A(vIn), .Z(DP_reg_in_n39) );
  BUF_X1 DP_reg_in_U2 ( .A(vIn), .Z(DP_reg_in_n38) );
  DFFR_X1 DP_reg_in_Q_reg_0_ ( .D(DP_reg_in_n25), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_0_), .QN(DP_reg_in_n13) );
  DFFR_X1 DP_reg_in_Q_reg_1_ ( .D(DP_reg_in_n26), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_1_), .QN(DP_reg_in_n14) );
  DFFR_X1 DP_reg_in_Q_reg_2_ ( .D(DP_reg_in_n27), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_2_), .QN(DP_reg_in_n15) );
  DFFR_X1 DP_reg_in_Q_reg_3_ ( .D(DP_reg_in_n28), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_3_), .QN(DP_reg_in_n16) );
  DFFR_X1 DP_reg_in_Q_reg_4_ ( .D(DP_reg_in_n29), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_4_), .QN(DP_reg_in_n17) );
  DFFR_X1 DP_reg_in_Q_reg_5_ ( .D(DP_reg_in_n30), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_5_), .QN(DP_reg_in_n18) );
  DFFR_X1 DP_reg_in_Q_reg_6_ ( .D(DP_reg_in_n31), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_6_), .QN(DP_reg_in_n19) );
  DFFR_X1 DP_reg_in_Q_reg_7_ ( .D(DP_reg_in_n32), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_7_), .QN(DP_reg_in_n20) );
  DFFR_X1 DP_reg_in_Q_reg_8_ ( .D(DP_reg_in_n33), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_8_), .QN(DP_reg_in_n21) );
  DFFR_X1 DP_reg_in_Q_reg_9_ ( .D(DP_reg_in_n34), .CK(clk), .RN(DP_reg_in_n36), 
        .Q(DP_x_9_), .QN(DP_reg_in_n22) );
  DFFR_X1 DP_reg_in_Q_reg_10_ ( .D(DP_reg_in_n35), .CK(clk), .RN(DP_reg_in_n36), .Q(DP_x_10_), .QN(DP_reg_in_n23) );
  DFFR_X1 DP_reg_in_Q_reg_11_ ( .D(DP_reg_in_n37), .CK(clk), .RN(DP_reg_in_n36), .Q(DP_x_11_), .QN(DP_reg_in_n24) );
  NAND2_X1 DP_reg_a_i_1_U28 ( .A1(a[22]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n66) );
  OAI21_X1 DP_reg_a_i_1_U27 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n54), 
        .A(DP_reg_a_i_1_n66), .ZN(DP_reg_a_i_1_n42) );
  NAND2_X1 DP_reg_a_i_1_U26 ( .A1(a[21]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n67) );
  OAI21_X1 DP_reg_a_i_1_U25 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n55), 
        .A(DP_reg_a_i_1_n67), .ZN(DP_reg_a_i_1_n43) );
  NAND2_X1 DP_reg_a_i_1_U24 ( .A1(a[20]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n68) );
  OAI21_X1 DP_reg_a_i_1_U23 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n56), 
        .A(DP_reg_a_i_1_n68), .ZN(DP_reg_a_i_1_n44) );
  NAND2_X1 DP_reg_a_i_1_U22 ( .A1(a[19]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n69) );
  OAI21_X1 DP_reg_a_i_1_U21 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n57), 
        .A(DP_reg_a_i_1_n69), .ZN(DP_reg_a_i_1_n45) );
  NAND2_X1 DP_reg_a_i_1_U20 ( .A1(a[18]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n70) );
  OAI21_X1 DP_reg_a_i_1_U19 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n58), 
        .A(DP_reg_a_i_1_n70), .ZN(DP_reg_a_i_1_n46) );
  NAND2_X1 DP_reg_a_i_1_U18 ( .A1(a[17]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n71) );
  OAI21_X1 DP_reg_a_i_1_U17 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n59), 
        .A(DP_reg_a_i_1_n71), .ZN(DP_reg_a_i_1_n47) );
  NAND2_X1 DP_reg_a_i_1_U16 ( .A1(a[16]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n72) );
  OAI21_X1 DP_reg_a_i_1_U15 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n60), 
        .A(DP_reg_a_i_1_n72), .ZN(DP_reg_a_i_1_n48) );
  NAND2_X1 DP_reg_a_i_1_U14 ( .A1(a[15]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n73) );
  OAI21_X1 DP_reg_a_i_1_U13 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n61), 
        .A(DP_reg_a_i_1_n73), .ZN(DP_reg_a_i_1_n49) );
  NAND2_X1 DP_reg_a_i_1_U12 ( .A1(a[14]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n74) );
  OAI21_X1 DP_reg_a_i_1_U11 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n62), 
        .A(DP_reg_a_i_1_n74), .ZN(DP_reg_a_i_1_n50) );
  NAND2_X1 DP_reg_a_i_1_U10 ( .A1(a[13]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n75) );
  OAI21_X1 DP_reg_a_i_1_U9 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n63), .A(
        DP_reg_a_i_1_n75), .ZN(DP_reg_a_i_1_n51) );
  NAND2_X1 DP_reg_a_i_1_U8 ( .A1(DP_reg_a_i_1_n39), .A2(a[12]), .ZN(
        DP_reg_a_i_1_n76) );
  OAI21_X1 DP_reg_a_i_1_U7 ( .B1(DP_reg_a_i_1_n39), .B2(DP_reg_a_i_1_n64), .A(
        DP_reg_a_i_1_n76), .ZN(DP_reg_a_i_1_n52) );
  NAND2_X1 DP_reg_a_i_1_U6 ( .A1(a[23]), .A2(DP_reg_a_i_1_n38), .ZN(
        DP_reg_a_i_1_n65) );
  OAI21_X1 DP_reg_a_i_1_U5 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n53), .A(
        DP_reg_a_i_1_n65), .ZN(DP_reg_a_i_1_n40) );
  INV_X1 DP_reg_a_i_1_U4 ( .A(regs_clr_int), .ZN(DP_reg_a_i_1_n41) );
  BUF_X1 DP_reg_a_i_1_U3 ( .A(vIn), .Z(DP_reg_a_i_1_n39) );
  BUF_X1 DP_reg_a_i_1_U2 ( .A(vIn), .Z(DP_reg_a_i_1_n38) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_0_ ( .D(DP_reg_a_i_1_n52), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[11]), .QN(DP_reg_a_i_1_n64) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_1_ ( .D(DP_reg_a_i_1_n51), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[10]), .QN(DP_reg_a_i_1_n63) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_2_ ( .D(DP_reg_a_i_1_n50), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[9]), .QN(DP_reg_a_i_1_n62) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_3_ ( .D(DP_reg_a_i_1_n49), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[8]), .QN(DP_reg_a_i_1_n61) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_4_ ( .D(DP_reg_a_i_1_n48), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[7]), .QN(DP_reg_a_i_1_n60) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_5_ ( .D(DP_reg_a_i_1_n47), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[6]), .QN(DP_reg_a_i_1_n59) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_6_ ( .D(DP_reg_a_i_1_n46), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[5]), .QN(DP_reg_a_i_1_n58) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_7_ ( .D(DP_reg_a_i_1_n45), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[4]), .QN(DP_reg_a_i_1_n57) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_8_ ( .D(DP_reg_a_i_1_n44), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[3]), .QN(DP_reg_a_i_1_n56) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_9_ ( .D(DP_reg_a_i_1_n43), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[2]), .QN(DP_reg_a_i_1_n55) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_10_ ( .D(DP_reg_a_i_1_n42), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[1]), .QN(DP_reg_a_i_1_n54) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_11_ ( .D(DP_reg_a_i_1_n40), .CK(clk), .RN(
        DP_reg_a_i_1_n41), .Q(DP_a_int[0]), .QN(DP_reg_a_i_1_n53) );
  OAI21_X1 DP_reg_a_i_2_U44 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n73), 
        .A(DP_reg_a_i_2_n85), .ZN(DP_reg_a_i_2_n61) );
  OAI21_X1 DP_reg_a_i_2_U43 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n77), 
        .A(DP_reg_a_i_2_n89), .ZN(DP_reg_a_i_2_n65) );
  OAI21_X1 DP_reg_a_i_2_U42 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n75), 
        .A(DP_reg_a_i_2_n87), .ZN(DP_reg_a_i_2_n63) );
  NAND2_X1 DP_reg_a_i_2_U41 ( .A1(a[10]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n82) );
  OAI21_X1 DP_reg_a_i_2_U40 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n70), 
        .A(DP_reg_a_i_2_n82), .ZN(DP_reg_a_i_2_n58) );
  NAND2_X1 DP_reg_a_i_2_U39 ( .A1(a[9]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n83) );
  OAI21_X1 DP_reg_a_i_2_U38 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n71), 
        .A(DP_reg_a_i_2_n83), .ZN(DP_reg_a_i_2_n59) );
  NAND2_X1 DP_reg_a_i_2_U37 ( .A1(a[8]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n84) );
  OAI21_X1 DP_reg_a_i_2_U36 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n72), 
        .A(DP_reg_a_i_2_n84), .ZN(DP_reg_a_i_2_n60) );
  NAND2_X1 DP_reg_a_i_2_U35 ( .A1(a[6]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n86) );
  OAI21_X1 DP_reg_a_i_2_U34 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n74), 
        .A(DP_reg_a_i_2_n86), .ZN(DP_reg_a_i_2_n62) );
  NAND2_X1 DP_reg_a_i_2_U33 ( .A1(a[4]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n88) );
  OAI21_X1 DP_reg_a_i_2_U32 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n76), 
        .A(DP_reg_a_i_2_n88), .ZN(DP_reg_a_i_2_n64) );
  NAND2_X1 DP_reg_a_i_2_U31 ( .A1(a[2]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n90) );
  OAI21_X1 DP_reg_a_i_2_U30 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n78), 
        .A(DP_reg_a_i_2_n90), .ZN(DP_reg_a_i_2_n66) );
  NAND2_X1 DP_reg_a_i_2_U29 ( .A1(a[1]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n91) );
  OAI21_X1 DP_reg_a_i_2_U28 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n79), 
        .A(DP_reg_a_i_2_n91), .ZN(DP_reg_a_i_2_n67) );
  NAND2_X1 DP_reg_a_i_2_U27 ( .A1(DP_reg_a_i_2_n55), .A2(a[0]), .ZN(
        DP_reg_a_i_2_n92) );
  OAI21_X1 DP_reg_a_i_2_U26 ( .B1(DP_reg_a_i_2_n55), .B2(DP_reg_a_i_2_n80), 
        .A(DP_reg_a_i_2_n92), .ZN(DP_reg_a_i_2_n68) );
  NAND2_X1 DP_reg_a_i_2_U25 ( .A1(a[11]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n81) );
  OAI21_X1 DP_reg_a_i_2_U24 ( .B1(DP_reg_a_i_2_n54), .B2(DP_reg_a_i_2_n69), 
        .A(DP_reg_a_i_2_n81), .ZN(DP_reg_a_i_2_n56) );
  NAND2_X1 DP_reg_a_i_2_U23 ( .A1(a[7]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n85) );
  NAND2_X1 DP_reg_a_i_2_U22 ( .A1(a[5]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n87) );
  NAND2_X1 DP_reg_a_i_2_U21 ( .A1(a[3]), .A2(DP_reg_a_i_2_n54), .ZN(
        DP_reg_a_i_2_n89) );
  INV_X1 DP_reg_a_i_2_U20 ( .A(regs_clr_int), .ZN(DP_reg_a_i_2_n57) );
  BUF_X1 DP_reg_a_i_2_U19 ( .A(vIn), .Z(DP_reg_a_i_2_n55) );
  BUF_X1 DP_reg_a_i_2_U18 ( .A(vIn), .Z(DP_reg_a_i_2_n54) );
  SDFFR_X1 DP_reg_a_i_2_Q_reg_0_ ( .D(1'b0), .SI(DP_reg_a_i_2_n68), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_a_i_2_n57), .Q(DP_a_int[23]), .QN(
        DP_reg_a_i_2_n80) );
  SDFFR_X1 DP_reg_a_i_2_Q_reg_6_ ( .D(1'b0), .SI(DP_reg_a_i_2_n62), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_a_i_2_n57), .Q(DP_a_int[17]), .QN(
        DP_reg_a_i_2_n74) );
  SDFFR_X1 DP_reg_a_i_2_Q_reg_5_ ( .D(1'b0), .SI(DP_reg_a_i_2_n63), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_a_i_2_n57), .Q(DP_a_int[18]), .QN(
        DP_reg_a_i_2_n75) );
  SDFFR_X1 DP_reg_a_i_2_Q_reg_9_ ( .D(1'b0), .SI(DP_reg_a_i_2_n59), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_a_i_2_n57), .Q(DP_a_int[14]), .QN(
        DP_reg_a_i_2_n71) );
  SDFFR_X1 DP_reg_a_i_2_Q_reg_7_ ( .D(1'b0), .SI(DP_reg_a_i_2_n61), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_a_i_2_n57), .Q(DP_a_int[16]), .QN(
        DP_reg_a_i_2_n73) );
  SDFFR_X1 DP_reg_a_i_2_Q_reg_3_ ( .D(1'b0), .SI(DP_reg_a_i_2_n65), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_a_i_2_n57), .Q(DP_a_int[20]), .QN(
        DP_reg_a_i_2_n77) );
  SDFFR_X1 DP_reg_a_i_2_Q_reg_4_ ( .D(1'b0), .SI(DP_reg_a_i_2_n64), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_a_i_2_n57), .Q(DP_a_int[19]), .QN(
        DP_reg_a_i_2_n76) );
  SDFFR_X1 DP_reg_a_i_2_Q_reg_1_ ( .D(1'b0), .SI(DP_reg_a_i_2_n67), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_a_i_2_n57), .Q(DP_a_int[22]), .QN(
        DP_reg_a_i_2_n79) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_2_ ( .D(DP_reg_a_i_2_n66), .CK(clk), .RN(
        DP_reg_a_i_2_n57), .Q(DP_a_int[21]), .QN(DP_reg_a_i_2_n78) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_8_ ( .D(DP_reg_a_i_2_n60), .CK(clk), .RN(
        DP_reg_a_i_2_n57), .Q(DP_a_int[15]), .QN(DP_reg_a_i_2_n72) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_10_ ( .D(DP_reg_a_i_2_n58), .CK(clk), .RN(
        DP_reg_a_i_2_n57), .Q(DP_a_int[13]), .QN(DP_reg_a_i_2_n70) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_11_ ( .D(DP_reg_a_i_2_n56), .CK(clk), .RN(
        DP_reg_a_i_2_n57), .Q(DP_a_int[12]), .QN(DP_reg_a_i_2_n69) );
  NAND2_X1 DP_reg_b_i_0_U28 ( .A1(b[34]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n66) );
  OAI21_X1 DP_reg_b_i_0_U27 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n54), 
        .A(DP_reg_b_i_0_n66), .ZN(DP_reg_b_i_0_n42) );
  NAND2_X1 DP_reg_b_i_0_U26 ( .A1(b[33]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n67) );
  OAI21_X1 DP_reg_b_i_0_U25 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n55), 
        .A(DP_reg_b_i_0_n67), .ZN(DP_reg_b_i_0_n43) );
  NAND2_X1 DP_reg_b_i_0_U24 ( .A1(b[32]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n68) );
  OAI21_X1 DP_reg_b_i_0_U23 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n56), 
        .A(DP_reg_b_i_0_n68), .ZN(DP_reg_b_i_0_n44) );
  NAND2_X1 DP_reg_b_i_0_U22 ( .A1(b[31]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n69) );
  OAI21_X1 DP_reg_b_i_0_U21 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n57), 
        .A(DP_reg_b_i_0_n69), .ZN(DP_reg_b_i_0_n45) );
  NAND2_X1 DP_reg_b_i_0_U20 ( .A1(b[30]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n70) );
  OAI21_X1 DP_reg_b_i_0_U19 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n58), 
        .A(DP_reg_b_i_0_n70), .ZN(DP_reg_b_i_0_n46) );
  NAND2_X1 DP_reg_b_i_0_U18 ( .A1(b[29]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n71) );
  OAI21_X1 DP_reg_b_i_0_U17 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n59), 
        .A(DP_reg_b_i_0_n71), .ZN(DP_reg_b_i_0_n47) );
  NAND2_X1 DP_reg_b_i_0_U16 ( .A1(b[28]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n72) );
  OAI21_X1 DP_reg_b_i_0_U15 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n60), 
        .A(DP_reg_b_i_0_n72), .ZN(DP_reg_b_i_0_n48) );
  NAND2_X1 DP_reg_b_i_0_U14 ( .A1(b[27]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n73) );
  OAI21_X1 DP_reg_b_i_0_U13 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n61), 
        .A(DP_reg_b_i_0_n73), .ZN(DP_reg_b_i_0_n49) );
  NAND2_X1 DP_reg_b_i_0_U12 ( .A1(b[26]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n74) );
  OAI21_X1 DP_reg_b_i_0_U11 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n62), 
        .A(DP_reg_b_i_0_n74), .ZN(DP_reg_b_i_0_n50) );
  NAND2_X1 DP_reg_b_i_0_U10 ( .A1(b[25]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n75) );
  OAI21_X1 DP_reg_b_i_0_U9 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n63), .A(
        DP_reg_b_i_0_n75), .ZN(DP_reg_b_i_0_n51) );
  NAND2_X1 DP_reg_b_i_0_U8 ( .A1(DP_reg_b_i_0_n39), .A2(b[24]), .ZN(
        DP_reg_b_i_0_n76) );
  OAI21_X1 DP_reg_b_i_0_U7 ( .B1(DP_reg_b_i_0_n39), .B2(DP_reg_b_i_0_n64), .A(
        DP_reg_b_i_0_n76), .ZN(DP_reg_b_i_0_n52) );
  NAND2_X1 DP_reg_b_i_0_U6 ( .A1(b[35]), .A2(DP_reg_b_i_0_n38), .ZN(
        DP_reg_b_i_0_n65) );
  OAI21_X1 DP_reg_b_i_0_U5 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n53), .A(
        DP_reg_b_i_0_n65), .ZN(DP_reg_b_i_0_n40) );
  INV_X1 DP_reg_b_i_0_U4 ( .A(regs_clr_int), .ZN(DP_reg_b_i_0_n41) );
  BUF_X1 DP_reg_b_i_0_U3 ( .A(vIn), .Z(DP_reg_b_i_0_n39) );
  BUF_X1 DP_reg_b_i_0_U2 ( .A(vIn), .Z(DP_reg_b_i_0_n38) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_0_ ( .D(DP_reg_b_i_0_n52), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[11]), .QN(DP_reg_b_i_0_n64) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_1_ ( .D(DP_reg_b_i_0_n51), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[10]), .QN(DP_reg_b_i_0_n63) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_2_ ( .D(DP_reg_b_i_0_n50), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[9]), .QN(DP_reg_b_i_0_n62) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_3_ ( .D(DP_reg_b_i_0_n49), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[8]), .QN(DP_reg_b_i_0_n61) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_4_ ( .D(DP_reg_b_i_0_n48), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[7]), .QN(DP_reg_b_i_0_n60) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_5_ ( .D(DP_reg_b_i_0_n47), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[6]), .QN(DP_reg_b_i_0_n59) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_6_ ( .D(DP_reg_b_i_0_n46), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[5]), .QN(DP_reg_b_i_0_n58) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_7_ ( .D(DP_reg_b_i_0_n45), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[4]), .QN(DP_reg_b_i_0_n57) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_8_ ( .D(DP_reg_b_i_0_n44), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[3]), .QN(DP_reg_b_i_0_n56) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_9_ ( .D(DP_reg_b_i_0_n43), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[2]), .QN(DP_reg_b_i_0_n55) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_10_ ( .D(DP_reg_b_i_0_n42), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[1]), .QN(DP_reg_b_i_0_n54) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_11_ ( .D(DP_reg_b_i_0_n40), .CK(clk), .RN(
        DP_reg_b_i_0_n41), .Q(DP_b_int[0]), .QN(DP_reg_b_i_0_n53) );
  NAND2_X1 DP_reg_b_i_1_U28 ( .A1(b[22]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n66) );
  OAI21_X1 DP_reg_b_i_1_U27 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n54), 
        .A(DP_reg_b_i_1_n66), .ZN(DP_reg_b_i_1_n42) );
  NAND2_X1 DP_reg_b_i_1_U26 ( .A1(b[21]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n67) );
  OAI21_X1 DP_reg_b_i_1_U25 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n55), 
        .A(DP_reg_b_i_1_n67), .ZN(DP_reg_b_i_1_n43) );
  NAND2_X1 DP_reg_b_i_1_U24 ( .A1(b[20]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n68) );
  OAI21_X1 DP_reg_b_i_1_U23 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n56), 
        .A(DP_reg_b_i_1_n68), .ZN(DP_reg_b_i_1_n44) );
  NAND2_X1 DP_reg_b_i_1_U22 ( .A1(b[19]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n69) );
  OAI21_X1 DP_reg_b_i_1_U21 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n57), 
        .A(DP_reg_b_i_1_n69), .ZN(DP_reg_b_i_1_n45) );
  NAND2_X1 DP_reg_b_i_1_U20 ( .A1(b[18]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n70) );
  OAI21_X1 DP_reg_b_i_1_U19 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n58), 
        .A(DP_reg_b_i_1_n70), .ZN(DP_reg_b_i_1_n46) );
  NAND2_X1 DP_reg_b_i_1_U18 ( .A1(b[17]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n71) );
  OAI21_X1 DP_reg_b_i_1_U17 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n59), 
        .A(DP_reg_b_i_1_n71), .ZN(DP_reg_b_i_1_n47) );
  NAND2_X1 DP_reg_b_i_1_U16 ( .A1(b[16]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n72) );
  OAI21_X1 DP_reg_b_i_1_U15 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n60), 
        .A(DP_reg_b_i_1_n72), .ZN(DP_reg_b_i_1_n48) );
  NAND2_X1 DP_reg_b_i_1_U14 ( .A1(b[15]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n73) );
  OAI21_X1 DP_reg_b_i_1_U13 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n61), 
        .A(DP_reg_b_i_1_n73), .ZN(DP_reg_b_i_1_n49) );
  NAND2_X1 DP_reg_b_i_1_U12 ( .A1(b[14]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n74) );
  OAI21_X1 DP_reg_b_i_1_U11 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n62), 
        .A(DP_reg_b_i_1_n74), .ZN(DP_reg_b_i_1_n50) );
  NAND2_X1 DP_reg_b_i_1_U10 ( .A1(b[13]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n75) );
  OAI21_X1 DP_reg_b_i_1_U9 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n63), .A(
        DP_reg_b_i_1_n75), .ZN(DP_reg_b_i_1_n51) );
  NAND2_X1 DP_reg_b_i_1_U8 ( .A1(DP_reg_b_i_1_n39), .A2(b[12]), .ZN(
        DP_reg_b_i_1_n76) );
  OAI21_X1 DP_reg_b_i_1_U7 ( .B1(DP_reg_b_i_1_n39), .B2(DP_reg_b_i_1_n64), .A(
        DP_reg_b_i_1_n76), .ZN(DP_reg_b_i_1_n52) );
  NAND2_X1 DP_reg_b_i_1_U6 ( .A1(b[23]), .A2(DP_reg_b_i_1_n38), .ZN(
        DP_reg_b_i_1_n65) );
  OAI21_X1 DP_reg_b_i_1_U5 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n53), .A(
        DP_reg_b_i_1_n65), .ZN(DP_reg_b_i_1_n40) );
  INV_X1 DP_reg_b_i_1_U4 ( .A(regs_clr_int), .ZN(DP_reg_b_i_1_n41) );
  BUF_X1 DP_reg_b_i_1_U3 ( .A(vIn), .Z(DP_reg_b_i_1_n39) );
  BUF_X1 DP_reg_b_i_1_U2 ( .A(vIn), .Z(DP_reg_b_i_1_n38) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_0_ ( .D(DP_reg_b_i_1_n52), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[23]), .QN(DP_reg_b_i_1_n64) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_1_ ( .D(DP_reg_b_i_1_n51), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[22]), .QN(DP_reg_b_i_1_n63) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_2_ ( .D(DP_reg_b_i_1_n50), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[21]), .QN(DP_reg_b_i_1_n62) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_3_ ( .D(DP_reg_b_i_1_n49), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[20]), .QN(DP_reg_b_i_1_n61) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_4_ ( .D(DP_reg_b_i_1_n48), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[19]), .QN(DP_reg_b_i_1_n60) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_5_ ( .D(DP_reg_b_i_1_n47), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[18]), .QN(DP_reg_b_i_1_n59) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_6_ ( .D(DP_reg_b_i_1_n46), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[17]), .QN(DP_reg_b_i_1_n58) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_7_ ( .D(DP_reg_b_i_1_n45), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[16]), .QN(DP_reg_b_i_1_n57) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_8_ ( .D(DP_reg_b_i_1_n44), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[15]), .QN(DP_reg_b_i_1_n56) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_9_ ( .D(DP_reg_b_i_1_n43), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[14]), .QN(DP_reg_b_i_1_n55) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_10_ ( .D(DP_reg_b_i_1_n42), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[13]), .QN(DP_reg_b_i_1_n54) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_11_ ( .D(DP_reg_b_i_1_n40), .CK(clk), .RN(
        DP_reg_b_i_1_n41), .Q(DP_b_int[12]), .QN(DP_reg_b_i_1_n53) );
  NAND2_X1 DP_reg_b_i_2_U28 ( .A1(b[10]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n66) );
  OAI21_X1 DP_reg_b_i_2_U27 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n54), 
        .A(DP_reg_b_i_2_n66), .ZN(DP_reg_b_i_2_n42) );
  NAND2_X1 DP_reg_b_i_2_U26 ( .A1(b[9]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n67) );
  OAI21_X1 DP_reg_b_i_2_U25 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n55), 
        .A(DP_reg_b_i_2_n67), .ZN(DP_reg_b_i_2_n43) );
  NAND2_X1 DP_reg_b_i_2_U24 ( .A1(b[8]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n68) );
  OAI21_X1 DP_reg_b_i_2_U23 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n56), 
        .A(DP_reg_b_i_2_n68), .ZN(DP_reg_b_i_2_n44) );
  NAND2_X1 DP_reg_b_i_2_U22 ( .A1(b[7]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n69) );
  OAI21_X1 DP_reg_b_i_2_U21 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n57), 
        .A(DP_reg_b_i_2_n69), .ZN(DP_reg_b_i_2_n45) );
  NAND2_X1 DP_reg_b_i_2_U20 ( .A1(b[6]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n70) );
  OAI21_X1 DP_reg_b_i_2_U19 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n58), 
        .A(DP_reg_b_i_2_n70), .ZN(DP_reg_b_i_2_n46) );
  NAND2_X1 DP_reg_b_i_2_U18 ( .A1(b[5]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n71) );
  OAI21_X1 DP_reg_b_i_2_U17 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n59), 
        .A(DP_reg_b_i_2_n71), .ZN(DP_reg_b_i_2_n47) );
  NAND2_X1 DP_reg_b_i_2_U16 ( .A1(b[4]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n72) );
  OAI21_X1 DP_reg_b_i_2_U15 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n60), 
        .A(DP_reg_b_i_2_n72), .ZN(DP_reg_b_i_2_n48) );
  NAND2_X1 DP_reg_b_i_2_U14 ( .A1(b[3]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n73) );
  OAI21_X1 DP_reg_b_i_2_U13 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n61), 
        .A(DP_reg_b_i_2_n73), .ZN(DP_reg_b_i_2_n49) );
  NAND2_X1 DP_reg_b_i_2_U12 ( .A1(b[2]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n74) );
  OAI21_X1 DP_reg_b_i_2_U11 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n62), 
        .A(DP_reg_b_i_2_n74), .ZN(DP_reg_b_i_2_n50) );
  NAND2_X1 DP_reg_b_i_2_U10 ( .A1(b[1]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n75) );
  OAI21_X1 DP_reg_b_i_2_U9 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n63), .A(
        DP_reg_b_i_2_n75), .ZN(DP_reg_b_i_2_n51) );
  NAND2_X1 DP_reg_b_i_2_U8 ( .A1(DP_reg_b_i_2_n39), .A2(b[0]), .ZN(
        DP_reg_b_i_2_n76) );
  OAI21_X1 DP_reg_b_i_2_U7 ( .B1(DP_reg_b_i_2_n39), .B2(DP_reg_b_i_2_n64), .A(
        DP_reg_b_i_2_n76), .ZN(DP_reg_b_i_2_n52) );
  NAND2_X1 DP_reg_b_i_2_U6 ( .A1(b[11]), .A2(DP_reg_b_i_2_n38), .ZN(
        DP_reg_b_i_2_n65) );
  OAI21_X1 DP_reg_b_i_2_U5 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n53), .A(
        DP_reg_b_i_2_n65), .ZN(DP_reg_b_i_2_n40) );
  INV_X1 DP_reg_b_i_2_U4 ( .A(regs_clr_int), .ZN(DP_reg_b_i_2_n41) );
  BUF_X1 DP_reg_b_i_2_U3 ( .A(vIn), .Z(DP_reg_b_i_2_n39) );
  BUF_X1 DP_reg_b_i_2_U2 ( .A(vIn), .Z(DP_reg_b_i_2_n38) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_0_ ( .D(DP_reg_b_i_2_n52), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[35]), .QN(DP_reg_b_i_2_n64) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_1_ ( .D(DP_reg_b_i_2_n51), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[34]), .QN(DP_reg_b_i_2_n63) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_2_ ( .D(DP_reg_b_i_2_n50), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[33]), .QN(DP_reg_b_i_2_n62) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_3_ ( .D(DP_reg_b_i_2_n49), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[32]), .QN(DP_reg_b_i_2_n61) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_4_ ( .D(DP_reg_b_i_2_n48), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[31]), .QN(DP_reg_b_i_2_n60) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_5_ ( .D(DP_reg_b_i_2_n47), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[30]), .QN(DP_reg_b_i_2_n59) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_6_ ( .D(DP_reg_b_i_2_n46), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[29]), .QN(DP_reg_b_i_2_n58) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_7_ ( .D(DP_reg_b_i_2_n45), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[28]), .QN(DP_reg_b_i_2_n57) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_8_ ( .D(DP_reg_b_i_2_n44), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[27]), .QN(DP_reg_b_i_2_n56) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_9_ ( .D(DP_reg_b_i_2_n43), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[26]), .QN(DP_reg_b_i_2_n55) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_10_ ( .D(DP_reg_b_i_2_n42), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[25]), .QN(DP_reg_b_i_2_n54) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_11_ ( .D(DP_reg_b_i_2_n40), .CK(clk), .RN(
        DP_reg_b_i_2_n41), .Q(DP_b_int[24]), .QN(DP_reg_b_i_2_n53) );
  NAND2_X1 DP_reg_sw0_U35 ( .A1(DP_n12), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n13) );
  NAND2_X1 DP_reg_sw0_U34 ( .A1(DP_n11), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n12) );
  NAND2_X1 DP_reg_sw0_U33 ( .A1(DP_n9), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n10) );
  NAND2_X1 DP_reg_sw0_U32 ( .A1(DP_w_8_), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n9) );
  NAND2_X1 DP_reg_sw0_U31 ( .A1(DP_w_5_), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n6) );
  OAI21_X1 DP_reg_sw0_U30 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n19), .A(
        DP_reg_sw0_n6), .ZN(DP_reg_sw0_n32) );
  NAND2_X1 DP_reg_sw0_U29 ( .A1(DP_w_4_), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n5) );
  OAI21_X1 DP_reg_sw0_U28 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n18), .A(
        DP_reg_sw0_n5), .ZN(DP_reg_sw0_n31) );
  NAND2_X1 DP_reg_sw0_U27 ( .A1(DP_w_3_), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n4) );
  OAI21_X1 DP_reg_sw0_U26 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n17), .A(
        DP_reg_sw0_n4), .ZN(DP_reg_sw0_n30) );
  NAND2_X1 DP_reg_sw0_U25 ( .A1(DP_w_2_), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n3) );
  OAI21_X1 DP_reg_sw0_U24 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n16), .A(
        DP_reg_sw0_n3), .ZN(DP_reg_sw0_n29) );
  NAND2_X1 DP_reg_sw0_U23 ( .A1(DP_w_1_), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n2) );
  OAI21_X1 DP_reg_sw0_U22 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n15), .A(
        DP_reg_sw0_n2), .ZN(DP_reg_sw0_n28) );
  NAND2_X1 DP_reg_sw0_U21 ( .A1(DP_reg_sw0_n47), .A2(DP_w_0_), .ZN(
        DP_reg_sw0_n1) );
  OAI21_X1 DP_reg_sw0_U20 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n14), .A(
        DP_reg_sw0_n1), .ZN(DP_reg_sw0_n27) );
  OAI21_X1 DP_reg_sw0_U19 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n26), .A(
        DP_reg_sw0_n13), .ZN(DP_reg_sw0_n40) );
  OAI21_X1 DP_reg_sw0_U18 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n25), .A(
        DP_reg_sw0_n12), .ZN(DP_reg_sw0_n38) );
  NAND2_X1 DP_reg_sw0_U17 ( .A1(DP_n13), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n11) );
  OAI21_X1 DP_reg_sw0_U16 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n24), .A(
        DP_reg_sw0_n11), .ZN(DP_reg_sw0_n37) );
  OAI21_X1 DP_reg_sw0_U15 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n23), .A(
        DP_reg_sw0_n10), .ZN(DP_reg_sw0_n36) );
  OAI21_X1 DP_reg_sw0_U14 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n22), .A(
        DP_reg_sw0_n9), .ZN(DP_reg_sw0_n35) );
  NAND2_X1 DP_reg_sw0_U13 ( .A1(DP_w_7_), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n8) );
  OAI21_X1 DP_reg_sw0_U12 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n21), .A(
        DP_reg_sw0_n8), .ZN(DP_reg_sw0_n34) );
  NAND2_X1 DP_reg_sw0_U11 ( .A1(DP_w_6_), .A2(DP_reg_sw0_n46), .ZN(
        DP_reg_sw0_n7) );
  OAI21_X1 DP_reg_sw0_U10 ( .B1(DP_reg_sw0_n47), .B2(DP_reg_sw0_n20), .A(
        DP_reg_sw0_n7), .ZN(DP_reg_sw0_n33) );
  INV_X1 DP_reg_sw0_U9 ( .A(regs_clr_int), .ZN(DP_reg_sw0_n39) );
  BUF_X1 DP_reg_sw0_U8 ( .A(reg_sw0_en_int), .Z(DP_reg_sw0_n46) );
  BUF_X1 DP_reg_sw0_U7 ( .A(reg_sw0_en_int), .Z(DP_reg_sw0_n47) );
  INV_X2 DP_reg_sw0_U6 ( .A(DP_reg_sw0_n20), .ZN(DP_sw0_6_) );
  INV_X2 DP_reg_sw0_U5 ( .A(DP_reg_sw0_n21), .ZN(DP_sw0_7_) );
  INV_X2 DP_reg_sw0_U4 ( .A(DP_reg_sw0_n19), .ZN(DP_sw0_5_) );
  INV_X2 DP_reg_sw0_U3 ( .A(DP_reg_sw0_n22), .ZN(DP_sw0_8_) );
  INV_X2 DP_reg_sw0_U2 ( .A(DP_reg_sw0_n16), .ZN(DP_sw0_2_) );
  DFFR_X1 DP_reg_sw0_Q_reg_2_ ( .D(DP_reg_sw0_n29), .CK(clk), .RN(
        DP_reg_sw0_n39), .QN(DP_reg_sw0_n16) );
  DFFR_X1 DP_reg_sw0_Q_reg_5_ ( .D(DP_reg_sw0_n32), .CK(clk), .RN(
        DP_reg_sw0_n39), .QN(DP_reg_sw0_n19) );
  DFFR_X1 DP_reg_sw0_Q_reg_0_ ( .D(DP_reg_sw0_n27), .CK(clk), .RN(
        DP_reg_sw0_n39), .Q(DP_sw0_0_), .QN(DP_reg_sw0_n14) );
  DFFR_X1 DP_reg_sw0_Q_reg_1_ ( .D(DP_reg_sw0_n28), .CK(clk), .RN(
        DP_reg_sw0_n39), .Q(DP_sw0_1_), .QN(DP_reg_sw0_n15) );
  DFFR_X1 DP_reg_sw0_Q_reg_3_ ( .D(DP_reg_sw0_n30), .CK(clk), .RN(
        DP_reg_sw0_n39), .Q(DP_sw0_3_), .QN(DP_reg_sw0_n17) );
  DFFR_X1 DP_reg_sw0_Q_reg_4_ ( .D(DP_reg_sw0_n31), .CK(clk), .RN(
        DP_reg_sw0_n39), .Q(DP_sw0_4_), .QN(DP_reg_sw0_n18) );
  DFFR_X1 DP_reg_sw0_Q_reg_6_ ( .D(DP_reg_sw0_n33), .CK(clk), .RN(
        DP_reg_sw0_n39), .QN(DP_reg_sw0_n20) );
  DFFR_X1 DP_reg_sw0_Q_reg_7_ ( .D(DP_reg_sw0_n34), .CK(clk), .RN(
        DP_reg_sw0_n39), .QN(DP_reg_sw0_n21) );
  DFFR_X1 DP_reg_sw0_Q_reg_8_ ( .D(DP_reg_sw0_n35), .CK(clk), .RN(
        DP_reg_sw0_n39), .QN(DP_reg_sw0_n22) );
  DFFR_X1 DP_reg_sw0_Q_reg_9_ ( .D(DP_reg_sw0_n36), .CK(clk), .RN(
        DP_reg_sw0_n39), .Q(DP_sw0_9_), .QN(DP_reg_sw0_n23) );
  DFFR_X1 DP_reg_sw0_Q_reg_10_ ( .D(DP_reg_sw0_n37), .CK(clk), .RN(
        DP_reg_sw0_n39), .Q(DP_sw0_10_), .QN(DP_reg_sw0_n24) );
  DFFR_X1 DP_reg_sw0_Q_reg_11_ ( .D(DP_reg_sw0_n38), .CK(clk), .RN(
        DP_reg_sw0_n39), .Q(DP_sw0_11_), .QN(DP_reg_sw0_n25) );
  DFFR_X1 DP_reg_sw0_Q_reg_12_ ( .D(DP_reg_sw0_n40), .CK(clk), .RN(
        DP_reg_sw0_n39), .Q(DP_sw0_12_), .QN(DP_reg_sw0_n26) );
  NAND2_X1 DP_reg_sw1_U38 ( .A1(DP_reg_sw1_n53), .A2(DP_sw0_0_), .ZN(
        DP_reg_sw1_n92) );
  OAI21_X1 DP_reg_sw1_U37 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n79), .A(
        DP_reg_sw1_n92), .ZN(DP_reg_sw1_n66) );
  OAI21_X1 DP_reg_sw1_U36 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n77), .A(
        DP_reg_sw1_n90), .ZN(DP_reg_sw1_n64) );
  OAI21_X1 DP_reg_sw1_U35 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n48), .A(
        DP_reg_sw1_n91), .ZN(DP_reg_sw1_n65) );
  INV_X2 DP_reg_sw1_U34 ( .A(DP_reg_sw1_n78), .ZN(DP_sw1_1_) );
  OAI21_X1 DP_reg_sw1_U33 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n72), .A(
        DP_reg_sw1_n85), .ZN(DP_reg_sw1_n60) );
  OAI21_X1 DP_reg_sw1_U32 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n46), .A(
        DP_reg_sw1_n84), .ZN(DP_reg_sw1_n59) );
  INV_X2 DP_reg_sw1_U31 ( .A(DP_reg_sw1_n71), .ZN(DP_sw1_8_) );
  INV_X1 DP_reg_sw1_U30 ( .A(DP_reg_sw1_n47), .ZN(DP_reg_sw1_n48) );
  NAND2_X1 DP_reg_sw1_U29 ( .A1(DP_sw0_12_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n80) );
  OAI21_X1 DP_reg_sw1_U28 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n67), .A(
        DP_reg_sw1_n80), .ZN(DP_reg_sw1_n54) );
  NAND2_X1 DP_reg_sw1_U27 ( .A1(DP_sw0_11_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n81) );
  OAI21_X1 DP_reg_sw1_U26 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n68), .A(
        DP_reg_sw1_n81), .ZN(DP_reg_sw1_n56) );
  NAND2_X1 DP_reg_sw1_U25 ( .A1(DP_sw0_10_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n82) );
  OAI21_X1 DP_reg_sw1_U24 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n69), .A(
        DP_reg_sw1_n82), .ZN(DP_reg_sw1_n57) );
  NAND2_X1 DP_reg_sw1_U23 ( .A1(DP_sw0_9_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n83) );
  OAI21_X1 DP_reg_sw1_U22 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n70), .A(
        DP_reg_sw1_n83), .ZN(DP_reg_sw1_n58) );
  NAND2_X1 DP_reg_sw1_U21 ( .A1(DP_sw0_6_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n86) );
  OAI21_X1 DP_reg_sw1_U20 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n73), .A(
        DP_reg_sw1_n86), .ZN(DP_reg_sw1_n61) );
  NAND2_X1 DP_reg_sw1_U19 ( .A1(DP_sw0_4_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n88) );
  OAI21_X1 DP_reg_sw1_U18 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n75), .A(
        DP_reg_sw1_n88), .ZN(DP_reg_sw1_n63) );
  NAND2_X1 DP_reg_sw1_U17 ( .A1(DP_sw0_3_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n89) );
  OAI21_X1 DP_reg_sw1_U16 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n76), .A(
        DP_reg_sw1_n89), .ZN(DP_reg_sw1_n41) );
  NAND2_X1 DP_reg_sw1_U15 ( .A1(DP_sw0_5_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n87) );
  OAI21_X1 DP_reg_sw1_U14 ( .B1(DP_reg_sw1_n53), .B2(DP_reg_sw1_n74), .A(
        DP_reg_sw1_n87), .ZN(DP_reg_sw1_n62) );
  NAND2_X1 DP_reg_sw1_U13 ( .A1(DP_sw0_8_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n84) );
  NAND2_X1 DP_reg_sw1_U12 ( .A1(DP_sw0_7_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n85) );
  NAND2_X1 DP_reg_sw1_U11 ( .A1(DP_sw0_2_), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n90) );
  NAND2_X1 DP_reg_sw1_U10 ( .A1(DP_n1), .A2(DP_reg_sw1_n52), .ZN(
        DP_reg_sw1_n91) );
  INV_X1 DP_reg_sw1_U9 ( .A(regs_clr_int), .ZN(DP_reg_sw1_n55) );
  BUF_X1 DP_reg_sw1_U8 ( .A(reg_sw0_en_int), .Z(DP_reg_sw1_n53) );
  BUF_X1 DP_reg_sw1_U7 ( .A(reg_sw0_en_int), .Z(DP_reg_sw1_n52) );
  INV_X1 DP_reg_sw1_U6 ( .A(DP_reg_sw1_n45), .ZN(DP_reg_sw1_n46) );
  INV_X1 DP_reg_sw1_U5 ( .A(DP_reg_sw1_n72), .ZN(DP_sw1_7_) );
  INV_X2 DP_reg_sw1_U2 ( .A(DP_reg_sw1_n74), .ZN(DP_sw1_5_) );
  DFFR_X1 DP_reg_sw1_Q_reg_5_ ( .D(DP_reg_sw1_n62), .CK(clk), .RN(
        DP_reg_sw1_n55), .QN(DP_reg_sw1_n74) );
  DFFR_X2 DP_reg_sw1_Q_reg_0_ ( .D(DP_reg_sw1_n66), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_sw1_0_), .QN(DP_reg_sw1_n79) );
  DFFR_X1 DP_reg_sw1_Q_reg_3_ ( .D(DP_reg_sw1_n41), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_sw1_3_), .QN(DP_reg_sw1_n76) );
  DFFR_X2 DP_reg_sw1_Q_reg_9_ ( .D(DP_reg_sw1_n58), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_sw1_9_), .QN(DP_reg_sw1_n70) );
  SDFFR_X1 DP_reg_sw1_Q_reg_2_ ( .D(1'b0), .SI(DP_reg_sw1_n64), .SE(1'b1), 
        .CK(clk), .RN(DP_reg_sw1_n55), .Q(DP_sw1_2_), .QN(DP_reg_sw1_n77) );
  DFFR_X1 DP_reg_sw1_Q_reg_1_ ( .D(DP_reg_sw1_n65), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_reg_sw1_n47), .QN(DP_reg_sw1_n78) );
  DFFR_X1 DP_reg_sw1_Q_reg_4_ ( .D(DP_reg_sw1_n63), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_sw1_4_), .QN(DP_reg_sw1_n75) );
  DFFR_X1 DP_reg_sw1_Q_reg_6_ ( .D(DP_reg_sw1_n61), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_sw1_6_), .QN(DP_reg_sw1_n73) );
  DFFR_X1 DP_reg_sw1_Q_reg_7_ ( .D(DP_reg_sw1_n60), .CK(clk), .RN(
        DP_reg_sw1_n55), .QN(DP_reg_sw1_n72) );
  DFFR_X1 DP_reg_sw1_Q_reg_8_ ( .D(DP_reg_sw1_n59), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_reg_sw1_n45), .QN(DP_reg_sw1_n71) );
  DFFR_X1 DP_reg_sw1_Q_reg_10_ ( .D(DP_reg_sw1_n57), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_sw1_10_), .QN(DP_reg_sw1_n69) );
  DFFR_X1 DP_reg_sw1_Q_reg_11_ ( .D(DP_reg_sw1_n56), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_sw1_11_), .QN(DP_reg_sw1_n68) );
  DFFR_X1 DP_reg_sw1_Q_reg_12_ ( .D(DP_reg_sw1_n54), .CK(clk), .RN(
        DP_reg_sw1_n55), .Q(DP_sw1_12_), .QN(DP_reg_sw1_n67) );
  MUX2_X1 DP_reg_out_U15 ( .A(dOut[11]), .B(DP_n15), .S(DP_reg_out_n9), .Z(
        DP_reg_out_n22) );
  MUX2_X1 DP_reg_out_U14 ( .A(dOut[10]), .B(DP_y_out_10_), .S(DP_reg_out_n9), 
        .Z(DP_reg_out_n24) );
  MUX2_X1 DP_reg_out_U13 ( .A(dOut[9]), .B(DP_y_out_9_), .S(DP_reg_out_n9), 
        .Z(DP_reg_out_n35) );
  MUX2_X1 DP_reg_out_U12 ( .A(dOut[8]), .B(DP_y_out_8_), .S(DP_reg_out_n9), 
        .Z(DP_reg_out_n36) );
  MUX2_X1 DP_reg_out_U11 ( .A(dOut[7]), .B(DP_y_out_7_), .S(DP_reg_out_n9), 
        .Z(DP_reg_out_n37) );
  MUX2_X1 DP_reg_out_U10 ( .A(dOut[6]), .B(DP_y_out_6_), .S(DP_reg_out_n9), 
        .Z(DP_reg_out_n38) );
  MUX2_X1 DP_reg_out_U9 ( .A(dOut[5]), .B(DP_y_out_5_), .S(DP_reg_out_n9), .Z(
        DP_reg_out_n39) );
  MUX2_X1 DP_reg_out_U8 ( .A(dOut[4]), .B(DP_y_out_4_), .S(DP_reg_out_n9), .Z(
        DP_reg_out_n40) );
  MUX2_X1 DP_reg_out_U7 ( .A(dOut[3]), .B(DP_y_out_3_), .S(DP_reg_out_n9), .Z(
        DP_reg_out_n41) );
  MUX2_X1 DP_reg_out_U6 ( .A(dOut[2]), .B(DP_y_out_2_), .S(DP_reg_out_n9), .Z(
        DP_reg_out_n42) );
  MUX2_X1 DP_reg_out_U5 ( .A(dOut[1]), .B(DP_y_out_1_), .S(DP_reg_out_n9), .Z(
        DP_reg_out_n43) );
  MUX2_X1 DP_reg_out_U4 ( .A(dOut[0]), .B(DP_y_out_0_), .S(DP_reg_out_n9), .Z(
        DP_reg_out_n44) );
  INV_X1 DP_reg_out_U3 ( .A(regs_clr_int), .ZN(DP_reg_out_n23) );
  BUF_X1 DP_reg_out_U2 ( .A(reg_sw0_en_int), .Z(DP_reg_out_n9) );
  DFFR_X1 DP_reg_out_Q_reg_1_ ( .D(DP_reg_out_n43), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[1]) );
  DFFR_X1 DP_reg_out_Q_reg_8_ ( .D(DP_reg_out_n36), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[8]) );
  DFFR_X1 DP_reg_out_Q_reg_10_ ( .D(DP_reg_out_n24), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[10]) );
  DFFR_X1 DP_reg_out_Q_reg_2_ ( .D(DP_reg_out_n42), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[2]) );
  DFFR_X1 DP_reg_out_Q_reg_3_ ( .D(DP_reg_out_n41), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[3]) );
  DFFR_X1 DP_reg_out_Q_reg_4_ ( .D(DP_reg_out_n40), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[4]) );
  DFFR_X1 DP_reg_out_Q_reg_5_ ( .D(DP_reg_out_n39), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[5]) );
  DFFR_X1 DP_reg_out_Q_reg_6_ ( .D(DP_reg_out_n38), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[6]) );
  DFFR_X1 DP_reg_out_Q_reg_0_ ( .D(DP_reg_out_n44), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[0]) );
  DFFR_X1 DP_reg_out_Q_reg_7_ ( .D(DP_reg_out_n37), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[7]) );
  DFFR_X1 DP_reg_out_Q_reg_9_ ( .D(DP_reg_out_n35), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[9]) );
  DFFR_X1 DP_reg_out_Q_reg_11_ ( .D(DP_reg_out_n22), .CK(clk), .RN(
        DP_reg_out_n23), .Q(dOut[11]) );
  XOR2_X1 DP_add_1_root_add_0_root_add_107_U2 ( .A(DP_sw0_b1_0_), .B(
        DP_sw1_b2_0_), .Z(DP_ff_0_) );
  AND2_X1 DP_add_1_root_add_0_root_add_107_U1 ( .A1(DP_sw1_b2_0_), .A2(
        DP_sw0_b1_0_), .ZN(DP_add_1_root_add_0_root_add_107_carry_1_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_1 ( .A(DP_sw1_b2_1_), .B(
        DP_sw0_b1_1_), .CI(DP_add_1_root_add_0_root_add_107_carry_1_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_2_), .S(DP_ff_1_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_2 ( .A(DP_sw1_b2_2_), .B(
        DP_sw0_b1_2_), .CI(DP_add_1_root_add_0_root_add_107_carry_2_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_3_), .S(DP_ff_2_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_3 ( .A(DP_sw1_b2_3_), .B(
        DP_sw0_b1_3_), .CI(DP_add_1_root_add_0_root_add_107_carry_3_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_4_), .S(DP_ff_3_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_4 ( .A(DP_sw1_b2_4_), .B(
        DP_sw0_b1_4_), .CI(DP_add_1_root_add_0_root_add_107_carry_4_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_5_), .S(DP_ff_4_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_5 ( .A(DP_sw1_b2_5_), .B(
        DP_sw0_b1_5_), .CI(DP_add_1_root_add_0_root_add_107_carry_5_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_6_), .S(DP_ff_5_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_6 ( .A(DP_sw1_b2_6_), .B(
        DP_sw0_b1_6_), .CI(DP_add_1_root_add_0_root_add_107_carry_6_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_7_), .S(DP_ff_6_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_7 ( .A(DP_sw1_b2_7_), .B(
        DP_sw0_b1_7_), .CI(DP_add_1_root_add_0_root_add_107_carry_7_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_8_), .S(DP_ff_7_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_8 ( .A(DP_sw1_b2_8_), .B(
        DP_sw0_b1_8_), .CI(DP_add_1_root_add_0_root_add_107_carry_8_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_9_), .S(DP_ff_8_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_9 ( .A(DP_sw1_b2_9_), .B(
        DP_sw0_b1_9_), .CI(DP_add_1_root_add_0_root_add_107_carry_9_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_10_), .S(DP_ff_9_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_10 ( .A(DP_sw1_b2_10_), .B(
        DP_sw0_b1_10_), .CI(DP_add_1_root_add_0_root_add_107_carry_10_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_11_), .S(DP_ff_10_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_11 ( .A(DP_sw1_b2_11_), .B(
        DP_sw0_b1_11_), .CI(DP_add_1_root_add_0_root_add_107_carry_11_), .CO(
        DP_add_1_root_add_0_root_add_107_carry_12_), .S(DP_ff_11_) );
  FA_X1 DP_add_1_root_add_0_root_add_107_U1_12 ( .A(DP_sw1_b2_11_), .B(
        DP_sw0_b1_11_), .CI(DP_add_1_root_add_0_root_add_107_carry_12_), .S(
        DP_ff_12_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U102 ( .A(DP_w_b0_0_), .B(DP_ff_0_), 
        .Z(DP_y_0_) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U101 ( .A1(
        DP_add_0_root_add_0_root_add_107_n81), .A2(
        DP_add_0_root_add_0_root_add_107_n82), .A3(
        DP_add_0_root_add_0_root_add_107_n80), .ZN(
        DP_add_0_root_add_0_root_add_107_carry_4_) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U100 ( .A1(DP_w_b0_3_), .A2(
        DP_ff_3_), .ZN(DP_add_0_root_add_0_root_add_107_n82) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U99 ( .A1(
        DP_add_0_root_add_0_root_add_107_n26), .A2(DP_ff_3_), .ZN(
        DP_add_0_root_add_0_root_add_107_n81) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U98 ( .A1(DP_w_b0_3_), .A2(
        DP_add_0_root_add_0_root_add_107_carry_3_), .ZN(
        DP_add_0_root_add_0_root_add_107_n80) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U97 ( .A(
        DP_add_0_root_add_0_root_add_107_n34), .B(
        DP_add_0_root_add_0_root_add_107_n79), .Z(DP_y_3_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U96 ( .A(DP_w_b0_3_), .B(DP_ff_3_), 
        .Z(DP_add_0_root_add_0_root_add_107_n79) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U95 ( .A1(DP_w_b0_10_), .A2(
        DP_ff_10_), .ZN(DP_add_0_root_add_0_root_add_107_n78) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U94 ( .A1(
        DP_add_0_root_add_0_root_add_107_n16), .A2(DP_ff_10_), .ZN(
        DP_add_0_root_add_0_root_add_107_n77) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U93 ( .A1(
        DP_add_0_root_add_0_root_add_107_n15), .A2(DP_w_b0_10_), .ZN(
        DP_add_0_root_add_0_root_add_107_n76) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U92 ( .A(
        DP_add_0_root_add_0_root_add_107_n11), .B(
        DP_add_0_root_add_0_root_add_107_n75), .Z(DP_y_10_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U91 ( .A(DP_w_b0_10_), .B(DP_ff_10_), .Z(DP_add_0_root_add_0_root_add_107_n75) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U90 ( .A1(DP_w_b0_7_), .A2(
        DP_ff_7_), .ZN(DP_add_0_root_add_0_root_add_107_n74) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U89 ( .A1(
        DP_add_0_root_add_0_root_add_107_n42), .A2(DP_ff_7_), .ZN(
        DP_add_0_root_add_0_root_add_107_n73) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U88 ( .A1(
        DP_add_0_root_add_0_root_add_107_n62), .A2(DP_w_b0_7_), .ZN(
        DP_add_0_root_add_0_root_add_107_n72) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U87 ( .A(
        DP_add_0_root_add_0_root_add_107_n43), .B(
        DP_add_0_root_add_0_root_add_107_n71), .Z(DP_y_7_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U86 ( .A(DP_w_b0_7_), .B(DP_ff_7_), 
        .Z(DP_add_0_root_add_0_root_add_107_n71) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U85 ( .A1(DP_w_b0_6_), .A2(
        DP_ff_6_), .ZN(DP_add_0_root_add_0_root_add_107_n70) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U84 ( .A1(
        DP_add_0_root_add_0_root_add_107_n54), .A2(DP_ff_6_), .ZN(
        DP_add_0_root_add_0_root_add_107_n69) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U83 ( .A1(
        DP_add_0_root_add_0_root_add_107_carry_6_), .A2(DP_w_b0_6_), .ZN(
        DP_add_0_root_add_0_root_add_107_n68) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U82 ( .A(
        DP_add_0_root_add_0_root_add_107_n60), .B(
        DP_add_0_root_add_0_root_add_107_n67), .Z(DP_y_6_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U81 ( .A(DP_w_b0_6_), .B(DP_ff_6_), 
        .Z(DP_add_0_root_add_0_root_add_107_n67) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U80 ( .A1(DP_w_b0_4_), .A2(
        DP_ff_4_), .ZN(DP_add_0_root_add_0_root_add_107_n66) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U79 ( .A1(
        DP_add_0_root_add_0_root_add_107_n55), .A2(DP_ff_4_), .ZN(
        DP_add_0_root_add_0_root_add_107_n65) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U78 ( .A1(
        DP_add_0_root_add_0_root_add_107_carry_4_), .A2(DP_w_b0_4_), .ZN(
        DP_add_0_root_add_0_root_add_107_n64) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U77 ( .A(
        DP_add_0_root_add_0_root_add_107_n61), .B(
        DP_add_0_root_add_0_root_add_107_n63), .Z(DP_y_4_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U76 ( .A(DP_w_b0_4_), .B(DP_ff_4_), 
        .Z(DP_add_0_root_add_0_root_add_107_n63) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U75 ( .A1(
        DP_add_0_root_add_0_root_add_107_n69), .A2(
        DP_add_0_root_add_0_root_add_107_n68), .A3(
        DP_add_0_root_add_0_root_add_107_n70), .ZN(
        DP_add_0_root_add_0_root_add_107_n62) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U74 ( .A(
        DP_add_0_root_add_0_root_add_107_n55), .Z(
        DP_add_0_root_add_0_root_add_107_n61) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U73 ( .A(
        DP_add_0_root_add_0_root_add_107_n54), .Z(
        DP_add_0_root_add_0_root_add_107_n60) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U72 ( .A1(
        DP_add_0_root_add_0_root_add_107_n57), .A2(
        DP_add_0_root_add_0_root_add_107_n58), .A3(
        DP_add_0_root_add_0_root_add_107_n59), .ZN(
        DP_add_0_root_add_0_root_add_107_carry_6_) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U71 ( .A1(DP_w_b0_5_), .A2(
        DP_ff_5_), .ZN(DP_add_0_root_add_0_root_add_107_n59) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U70 ( .A1(
        DP_add_0_root_add_0_root_add_107_n35), .A2(DP_ff_5_), .ZN(
        DP_add_0_root_add_0_root_add_107_n58) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U69 ( .A1(
        DP_add_0_root_add_0_root_add_107_n24), .A2(DP_w_b0_5_), .ZN(
        DP_add_0_root_add_0_root_add_107_n57) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U68 ( .A(
        DP_add_0_root_add_0_root_add_107_n56), .B(
        DP_add_0_root_add_0_root_add_107_n10), .Z(DP_y_5_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U67 ( .A(DP_w_b0_5_), .B(DP_ff_5_), 
        .Z(DP_add_0_root_add_0_root_add_107_n56) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U66 ( .A1(
        DP_add_0_root_add_0_root_add_107_n81), .A2(
        DP_add_0_root_add_0_root_add_107_n82), .A3(
        DP_add_0_root_add_0_root_add_107_n80), .ZN(
        DP_add_0_root_add_0_root_add_107_n55) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U65 ( .A1(
        DP_add_0_root_add_0_root_add_107_n58), .A2(
        DP_add_0_root_add_0_root_add_107_n57), .A3(
        DP_add_0_root_add_0_root_add_107_n59), .ZN(
        DP_add_0_root_add_0_root_add_107_n54) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U64 ( .A1(
        DP_add_0_root_add_0_root_add_107_n52), .A2(
        DP_add_0_root_add_0_root_add_107_n51), .A3(
        DP_add_0_root_add_0_root_add_107_n53), .ZN(
        DP_add_0_root_add_0_root_add_107_carry_9_) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U63 ( .A1(DP_w_b0_8_), .A2(
        DP_ff_8_), .ZN(DP_add_0_root_add_0_root_add_107_n53) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U62 ( .A1(
        DP_add_0_root_add_0_root_add_107_n14), .A2(DP_ff_8_), .ZN(
        DP_add_0_root_add_0_root_add_107_n52) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U61 ( .A1(
        DP_add_0_root_add_0_root_add_107_n48), .A2(DP_w_b0_8_), .ZN(
        DP_add_0_root_add_0_root_add_107_n51) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U60 ( .A(
        DP_add_0_root_add_0_root_add_107_n49), .B(
        DP_add_0_root_add_0_root_add_107_n50), .Z(DP_y_8_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U59 ( .A(DP_w_b0_8_), .B(DP_ff_8_), 
        .Z(DP_add_0_root_add_0_root_add_107_n50) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U58 ( .A1(
        DP_add_0_root_add_0_root_add_107_n73), .A2(
        DP_add_0_root_add_0_root_add_107_n72), .A3(
        DP_add_0_root_add_0_root_add_107_n74), .ZN(
        DP_add_0_root_add_0_root_add_107_n48) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U57 ( .A1(
        DP_add_0_root_add_0_root_add_107_n25), .A2(
        DP_add_0_root_add_0_root_add_107_n36), .A3(
        DP_add_0_root_add_0_root_add_107_n74), .ZN(
        DP_add_0_root_add_0_root_add_107_n49) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U56 ( .A1(
        DP_add_0_root_add_0_root_add_107_n46), .A2(
        DP_add_0_root_add_0_root_add_107_n45), .A3(
        DP_add_0_root_add_0_root_add_107_n47), .ZN(
        DP_add_0_root_add_0_root_add_107_carry_12_) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U55 ( .A1(DP_w_b0_11_), .A2(
        DP_ff_11_), .ZN(DP_add_0_root_add_0_root_add_107_n47) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U54 ( .A1(
        DP_add_0_root_add_0_root_add_107_n13), .A2(DP_ff_11_), .ZN(
        DP_add_0_root_add_0_root_add_107_n46) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U53 ( .A1(
        DP_add_0_root_add_0_root_add_107_n32), .A2(DP_w_b0_11_), .ZN(
        DP_add_0_root_add_0_root_add_107_n45) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U52 ( .A(
        DP_add_0_root_add_0_root_add_107_n33), .B(
        DP_add_0_root_add_0_root_add_107_n44), .Z(DP_y_11_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U51 ( .A(DP_w_b0_11_), .B(DP_ff_11_), .Z(DP_add_0_root_add_0_root_add_107_n44) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U50 ( .A1(
        DP_add_0_root_add_0_root_add_107_n69), .A2(
        DP_add_0_root_add_0_root_add_107_n68), .A3(
        DP_add_0_root_add_0_root_add_107_n70), .ZN(
        DP_add_0_root_add_0_root_add_107_n42) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U49 ( .A1(
        DP_add_0_root_add_0_root_add_107_n6), .A2(
        DP_add_0_root_add_0_root_add_107_n68), .A3(
        DP_add_0_root_add_0_root_add_107_n70), .ZN(
        DP_add_0_root_add_0_root_add_107_n43) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U48 ( .A(DP_w_b0_1_), .Z(
        DP_add_0_root_add_0_root_add_107_n41) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U47 ( .A1(
        DP_add_0_root_add_0_root_add_107_n38), .A2(
        DP_add_0_root_add_0_root_add_107_n39), .A3(
        DP_add_0_root_add_0_root_add_107_n40), .ZN(
        DP_add_0_root_add_0_root_add_107_carry_2_) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U46 ( .A1(
        DP_add_0_root_add_0_root_add_107_carry_1_), .A2(DP_ff_1_), .ZN(
        DP_add_0_root_add_0_root_add_107_n40) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U45 ( .A1(DP_w_b0_1_), .A2(
        DP_ff_1_), .ZN(DP_add_0_root_add_0_root_add_107_n39) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U44 ( .A1(DP_w_b0_1_), .A2(
        DP_add_0_root_add_0_root_add_107_carry_1_), .ZN(
        DP_add_0_root_add_0_root_add_107_n38) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U43 ( .A(
        DP_add_0_root_add_0_root_add_107_n41), .B(
        DP_add_0_root_add_0_root_add_107_n37), .Z(DP_y_1_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U42 ( .A(
        DP_add_0_root_add_0_root_add_107_carry_1_), .B(DP_ff_1_), .Z(
        DP_add_0_root_add_0_root_add_107_n37) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U41 ( .A(
        DP_add_0_root_add_0_root_add_107_n9), .Z(
        DP_add_0_root_add_0_root_add_107_n36) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U40 ( .A1(
        DP_add_0_root_add_0_root_add_107_n65), .A2(
        DP_add_0_root_add_0_root_add_107_n64), .A3(
        DP_add_0_root_add_0_root_add_107_n66), .ZN(
        DP_add_0_root_add_0_root_add_107_n35) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U39 ( .A(
        DP_add_0_root_add_0_root_add_107_n26), .Z(
        DP_add_0_root_add_0_root_add_107_n34) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U38 ( .A1(
        DP_add_0_root_add_0_root_add_107_n77), .A2(
        DP_add_0_root_add_0_root_add_107_n76), .A3(
        DP_add_0_root_add_0_root_add_107_n78), .ZN(
        DP_add_0_root_add_0_root_add_107_n32) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U37 ( .A1(
        DP_add_0_root_add_0_root_add_107_n77), .A2(
        DP_add_0_root_add_0_root_add_107_n2), .A3(
        DP_add_0_root_add_0_root_add_107_n78), .ZN(
        DP_add_0_root_add_0_root_add_107_n33) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U36 ( .A1(
        DP_add_0_root_add_0_root_add_107_n29), .A2(
        DP_add_0_root_add_0_root_add_107_n31), .A3(
        DP_add_0_root_add_0_root_add_107_n30), .ZN(
        DP_add_0_root_add_0_root_add_107_carry_3_) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U35 ( .A1(DP_w_b0_2_), .A2(
        DP_ff_2_), .ZN(DP_add_0_root_add_0_root_add_107_n31) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U34 ( .A1(
        DP_add_0_root_add_0_root_add_107_carry_2_), .A2(DP_ff_2_), .ZN(
        DP_add_0_root_add_0_root_add_107_n30) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U33 ( .A1(
        DP_add_0_root_add_0_root_add_107_n27), .A2(DP_w_b0_2_), .ZN(
        DP_add_0_root_add_0_root_add_107_n29) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U32 ( .A(
        DP_add_0_root_add_0_root_add_107_n17), .B(
        DP_add_0_root_add_0_root_add_107_n28), .Z(DP_y_2_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U31 ( .A(
        DP_add_0_root_add_0_root_add_107_n8), .B(DP_ff_2_), .Z(
        DP_add_0_root_add_0_root_add_107_n28) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U30 ( .A1(
        DP_add_0_root_add_0_root_add_107_n39), .A2(
        DP_add_0_root_add_0_root_add_107_n38), .A3(
        DP_add_0_root_add_0_root_add_107_n40), .ZN(
        DP_add_0_root_add_0_root_add_107_n27) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U29 ( .A1(
        DP_add_0_root_add_0_root_add_107_n29), .A2(
        DP_add_0_root_add_0_root_add_107_n31), .A3(
        DP_add_0_root_add_0_root_add_107_n30), .ZN(
        DP_add_0_root_add_0_root_add_107_n26) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U28 ( .A(
        DP_add_0_root_add_0_root_add_107_n73), .Z(
        DP_add_0_root_add_0_root_add_107_n25) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U27 ( .A1(
        DP_add_0_root_add_0_root_add_107_n65), .A2(
        DP_add_0_root_add_0_root_add_107_n64), .A3(
        DP_add_0_root_add_0_root_add_107_n66), .ZN(
        DP_add_0_root_add_0_root_add_107_n24) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U26 ( .A1(DP_w_b0_9_), .A2(
        DP_ff_9_), .ZN(DP_add_0_root_add_0_root_add_107_n23) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U25 ( .A1(
        DP_add_0_root_add_0_root_add_107_carry_9_), .A2(DP_ff_9_), .ZN(
        DP_add_0_root_add_0_root_add_107_n22) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U24 ( .A1(
        DP_add_0_root_add_0_root_add_107_n18), .A2(DP_w_b0_9_), .ZN(
        DP_add_0_root_add_0_root_add_107_n21) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U23 ( .A(
        DP_add_0_root_add_0_root_add_107_n12), .B(
        DP_add_0_root_add_0_root_add_107_n20), .Z(DP_y_9_) );
  XOR2_X1 DP_add_0_root_add_0_root_add_107_U22 ( .A(DP_w_b0_9_), .B(DP_ff_9_), 
        .Z(DP_add_0_root_add_0_root_add_107_n20) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_107_U21 ( .A(DP_w_b0_11_), .B(
        DP_ff_12_), .ZN(DP_add_0_root_add_0_root_add_107_n19) );
  XNOR2_X1 DP_add_0_root_add_0_root_add_107_U20 ( .A(
        DP_add_0_root_add_0_root_add_107_carry_12_), .B(
        DP_add_0_root_add_0_root_add_107_n19), .ZN(DP_y_out_11_) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U19 ( .A1(
        DP_add_0_root_add_0_root_add_107_n52), .A2(
        DP_add_0_root_add_0_root_add_107_n51), .A3(
        DP_add_0_root_add_0_root_add_107_n53), .ZN(
        DP_add_0_root_add_0_root_add_107_n18) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U18 ( .A(
        DP_add_0_root_add_0_root_add_107_n27), .Z(
        DP_add_0_root_add_0_root_add_107_n17) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U17 ( .A1(
        DP_add_0_root_add_0_root_add_107_n21), .A2(
        DP_add_0_root_add_0_root_add_107_n22), .A3(
        DP_add_0_root_add_0_root_add_107_n23), .ZN(
        DP_add_0_root_add_0_root_add_107_n15) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U16 ( .A1(
        DP_add_0_root_add_0_root_add_107_n21), .A2(
        DP_add_0_root_add_0_root_add_107_n22), .A3(
        DP_add_0_root_add_0_root_add_107_n23), .ZN(
        DP_add_0_root_add_0_root_add_107_n16) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U15 ( .A1(
        DP_add_0_root_add_0_root_add_107_n9), .A2(
        DP_add_0_root_add_0_root_add_107_n73), .A3(
        DP_add_0_root_add_0_root_add_107_n74), .ZN(
        DP_add_0_root_add_0_root_add_107_n14) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U14 ( .A1(
        DP_add_0_root_add_0_root_add_107_n2), .A2(
        DP_add_0_root_add_0_root_add_107_n77), .A3(
        DP_add_0_root_add_0_root_add_107_n78), .ZN(
        DP_add_0_root_add_0_root_add_107_n13) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U13 ( .A1(
        DP_add_0_root_add_0_root_add_107_n3), .A2(
        DP_add_0_root_add_0_root_add_107_n4), .A3(
        DP_add_0_root_add_0_root_add_107_n53), .ZN(
        DP_add_0_root_add_0_root_add_107_n12) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U12 ( .A1(
        DP_add_0_root_add_0_root_add_107_n21), .A2(
        DP_add_0_root_add_0_root_add_107_n7), .A3(
        DP_add_0_root_add_0_root_add_107_n23), .ZN(
        DP_add_0_root_add_0_root_add_107_n11) );
  NAND3_X1 DP_add_0_root_add_0_root_add_107_U11 ( .A1(
        DP_add_0_root_add_0_root_add_107_n5), .A2(
        DP_add_0_root_add_0_root_add_107_n1), .A3(
        DP_add_0_root_add_0_root_add_107_n66), .ZN(
        DP_add_0_root_add_0_root_add_107_n10) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U10 ( .A1(
        DP_add_0_root_add_0_root_add_107_n62), .A2(DP_w_b0_7_), .ZN(
        DP_add_0_root_add_0_root_add_107_n9) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U9 ( .A(DP_w_b0_2_), .Z(
        DP_add_0_root_add_0_root_add_107_n8) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U8 ( .A(
        DP_add_0_root_add_0_root_add_107_n22), .Z(
        DP_add_0_root_add_0_root_add_107_n7) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U7 ( .A(
        DP_add_0_root_add_0_root_add_107_n69), .Z(
        DP_add_0_root_add_0_root_add_107_n6) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U6 ( .A(
        DP_add_0_root_add_0_root_add_107_n65), .Z(
        DP_add_0_root_add_0_root_add_107_n5) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U5 ( .A(
        DP_add_0_root_add_0_root_add_107_n51), .Z(
        DP_add_0_root_add_0_root_add_107_n4) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U4 ( .A(
        DP_add_0_root_add_0_root_add_107_n52), .Z(
        DP_add_0_root_add_0_root_add_107_n3) );
  NAND2_X1 DP_add_0_root_add_0_root_add_107_U3 ( .A1(
        DP_add_0_root_add_0_root_add_107_n15), .A2(DP_w_b0_10_), .ZN(
        DP_add_0_root_add_0_root_add_107_n2) );
  CLKBUF_X1 DP_add_0_root_add_0_root_add_107_U2 ( .A(
        DP_add_0_root_add_0_root_add_107_n64), .Z(
        DP_add_0_root_add_0_root_add_107_n1) );
  AND2_X2 DP_add_0_root_add_0_root_add_107_U1 ( .A1(DP_ff_0_), .A2(DP_w_b0_0_), 
        .ZN(DP_add_0_root_add_0_root_add_107_carry_1_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U117 ( .A(DP_sw0_a1_0_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_0_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U116 ( .A(DP_sw0_a1_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_10_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U115 ( .A(DP_sw0_a1_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_1_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U114 ( .A(DP_sw0_a1_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_2_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U113 ( .A(DP_sw0_a1_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_3_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U112 ( .A(DP_sw0_a1_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_4_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U111 ( .A(DP_sw0_a1_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_5_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U110 ( .A(DP_sw0_a1_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_6_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U109 ( .A(DP_sw0_a1_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_7_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U108 ( .A(DP_sw0_a1_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_8_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U107 ( .A(DP_sw0_a1_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_9_) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U106 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n6), .B(
        DP_sub_0_root_sub_0_root_sub_104_n1), .ZN(DP_w_0_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U105 ( .A1(DP_fb_10_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n82) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U104 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_10_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n81) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U103 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n19), .A2(DP_fb_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n80) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U102 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n78), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n79), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n77), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_5_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U101 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n35), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n79) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U100 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_4_), .A2(DP_fb_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n78) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U99 ( .A1(DP_fb_4_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n77) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U98 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n76), .B(
        DP_sub_0_root_sub_0_root_sub_104_n34), .Z(DP_w_4_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U97 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n53), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_4_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n76) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U96 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n75), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n74), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n73), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_4_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U95 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n21), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n75) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U94 ( .A1(DP_fb_3_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_carry_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n74) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U93 ( .A1(DP_fb_3_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n73) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U92 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n72), .B(
        DP_sub_0_root_sub_0_root_sub_104_n59), .Z(DP_w_3_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U91 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n14), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_3_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n72) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U90 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n4), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n70), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n69), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_9_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U89 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n12), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n71) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U88 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_8_), .A2(DP_fb_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n70) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U87 ( .A1(DP_fb_8_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n69) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U86 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n68), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n67), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n66), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_8_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U85 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n42), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n68) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U84 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_7_), .A2(DP_fb_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n67) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U83 ( .A1(DP_fb_7_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n66) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U82 ( .A(DP_fb_7_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_7_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n65) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U81 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n37), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n9), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n66), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n64) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U80 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n61), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n62), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n63), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_12_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U79 ( .A1(DP_fb_11_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_12_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n63) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U78 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n60), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_12_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n62) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U77 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n60), .A2(DP_fb_11_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n61) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U76 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n81), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n80), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n82), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n60) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U75 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n21), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n59) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U74 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n57), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n58), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n56), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_2_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U73 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n7), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n58) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U72 ( .A1(DP_fb_1_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n57) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U71 ( .A1(DP_fb_1_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n7), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n56) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U70 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n23), .B(
        DP_sub_0_root_sub_0_root_sub_104_n55), .Z(DP_w_1_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U69 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n8), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_1_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n55) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U68 ( .A(DP_fb_10_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n54) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U67 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n20), .B(
        DP_sub_0_root_sub_0_root_sub_104_n54), .ZN(DP_w_10_) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U66 ( .A(DP_fb_4_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n53) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U65 ( .A(DP_fb_11_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_12_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n52) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U64 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n49), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n50), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n48), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_7_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U63 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_6_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n50) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U62 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n40), .A2(DP_fb_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n49) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U61 ( .A1(DP_fb_6_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n48) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U60 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n47), .B(
        DP_sub_0_root_sub_0_root_sub_104_n41), .Z(DP_w_6_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U59 ( .A(DP_fb_6_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_6_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n47) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U58 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n10), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n45), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n44), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_6_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U57 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_5_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n46) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U56 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n11), .A2(DP_fb_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n45) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U55 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_B_not_5_), .A2(DP_fb_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n44) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U54 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n43), .B(
        DP_sub_0_root_sub_0_root_sub_104_n33), .Z(DP_w_5_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U53 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n5), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_5_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n43) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U52 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n50), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n49), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n48), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n42) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U51 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n45), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n44), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n46), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n40) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U50 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n44), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n36), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n39), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n41) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U49 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n42), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n38) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U48 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n68), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n37) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U47 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n45), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n36) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U46 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n10), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n39) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U45 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n75), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n74), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n73), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n35) );
  AND3_X1 DP_sub_0_root_sub_0_root_sub_104_U44 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n80), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n81), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n82), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n51) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U43 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_carry_4_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n34) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U42 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_carry_12_), .B(
        DP_sub_0_root_sub_0_root_sub_104_n2), .ZN(DP_w_12_) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U41 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n17), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n79), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n77), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n33) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U40 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n30), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n31), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n32), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_10_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U39 ( .A1(DP_fb_9_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n32) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U38 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n28), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n31) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U37 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_9_), .A2(DP_fb_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n30) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U36 ( .A(DP_fb_9_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_9_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n29) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U35 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n70), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n71), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n69), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n28) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U34 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n25), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n26), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n27), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_carry_3_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U33 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_2_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n27) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U32 ( .A1(DP_fb_2_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n26) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U31 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n22), .A2(DP_fb_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n25) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U30 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n13), .B(
        DP_sub_0_root_sub_0_root_sub_104_n24), .Z(DP_w_2_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U29 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n15), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_2_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n24) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U28 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n51), .B(
        DP_sub_0_root_sub_0_root_sub_104_n52), .ZN(DP_w_11_) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U27 ( .A(DP_fb_1_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n23) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U26 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n56), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n57), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n58), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n22) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U25 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n25), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n26), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n27), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n21) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U24 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n30), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n3), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n32), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n19) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U23 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n30), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n3), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n32), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n20) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U22 ( .A(DP_fb_8_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n18) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U21 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n18), .B(
        DP_sub_0_root_sub_0_root_sub_104_n64), .ZN(DP_w_8_) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U20 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n78), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n17) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U19 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n70), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n4), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n69), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n16) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U18 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n22), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n15) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U17 ( .A(DP_fb_3_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n14) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U16 ( .A(DP_fb_2_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n13) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U15 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n68), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n67), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n66), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n12) );
  NAND3_X1 DP_sub_0_root_sub_0_root_sub_104_U14 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n78), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n79), .A3(
        DP_sub_0_root_sub_0_root_sub_104_n77), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n11) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U13 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_carry_5_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n10) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U12 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n67), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n9) );
  OR2_X1 DP_sub_0_root_sub_0_root_sub_104_U11 ( .A1(DP_fb_0_), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_0_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n7) );
  OR2_X1 DP_sub_0_root_sub_0_root_sub_104_U10 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n6), .A2(
        DP_sub_0_root_sub_0_root_sub_104_n1), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n8) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U9 ( .A(DP_fb_0_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n6) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U8 ( .A(DP_fb_5_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n5) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U7 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n12), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n4) );
  XOR2_X2 DP_sub_0_root_sub_0_root_sub_104_U6 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n16), .B(
        DP_sub_0_root_sub_0_root_sub_104_n29), .Z(DP_w_9_) );
  NAND2_X1 DP_sub_0_root_sub_0_root_sub_104_U5 ( .A1(
        DP_sub_0_root_sub_0_root_sub_104_n28), .A2(
        DP_sub_0_root_sub_0_root_sub_104_B_not_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n3) );
  XNOR2_X1 DP_sub_0_root_sub_0_root_sub_104_U4 ( .A(DP_fb_12_), .B(
        DP_sub_0_root_sub_0_root_sub_104_B_not_12_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_n2) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_104_U3 ( .A(DP_sw0_a1_11_), .ZN(
        DP_sub_0_root_sub_0_root_sub_104_B_not_12_) );
  CLKBUF_X1 DP_sub_0_root_sub_0_root_sub_104_U2 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_B_not_0_), .Z(
        DP_sub_0_root_sub_0_root_sub_104_n1) );
  XOR2_X2 DP_sub_0_root_sub_0_root_sub_104_U1 ( .A(
        DP_sub_0_root_sub_0_root_sub_104_n65), .B(
        DP_sub_0_root_sub_0_root_sub_104_n38), .Z(DP_w_7_) );
  XOR2_X1 DP_mult_99_U563 ( .A(DP_b_int[33]), .B(DP_b_int[34]), .Z(
        DP_mult_99_n653) );
  INV_X1 DP_mult_99_U562 ( .A(DP_b_int[34]), .ZN(DP_mult_99_n543) );
  NOR2_X1 DP_mult_99_U561 ( .A1(DP_mult_99_n543), .A2(DP_sw1_1_), .ZN(
        DP_mult_99_n658) );
  INV_X1 DP_mult_99_U560 ( .A(DP_mult_99_n658), .ZN(DP_mult_99_n660) );
  NAND2_X1 DP_mult_99_U559 ( .A1(DP_b_int[34]), .A2(DP_mult_99_n532), .ZN(
        DP_mult_99_n530) );
  XNOR2_X1 DP_mult_99_U558 ( .A(DP_n14), .B(DP_b_int[34]), .ZN(DP_mult_99_n529) );
  OAI22_X1 DP_mult_99_U557 ( .A1(DP_mult_99_n660), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n529), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n659) );
  NAND2_X1 DP_mult_99_U556 ( .A1(DP_mult_99_n653), .A2(DP_mult_99_n659), .ZN(
        DP_mult_99_n656) );
  NAND2_X1 DP_mult_99_U555 ( .A1(DP_mult_99_n658), .A2(DP_mult_99_n659), .ZN(
        DP_mult_99_n657) );
  INV_X1 DP_mult_99_U554 ( .A(DP_n3), .ZN(DP_mult_99_n560) );
  MUX2_X1 DP_mult_99_U553 ( .A(DP_mult_99_n656), .B(DP_mult_99_n657), .S(
        DP_mult_99_n560), .Z(DP_mult_99_n655) );
  INV_X1 DP_mult_99_U552 ( .A(DP_mult_99_n655), .ZN(DP_mult_99_n650) );
  INV_X1 DP_mult_99_U551 ( .A(DP_b_int[32]), .ZN(DP_mult_99_n632) );
  XNOR2_X1 DP_mult_99_U550 ( .A(DP_mult_99_n632), .B(DP_b_int[33]), .ZN(
        DP_mult_99_n654) );
  NAND2_X1 DP_mult_99_U549 ( .A1(DP_mult_99_n546), .A2(DP_mult_99_n654), .ZN(
        DP_mult_99_n545) );
  NAND3_X1 DP_mult_99_U548 ( .A1(DP_mult_99_n653), .A2(DP_mult_99_n560), .A3(
        DP_b_int[32]), .ZN(DP_mult_99_n652) );
  OAI21_X1 DP_mult_99_U547 ( .B1(DP_mult_99_n632), .B2(DP_mult_99_n545), .A(
        DP_mult_99_n652), .ZN(DP_mult_99_n651) );
  AOI222_X1 DP_mult_99_U546 ( .A1(DP_mult_99_n650), .A2(DP_mult_99_n255), .B1(
        DP_mult_99_n651), .B2(DP_mult_99_n650), .C1(DP_mult_99_n651), .C2(
        DP_mult_99_n255), .ZN(DP_mult_99_n649) );
  INV_X1 DP_mult_99_U545 ( .A(DP_mult_99_n649), .ZN(DP_mult_99_n648) );
  AOI222_X1 DP_mult_99_U544 ( .A1(DP_mult_99_n648), .A2(DP_mult_99_n253), .B1(
        DP_mult_99_n648), .B2(DP_mult_99_n254), .C1(DP_mult_99_n254), .C2(
        DP_mult_99_n253), .ZN(DP_mult_99_n647) );
  INV_X1 DP_mult_99_U543 ( .A(DP_mult_99_n647), .ZN(DP_mult_99_n646) );
  AOI222_X1 DP_mult_99_U542 ( .A1(DP_mult_99_n646), .A2(DP_mult_99_n249), .B1(
        DP_mult_99_n646), .B2(DP_mult_99_n252), .C1(DP_mult_99_n252), .C2(
        DP_mult_99_n249), .ZN(DP_mult_99_n645) );
  INV_X1 DP_mult_99_U541 ( .A(DP_mult_99_n645), .ZN(DP_mult_99_n644) );
  AOI222_X1 DP_mult_99_U540 ( .A1(DP_mult_99_n644), .A2(DP_mult_99_n245), .B1(
        DP_mult_99_n644), .B2(DP_mult_99_n248), .C1(DP_mult_99_n248), .C2(
        DP_mult_99_n245), .ZN(DP_mult_99_n643) );
  INV_X1 DP_mult_99_U539 ( .A(DP_mult_99_n643), .ZN(DP_mult_99_n642) );
  AOI222_X1 DP_mult_99_U538 ( .A1(DP_mult_99_n642), .A2(DP_mult_99_n239), .B1(
        DP_mult_99_n642), .B2(DP_mult_99_n244), .C1(DP_mult_99_n244), .C2(
        DP_mult_99_n239), .ZN(DP_mult_99_n639) );
  INV_X1 DP_mult_99_U537 ( .A(DP_mult_99_n233), .ZN(DP_mult_99_n640) );
  INV_X1 DP_mult_99_U536 ( .A(DP_mult_99_n238), .ZN(DP_mult_99_n641) );
  OAI222_X1 DP_mult_99_U535 ( .A1(DP_mult_99_n639), .A2(DP_mult_99_n640), .B1(
        DP_mult_99_n639), .B2(DP_mult_99_n641), .C1(DP_mult_99_n641), .C2(
        DP_mult_99_n640), .ZN(DP_mult_99_n638) );
  AOI222_X1 DP_mult_99_U534 ( .A1(DP_mult_99_n638), .A2(DP_mult_99_n225), .B1(
        DP_mult_99_n638), .B2(DP_mult_99_n232), .C1(DP_mult_99_n232), .C2(
        DP_mult_99_n225), .ZN(DP_mult_99_n635) );
  INV_X1 DP_mult_99_U533 ( .A(DP_mult_99_n217), .ZN(DP_mult_99_n636) );
  INV_X1 DP_mult_99_U532 ( .A(DP_mult_99_n224), .ZN(DP_mult_99_n637) );
  OAI222_X1 DP_mult_99_U531 ( .A1(DP_mult_99_n635), .A2(DP_mult_99_n636), .B1(
        DP_mult_99_n635), .B2(DP_mult_99_n637), .C1(DP_mult_99_n637), .C2(
        DP_mult_99_n636), .ZN(DP_mult_99_n126) );
  XNOR2_X1 DP_mult_99_U530 ( .A(DP_n6), .B(DP_b_int[26]), .ZN(DP_mult_99_n606)
         );
  INV_X1 DP_mult_99_U529 ( .A(DP_b_int[28]), .ZN(DP_mult_99_n622) );
  INV_X1 DP_mult_99_U528 ( .A(DP_b_int[26]), .ZN(DP_mult_99_n624) );
  XNOR2_X1 DP_mult_99_U527 ( .A(DP_mult_99_n624), .B(DP_b_int[27]), .ZN(
        DP_mult_99_n634) );
  NAND2_X1 DP_mult_99_U526 ( .A1(DP_mult_99_n593), .A2(DP_mult_99_n634), .ZN(
        DP_mult_99_n595) );
  XNOR2_X1 DP_mult_99_U525 ( .A(DP_sw1_12_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n608) );
  OAI22_X1 DP_mult_99_U524 ( .A1(DP_mult_99_n606), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n608), .ZN(DP_mult_99_n142) );
  INV_X1 DP_mult_99_U523 ( .A(DP_mult_99_n142), .ZN(DP_mult_99_n143) );
  XNOR2_X1 DP_mult_99_U522 ( .A(DP_n6), .B(DP_b_int[28]), .ZN(DP_mult_99_n590)
         );
  INV_X1 DP_mult_99_U521 ( .A(DP_b_int[30]), .ZN(DP_mult_99_n620) );
  XNOR2_X1 DP_mult_99_U520 ( .A(DP_mult_99_n622), .B(DP_b_int[29]), .ZN(
        DP_mult_99_n633) );
  NAND2_X1 DP_mult_99_U519 ( .A1(DP_mult_99_n577), .A2(DP_mult_99_n633), .ZN(
        DP_mult_99_n579) );
  XNOR2_X1 DP_mult_99_U518 ( .A(DP_sw1_12_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n592) );
  OAI22_X1 DP_mult_99_U517 ( .A1(DP_mult_99_n590), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n592), .ZN(DP_mult_99_n152) );
  INV_X1 DP_mult_99_U516 ( .A(DP_mult_99_n152), .ZN(DP_mult_99_n153) );
  XNOR2_X1 DP_mult_99_U515 ( .A(DP_n6), .B(DP_b_int[30]), .ZN(DP_mult_99_n574)
         );
  XNOR2_X1 DP_mult_99_U514 ( .A(DP_mult_99_n620), .B(DP_b_int[31]), .ZN(
        DP_mult_99_n631) );
  NAND2_X1 DP_mult_99_U513 ( .A1(DP_mult_99_n561), .A2(DP_mult_99_n631), .ZN(
        DP_mult_99_n563) );
  XNOR2_X1 DP_mult_99_U512 ( .A(DP_sw1_12_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n576) );
  OAI22_X1 DP_mult_99_U511 ( .A1(DP_mult_99_n574), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n576), .ZN(DP_mult_99_n166) );
  INV_X1 DP_mult_99_U510 ( .A(DP_mult_99_n166), .ZN(DP_mult_99_n167) );
  XNOR2_X1 DP_mult_99_U509 ( .A(DP_n6), .B(DP_b_int[32]), .ZN(DP_mult_99_n557)
         );
  XNOR2_X1 DP_mult_99_U508 ( .A(DP_sw1_12_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n559) );
  OAI22_X1 DP_mult_99_U507 ( .A1(DP_mult_99_n557), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n559), .ZN(DP_mult_99_n184) );
  INV_X1 DP_mult_99_U506 ( .A(DP_mult_99_n184), .ZN(DP_mult_99_n185) );
  XNOR2_X1 DP_mult_99_U505 ( .A(DP_n5), .B(DP_b_int[26]), .ZN(DP_mult_99_n599)
         );
  XNOR2_X1 DP_mult_99_U504 ( .A(DP_sw1_5_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n600) );
  OAI22_X1 DP_mult_99_U503 ( .A1(DP_mult_99_n599), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n600), .ZN(DP_mult_99_n629) );
  XNOR2_X1 DP_mult_99_U502 ( .A(DP_sw1_8_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n571) );
  XNOR2_X1 DP_mult_99_U501 ( .A(DP_sw1_9_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n572) );
  OAI22_X1 DP_mult_99_U500 ( .A1(DP_mult_99_n571), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n572), .ZN(DP_mult_99_n630) );
  OR2_X1 DP_mult_99_U499 ( .A1(DP_mult_99_n629), .A2(DP_mult_99_n630), .ZN(
        DP_mult_99_n194) );
  XNOR2_X1 DP_mult_99_U498 ( .A(DP_mult_99_n629), .B(DP_mult_99_n630), .ZN(
        DP_mult_99_n195) );
  INV_X1 DP_mult_99_U497 ( .A(DP_b_int[24]), .ZN(DP_mult_99_n626) );
  XNOR2_X1 DP_mult_99_U496 ( .A(DP_mult_99_n626), .B(DP_b_int[25]), .ZN(
        DP_mult_99_n628) );
  NAND2_X1 DP_mult_99_U495 ( .A1(DP_mult_99_n526), .A2(DP_mult_99_n628), .ZN(
        DP_mult_99_n525) );
  OR3_X1 DP_mult_99_U494 ( .A1(DP_mult_99_n526), .A2(DP_n3), .A3(
        DP_mult_99_n626), .ZN(DP_mult_99_n627) );
  OAI21_X1 DP_mult_99_U493 ( .B1(DP_mult_99_n626), .B2(DP_mult_99_n525), .A(
        DP_mult_99_n627), .ZN(DP_mult_99_n256) );
  OR3_X1 DP_mult_99_U492 ( .A1(DP_mult_99_n593), .A2(DP_n3), .A3(
        DP_mult_99_n624), .ZN(DP_mult_99_n625) );
  OAI21_X1 DP_mult_99_U491 ( .B1(DP_mult_99_n624), .B2(DP_mult_99_n595), .A(
        DP_mult_99_n625), .ZN(DP_mult_99_n257) );
  OR3_X1 DP_mult_99_U490 ( .A1(DP_mult_99_n577), .A2(DP_n3), .A3(
        DP_mult_99_n622), .ZN(DP_mult_99_n623) );
  OAI21_X1 DP_mult_99_U489 ( .B1(DP_mult_99_n622), .B2(DP_mult_99_n579), .A(
        DP_mult_99_n623), .ZN(DP_mult_99_n258) );
  OR3_X1 DP_mult_99_U488 ( .A1(DP_mult_99_n561), .A2(DP_n3), .A3(
        DP_mult_99_n620), .ZN(DP_mult_99_n621) );
  OAI21_X1 DP_mult_99_U487 ( .B1(DP_mult_99_n620), .B2(DP_mult_99_n563), .A(
        DP_mult_99_n621), .ZN(DP_mult_99_n259) );
  XNOR2_X1 DP_mult_99_U486 ( .A(DP_n7), .B(DP_b_int[24]), .ZN(DP_mult_99_n619)
         );
  XNOR2_X1 DP_mult_99_U485 ( .A(DP_n6), .B(DP_b_int[24]), .ZN(DP_mult_99_n528)
         );
  OAI22_X1 DP_mult_99_U484 ( .A1(DP_mult_99_n619), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n528), .ZN(DP_mult_99_n263) );
  XNOR2_X1 DP_mult_99_U483 ( .A(DP_sw1_9_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n618) );
  OAI22_X1 DP_mult_99_U482 ( .A1(DP_mult_99_n618), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n619), .ZN(DP_mult_99_n264) );
  XNOR2_X1 DP_mult_99_U481 ( .A(DP_sw1_8_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n617) );
  OAI22_X1 DP_mult_99_U480 ( .A1(DP_mult_99_n617), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n618), .ZN(DP_mult_99_n265) );
  XNOR2_X1 DP_mult_99_U479 ( .A(DP_n8), .B(DP_b_int[24]), .ZN(DP_mult_99_n616)
         );
  OAI22_X1 DP_mult_99_U478 ( .A1(DP_mult_99_n616), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n617), .ZN(DP_mult_99_n266) );
  XNOR2_X1 DP_mult_99_U477 ( .A(DP_n10), .B(DP_b_int[24]), .ZN(DP_mult_99_n615) );
  OAI22_X1 DP_mult_99_U476 ( .A1(DP_mult_99_n615), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n616), .ZN(DP_mult_99_n267) );
  XNOR2_X1 DP_mult_99_U475 ( .A(DP_sw1_5_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n614) );
  OAI22_X1 DP_mult_99_U474 ( .A1(DP_mult_99_n614), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n615), .ZN(DP_mult_99_n268) );
  XNOR2_X1 DP_mult_99_U473 ( .A(DP_n5), .B(DP_b_int[24]), .ZN(DP_mult_99_n613)
         );
  OAI22_X1 DP_mult_99_U472 ( .A1(DP_mult_99_n613), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n614), .ZN(DP_mult_99_n269) );
  XNOR2_X1 DP_mult_99_U471 ( .A(DP_n16), .B(DP_b_int[24]), .ZN(DP_mult_99_n612) );
  OAI22_X1 DP_mult_99_U470 ( .A1(DP_mult_99_n612), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n613), .ZN(DP_mult_99_n270) );
  XNOR2_X1 DP_mult_99_U469 ( .A(DP_n14), .B(DP_b_int[24]), .ZN(DP_mult_99_n611) );
  OAI22_X1 DP_mult_99_U468 ( .A1(DP_mult_99_n611), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n612), .ZN(DP_mult_99_n271) );
  XNOR2_X1 DP_mult_99_U467 ( .A(DP_sw1_1_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n610) );
  OAI22_X1 DP_mult_99_U466 ( .A1(DP_mult_99_n610), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n611), .ZN(DP_mult_99_n272) );
  XNOR2_X1 DP_mult_99_U465 ( .A(DP_n3), .B(DP_b_int[24]), .ZN(DP_mult_99_n609)
         );
  OAI22_X1 DP_mult_99_U464 ( .A1(DP_mult_99_n609), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n610), .ZN(DP_mult_99_n273) );
  NOR2_X1 DP_mult_99_U463 ( .A1(DP_mult_99_n560), .A2(DP_mult_99_n526), .ZN(
        DP_mult_99_n274) );
  AOI21_X1 DP_mult_99_U462 ( .B1(DP_mult_99_n595), .B2(DP_mult_99_n593), .A(
        DP_mult_99_n608), .ZN(DP_mult_99_n607) );
  INV_X1 DP_mult_99_U461 ( .A(DP_mult_99_n607), .ZN(DP_mult_99_n275) );
  XNOR2_X1 DP_mult_99_U460 ( .A(DP_n7), .B(DP_b_int[26]), .ZN(DP_mult_99_n605)
         );
  OAI22_X1 DP_mult_99_U459 ( .A1(DP_mult_99_n605), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n606), .ZN(DP_mult_99_n276) );
  XNOR2_X1 DP_mult_99_U458 ( .A(DP_sw1_9_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n604) );
  OAI22_X1 DP_mult_99_U457 ( .A1(DP_mult_99_n604), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n605), .ZN(DP_mult_99_n277) );
  XNOR2_X1 DP_mult_99_U456 ( .A(DP_sw1_8_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n603) );
  OAI22_X1 DP_mult_99_U455 ( .A1(DP_mult_99_n603), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n604), .ZN(DP_mult_99_n278) );
  XNOR2_X1 DP_mult_99_U454 ( .A(DP_n8), .B(DP_b_int[26]), .ZN(DP_mult_99_n602)
         );
  OAI22_X1 DP_mult_99_U453 ( .A1(DP_mult_99_n602), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n603), .ZN(DP_mult_99_n279) );
  XNOR2_X1 DP_mult_99_U452 ( .A(DP_n10), .B(DP_b_int[26]), .ZN(DP_mult_99_n601) );
  OAI22_X1 DP_mult_99_U451 ( .A1(DP_mult_99_n601), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n602), .ZN(DP_mult_99_n280) );
  OAI22_X1 DP_mult_99_U450 ( .A1(DP_mult_99_n600), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n601), .ZN(DP_mult_99_n281) );
  XNOR2_X1 DP_mult_99_U449 ( .A(DP_n16), .B(DP_b_int[26]), .ZN(DP_mult_99_n598) );
  OAI22_X1 DP_mult_99_U448 ( .A1(DP_mult_99_n598), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n599), .ZN(DP_mult_99_n283) );
  XNOR2_X1 DP_mult_99_U447 ( .A(DP_n14), .B(DP_b_int[26]), .ZN(DP_mult_99_n597) );
  OAI22_X1 DP_mult_99_U446 ( .A1(DP_mult_99_n597), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n598), .ZN(DP_mult_99_n284) );
  XNOR2_X1 DP_mult_99_U445 ( .A(DP_sw1_1_), .B(DP_b_int[26]), .ZN(
        DP_mult_99_n596) );
  OAI22_X1 DP_mult_99_U444 ( .A1(DP_mult_99_n596), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n597), .ZN(DP_mult_99_n285) );
  XNOR2_X1 DP_mult_99_U443 ( .A(DP_n3), .B(DP_b_int[26]), .ZN(DP_mult_99_n594)
         );
  OAI22_X1 DP_mult_99_U442 ( .A1(DP_mult_99_n594), .A2(DP_mult_99_n595), .B1(
        DP_mult_99_n593), .B2(DP_mult_99_n596), .ZN(DP_mult_99_n286) );
  NOR2_X1 DP_mult_99_U441 ( .A1(DP_mult_99_n560), .A2(DP_mult_99_n593), .ZN(
        DP_mult_99_n287) );
  AOI21_X1 DP_mult_99_U440 ( .B1(DP_mult_99_n579), .B2(DP_mult_99_n577), .A(
        DP_mult_99_n592), .ZN(DP_mult_99_n591) );
  INV_X1 DP_mult_99_U439 ( .A(DP_mult_99_n591), .ZN(DP_mult_99_n288) );
  XNOR2_X1 DP_mult_99_U438 ( .A(DP_n7), .B(DP_b_int[28]), .ZN(DP_mult_99_n589)
         );
  OAI22_X1 DP_mult_99_U437 ( .A1(DP_mult_99_n589), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n590), .ZN(DP_mult_99_n289) );
  XNOR2_X1 DP_mult_99_U436 ( .A(DP_sw1_9_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n588) );
  OAI22_X1 DP_mult_99_U435 ( .A1(DP_mult_99_n588), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n589), .ZN(DP_mult_99_n290) );
  XNOR2_X1 DP_mult_99_U434 ( .A(DP_sw1_8_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n587) );
  OAI22_X1 DP_mult_99_U433 ( .A1(DP_mult_99_n587), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n588), .ZN(DP_mult_99_n291) );
  XNOR2_X1 DP_mult_99_U432 ( .A(DP_n8), .B(DP_b_int[28]), .ZN(DP_mult_99_n586)
         );
  OAI22_X1 DP_mult_99_U431 ( .A1(DP_mult_99_n586), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n587), .ZN(DP_mult_99_n292) );
  XNOR2_X1 DP_mult_99_U430 ( .A(DP_n10), .B(DP_b_int[28]), .ZN(DP_mult_99_n585) );
  OAI22_X1 DP_mult_99_U429 ( .A1(DP_mult_99_n585), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n586), .ZN(DP_mult_99_n293) );
  XNOR2_X1 DP_mult_99_U428 ( .A(DP_sw1_5_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n584) );
  OAI22_X1 DP_mult_99_U427 ( .A1(DP_mult_99_n584), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n585), .ZN(DP_mult_99_n294) );
  XNOR2_X1 DP_mult_99_U426 ( .A(DP_n5), .B(DP_b_int[28]), .ZN(DP_mult_99_n583)
         );
  OAI22_X1 DP_mult_99_U425 ( .A1(DP_mult_99_n583), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n584), .ZN(DP_mult_99_n295) );
  XNOR2_X1 DP_mult_99_U424 ( .A(DP_n16), .B(DP_b_int[28]), .ZN(DP_mult_99_n582) );
  OAI22_X1 DP_mult_99_U423 ( .A1(DP_mult_99_n582), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n583), .ZN(DP_mult_99_n296) );
  XNOR2_X1 DP_mult_99_U422 ( .A(DP_n14), .B(DP_b_int[28]), .ZN(DP_mult_99_n581) );
  OAI22_X1 DP_mult_99_U421 ( .A1(DP_mult_99_n581), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n582), .ZN(DP_mult_99_n297) );
  XNOR2_X1 DP_mult_99_U420 ( .A(DP_sw1_1_), .B(DP_b_int[28]), .ZN(
        DP_mult_99_n580) );
  OAI22_X1 DP_mult_99_U419 ( .A1(DP_mult_99_n580), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n581), .ZN(DP_mult_99_n298) );
  XNOR2_X1 DP_mult_99_U418 ( .A(DP_n3), .B(DP_b_int[28]), .ZN(DP_mult_99_n578)
         );
  OAI22_X1 DP_mult_99_U417 ( .A1(DP_mult_99_n578), .A2(DP_mult_99_n579), .B1(
        DP_mult_99_n577), .B2(DP_mult_99_n580), .ZN(DP_mult_99_n299) );
  NOR2_X1 DP_mult_99_U416 ( .A1(DP_mult_99_n560), .A2(DP_mult_99_n577), .ZN(
        DP_mult_99_n300) );
  AOI21_X1 DP_mult_99_U415 ( .B1(DP_mult_99_n563), .B2(DP_mult_99_n561), .A(
        DP_mult_99_n576), .ZN(DP_mult_99_n575) );
  INV_X1 DP_mult_99_U414 ( .A(DP_mult_99_n575), .ZN(DP_mult_99_n301) );
  XNOR2_X1 DP_mult_99_U413 ( .A(DP_n7), .B(DP_b_int[30]), .ZN(DP_mult_99_n573)
         );
  OAI22_X1 DP_mult_99_U412 ( .A1(DP_mult_99_n573), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n574), .ZN(DP_mult_99_n302) );
  OAI22_X1 DP_mult_99_U411 ( .A1(DP_mult_99_n572), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n573), .ZN(DP_mult_99_n303) );
  XNOR2_X1 DP_mult_99_U410 ( .A(DP_n8), .B(DP_b_int[30]), .ZN(DP_mult_99_n570)
         );
  OAI22_X1 DP_mult_99_U409 ( .A1(DP_mult_99_n570), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n571), .ZN(DP_mult_99_n305) );
  XNOR2_X1 DP_mult_99_U408 ( .A(DP_n10), .B(DP_b_int[30]), .ZN(DP_mult_99_n569) );
  OAI22_X1 DP_mult_99_U407 ( .A1(DP_mult_99_n569), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n570), .ZN(DP_mult_99_n306) );
  XNOR2_X1 DP_mult_99_U406 ( .A(DP_sw1_5_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n568) );
  OAI22_X1 DP_mult_99_U405 ( .A1(DP_mult_99_n568), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n569), .ZN(DP_mult_99_n307) );
  XNOR2_X1 DP_mult_99_U404 ( .A(DP_n5), .B(DP_b_int[30]), .ZN(DP_mult_99_n567)
         );
  OAI22_X1 DP_mult_99_U403 ( .A1(DP_mult_99_n567), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n568), .ZN(DP_mult_99_n308) );
  XNOR2_X1 DP_mult_99_U402 ( .A(DP_n16), .B(DP_b_int[30]), .ZN(DP_mult_99_n566) );
  OAI22_X1 DP_mult_99_U401 ( .A1(DP_mult_99_n566), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n567), .ZN(DP_mult_99_n309) );
  XNOR2_X1 DP_mult_99_U400 ( .A(DP_n14), .B(DP_b_int[30]), .ZN(DP_mult_99_n565) );
  OAI22_X1 DP_mult_99_U399 ( .A1(DP_mult_99_n565), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n566), .ZN(DP_mult_99_n310) );
  XNOR2_X1 DP_mult_99_U398 ( .A(DP_sw1_1_), .B(DP_b_int[30]), .ZN(
        DP_mult_99_n564) );
  OAI22_X1 DP_mult_99_U397 ( .A1(DP_mult_99_n564), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n565), .ZN(DP_mult_99_n311) );
  XNOR2_X1 DP_mult_99_U396 ( .A(DP_n3), .B(DP_b_int[30]), .ZN(DP_mult_99_n562)
         );
  OAI22_X1 DP_mult_99_U395 ( .A1(DP_mult_99_n562), .A2(DP_mult_99_n563), .B1(
        DP_mult_99_n561), .B2(DP_mult_99_n564), .ZN(DP_mult_99_n312) );
  NOR2_X1 DP_mult_99_U394 ( .A1(DP_mult_99_n560), .A2(DP_mult_99_n561), .ZN(
        DP_mult_99_n313) );
  AOI21_X1 DP_mult_99_U393 ( .B1(DP_mult_99_n545), .B2(DP_mult_99_n546), .A(
        DP_mult_99_n559), .ZN(DP_mult_99_n558) );
  INV_X1 DP_mult_99_U392 ( .A(DP_mult_99_n558), .ZN(DP_mult_99_n314) );
  XNOR2_X1 DP_mult_99_U391 ( .A(DP_n7), .B(DP_b_int[32]), .ZN(DP_mult_99_n556)
         );
  OAI22_X1 DP_mult_99_U390 ( .A1(DP_mult_99_n556), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n557), .ZN(DP_mult_99_n315) );
  XNOR2_X1 DP_mult_99_U389 ( .A(DP_sw1_9_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n555) );
  OAI22_X1 DP_mult_99_U388 ( .A1(DP_mult_99_n555), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n556), .ZN(DP_mult_99_n316) );
  XNOR2_X1 DP_mult_99_U387 ( .A(DP_sw1_8_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n554) );
  OAI22_X1 DP_mult_99_U386 ( .A1(DP_mult_99_n554), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n555), .ZN(DP_mult_99_n317) );
  XNOR2_X1 DP_mult_99_U385 ( .A(DP_n8), .B(DP_b_int[32]), .ZN(DP_mult_99_n553)
         );
  OAI22_X1 DP_mult_99_U384 ( .A1(DP_mult_99_n553), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n554), .ZN(DP_mult_99_n318) );
  XNOR2_X1 DP_mult_99_U383 ( .A(DP_n10), .B(DP_b_int[32]), .ZN(DP_mult_99_n552) );
  OAI22_X1 DP_mult_99_U382 ( .A1(DP_mult_99_n552), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n553), .ZN(DP_mult_99_n319) );
  XNOR2_X1 DP_mult_99_U381 ( .A(DP_sw1_5_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n551) );
  OAI22_X1 DP_mult_99_U380 ( .A1(DP_mult_99_n551), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n552), .ZN(DP_mult_99_n320) );
  XNOR2_X1 DP_mult_99_U379 ( .A(DP_n5), .B(DP_b_int[32]), .ZN(DP_mult_99_n550)
         );
  OAI22_X1 DP_mult_99_U378 ( .A1(DP_mult_99_n550), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n551), .ZN(DP_mult_99_n321) );
  XNOR2_X1 DP_mult_99_U377 ( .A(DP_n16), .B(DP_b_int[32]), .ZN(DP_mult_99_n549) );
  OAI22_X1 DP_mult_99_U376 ( .A1(DP_mult_99_n549), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n550), .ZN(DP_mult_99_n322) );
  XNOR2_X1 DP_mult_99_U375 ( .A(DP_n14), .B(DP_b_int[32]), .ZN(DP_mult_99_n548) );
  OAI22_X1 DP_mult_99_U374 ( .A1(DP_mult_99_n548), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n549), .ZN(DP_mult_99_n323) );
  XNOR2_X1 DP_mult_99_U373 ( .A(DP_sw1_1_), .B(DP_b_int[32]), .ZN(
        DP_mult_99_n547) );
  OAI22_X1 DP_mult_99_U372 ( .A1(DP_mult_99_n547), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n548), .ZN(DP_mult_99_n324) );
  XNOR2_X1 DP_mult_99_U371 ( .A(DP_n3), .B(DP_b_int[32]), .ZN(DP_mult_99_n544)
         );
  OAI22_X1 DP_mult_99_U370 ( .A1(DP_mult_99_n544), .A2(DP_mult_99_n545), .B1(
        DP_mult_99_n546), .B2(DP_mult_99_n547), .ZN(DP_mult_99_n325) );
  XOR2_X1 DP_mult_99_U369 ( .A(DP_sw1_12_), .B(DP_mult_99_n543), .Z(
        DP_mult_99_n541) );
  AOI21_X1 DP_mult_99_U368 ( .B1(DP_mult_99_n530), .B2(DP_mult_99_n532), .A(
        DP_mult_99_n541), .ZN(DP_mult_99_n542) );
  INV_X1 DP_mult_99_U367 ( .A(DP_mult_99_n542), .ZN(DP_mult_99_n327) );
  XNOR2_X1 DP_mult_99_U366 ( .A(DP_n6), .B(DP_b_int[34]), .ZN(DP_mult_99_n540)
         );
  OAI22_X1 DP_mult_99_U365 ( .A1(DP_mult_99_n540), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n541), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n328) );
  XNOR2_X1 DP_mult_99_U364 ( .A(DP_n7), .B(DP_b_int[34]), .ZN(DP_mult_99_n539)
         );
  OAI22_X1 DP_mult_99_U363 ( .A1(DP_mult_99_n539), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n540), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n329) );
  XNOR2_X1 DP_mult_99_U362 ( .A(DP_sw1_9_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n538) );
  OAI22_X1 DP_mult_99_U361 ( .A1(DP_mult_99_n538), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n539), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n330) );
  XNOR2_X1 DP_mult_99_U360 ( .A(DP_sw1_8_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n537) );
  OAI22_X1 DP_mult_99_U359 ( .A1(DP_mult_99_n537), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n538), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n331) );
  XNOR2_X1 DP_mult_99_U358 ( .A(DP_n8), .B(DP_b_int[34]), .ZN(DP_mult_99_n536)
         );
  OAI22_X1 DP_mult_99_U357 ( .A1(DP_mult_99_n536), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n537), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n332) );
  XNOR2_X1 DP_mult_99_U356 ( .A(DP_n10), .B(DP_b_int[34]), .ZN(DP_mult_99_n535) );
  OAI22_X1 DP_mult_99_U355 ( .A1(DP_mult_99_n535), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n536), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n333) );
  XNOR2_X1 DP_mult_99_U354 ( .A(DP_sw1_5_), .B(DP_b_int[34]), .ZN(
        DP_mult_99_n534) );
  OAI22_X1 DP_mult_99_U353 ( .A1(DP_mult_99_n534), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n535), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n334) );
  XNOR2_X1 DP_mult_99_U352 ( .A(DP_n5), .B(DP_b_int[34]), .ZN(DP_mult_99_n533)
         );
  OAI22_X1 DP_mult_99_U351 ( .A1(DP_mult_99_n533), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n534), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n335) );
  XNOR2_X1 DP_mult_99_U350 ( .A(DP_n16), .B(DP_b_int[34]), .ZN(DP_mult_99_n531) );
  OAI22_X1 DP_mult_99_U349 ( .A1(DP_mult_99_n531), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n533), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n336) );
  OAI22_X1 DP_mult_99_U348 ( .A1(DP_mult_99_n529), .A2(DP_mult_99_n530), .B1(
        DP_mult_99_n531), .B2(DP_mult_99_n532), .ZN(DP_mult_99_n337) );
  XNOR2_X1 DP_mult_99_U347 ( .A(DP_sw1_12_), .B(DP_b_int[24]), .ZN(
        DP_mult_99_n527) );
  OAI22_X1 DP_mult_99_U346 ( .A1(DP_mult_99_n528), .A2(DP_mult_99_n525), .B1(
        DP_mult_99_n526), .B2(DP_mult_99_n527), .ZN(DP_mult_99_n519) );
  AOI21_X1 DP_mult_99_U345 ( .B1(DP_mult_99_n525), .B2(DP_mult_99_n526), .A(
        DP_mult_99_n527), .ZN(DP_mult_99_n522) );
  INV_X1 DP_mult_99_U344 ( .A(DP_mult_99_n522), .ZN(DP_mult_99_n520) );
  INV_X1 DP_mult_99_U343 ( .A(DP_mult_99_n519), .ZN(DP_mult_99_n524) );
  AOI222_X1 DP_mult_99_U342 ( .A1(DP_mult_99_n115), .A2(DP_mult_99_n138), .B1(
        DP_mult_99_n524), .B2(DP_mult_99_n115), .C1(DP_mult_99_n524), .C2(
        DP_mult_99_n138), .ZN(DP_mult_99_n523) );
  OAI22_X1 DP_mult_99_U341 ( .A1(DP_mult_99_n522), .A2(DP_mult_99_n523), .B1(
        DP_mult_99_n524), .B2(DP_mult_99_n523), .ZN(DP_mult_99_n521) );
  AOI21_X1 DP_mult_99_U340 ( .B1(DP_mult_99_n519), .B2(DP_mult_99_n520), .A(
        DP_mult_99_n521), .ZN(DP_sw1_b2_11_) );
  XOR2_X2 DP_mult_99_U339 ( .A(DP_b_int[27]), .B(DP_mult_99_n622), .Z(
        DP_mult_99_n593) );
  XOR2_X2 DP_mult_99_U338 ( .A(DP_b_int[29]), .B(DP_mult_99_n620), .Z(
        DP_mult_99_n577) );
  XOR2_X2 DP_mult_99_U337 ( .A(DP_b_int[31]), .B(DP_mult_99_n632), .Z(
        DP_mult_99_n561) );
  XOR2_X2 DP_mult_99_U336 ( .A(DP_b_int[25]), .B(DP_mult_99_n624), .Z(
        DP_mult_99_n526) );
  INV_X1 DP_mult_99_U335 ( .A(DP_b_int[35]), .ZN(DP_mult_99_n532) );
  INV_X1 DP_mult_99_U334 ( .A(DP_mult_99_n653), .ZN(DP_mult_99_n546) );
  HA_X1 DP_mult_99_U120 ( .A(DP_mult_99_n325), .B(DP_mult_99_n337), .CO(
        DP_mult_99_n254), .S(DP_mult_99_n255) );
  FA_X1 DP_mult_99_U119 ( .A(DP_mult_99_n336), .B(DP_mult_99_n313), .CI(
        DP_mult_99_n324), .CO(DP_mult_99_n252), .S(DP_mult_99_n253) );
  HA_X1 DP_mult_99_U118 ( .A(DP_mult_99_n259), .B(DP_mult_99_n312), .CO(
        DP_mult_99_n250), .S(DP_mult_99_n251) );
  FA_X1 DP_mult_99_U117 ( .A(DP_mult_99_n323), .B(DP_mult_99_n335), .CI(
        DP_mult_99_n251), .CO(DP_mult_99_n248), .S(DP_mult_99_n249) );
  FA_X1 DP_mult_99_U109 ( .A(DP_mult_99_n334), .B(DP_mult_99_n300), .CI(
        DP_mult_99_n322), .CO(DP_mult_99_n246), .S(DP_mult_99_n247) );
  FA_X1 DP_mult_99_U108 ( .A(DP_mult_99_n250), .B(DP_mult_99_n311), .CI(
        DP_mult_99_n247), .CO(DP_mult_99_n244), .S(DP_mult_99_n245) );
  HA_X1 DP_mult_99_U107 ( .A(DP_mult_99_n258), .B(DP_mult_99_n299), .CO(
        DP_mult_99_n242), .S(DP_mult_99_n243) );
  FA_X1 DP_mult_99_U106 ( .A(DP_mult_99_n310), .B(DP_mult_99_n333), .CI(
        DP_mult_99_n321), .CO(DP_mult_99_n240), .S(DP_mult_99_n241) );
  FA_X1 DP_mult_99_U105 ( .A(DP_mult_99_n246), .B(DP_mult_99_n243), .CI(
        DP_mult_99_n241), .CO(DP_mult_99_n238), .S(DP_mult_99_n239) );
  FA_X1 DP_mult_99_U104 ( .A(DP_mult_99_n309), .B(DP_mult_99_n287), .CI(
        DP_mult_99_n332), .CO(DP_mult_99_n236), .S(DP_mult_99_n237) );
  FA_X1 DP_mult_99_U103 ( .A(DP_mult_99_n298), .B(DP_mult_99_n320), .CI(
        DP_mult_99_n242), .CO(DP_mult_99_n234), .S(DP_mult_99_n235) );
  FA_X1 DP_mult_99_U102 ( .A(DP_mult_99_n237), .B(DP_mult_99_n240), .CI(
        DP_mult_99_n235), .CO(DP_mult_99_n232), .S(DP_mult_99_n233) );
  HA_X1 DP_mult_99_U101 ( .A(DP_mult_99_n257), .B(DP_mult_99_n286), .CO(
        DP_mult_99_n230), .S(DP_mult_99_n231) );
  FA_X1 DP_mult_99_U100 ( .A(DP_mult_99_n297), .B(DP_mult_99_n308), .CI(
        DP_mult_99_n319), .CO(DP_mult_99_n228), .S(DP_mult_99_n229) );
  FA_X1 DP_mult_99_U99 ( .A(DP_mult_99_n231), .B(DP_mult_99_n331), .CI(
        DP_mult_99_n236), .CO(DP_mult_99_n226), .S(DP_mult_99_n227) );
  FA_X1 DP_mult_99_U98 ( .A(DP_mult_99_n229), .B(DP_mult_99_n234), .CI(
        DP_mult_99_n227), .CO(DP_mult_99_n224), .S(DP_mult_99_n225) );
  FA_X1 DP_mult_99_U97 ( .A(DP_mult_99_n296), .B(DP_mult_99_n274), .CI(
        DP_mult_99_n330), .CO(DP_mult_99_n222), .S(DP_mult_99_n223) );
  FA_X1 DP_mult_99_U96 ( .A(DP_mult_99_n285), .B(DP_mult_99_n318), .CI(
        DP_mult_99_n307), .CO(DP_mult_99_n220), .S(DP_mult_99_n221) );
  FA_X1 DP_mult_99_U95 ( .A(DP_mult_99_n228), .B(DP_mult_99_n230), .CI(
        DP_mult_99_n223), .CO(DP_mult_99_n218), .S(DP_mult_99_n219) );
  FA_X1 DP_mult_99_U94 ( .A(DP_mult_99_n226), .B(DP_mult_99_n221), .CI(
        DP_mult_99_n219), .CO(DP_mult_99_n216), .S(DP_mult_99_n217) );
  HA_X1 DP_mult_99_U93 ( .A(DP_mult_99_n256), .B(DP_mult_99_n273), .CO(
        DP_mult_99_n214), .S(DP_mult_99_n215) );
  FA_X1 DP_mult_99_U92 ( .A(DP_mult_99_n284), .B(DP_mult_99_n306), .CI(
        DP_mult_99_n329), .CO(DP_mult_99_n212), .S(DP_mult_99_n213) );
  FA_X1 DP_mult_99_U91 ( .A(DP_mult_99_n295), .B(DP_mult_99_n317), .CI(
        DP_mult_99_n215), .CO(DP_mult_99_n210), .S(DP_mult_99_n211) );
  FA_X1 DP_mult_99_U90 ( .A(DP_mult_99_n220), .B(DP_mult_99_n222), .CI(
        DP_mult_99_n213), .CO(DP_mult_99_n208), .S(DP_mult_99_n209) );
  FA_X1 DP_mult_99_U89 ( .A(DP_mult_99_n218), .B(DP_mult_99_n211), .CI(
        DP_mult_99_n209), .CO(DP_mult_99_n206), .S(DP_mult_99_n207) );
  HA_X1 DP_mult_99_U88 ( .A(DP_mult_99_n272), .B(DP_mult_99_n283), .CO(
        DP_mult_99_n204), .S(DP_mult_99_n205) );
  FA_X1 DP_mult_99_U87 ( .A(DP_mult_99_n328), .B(DP_mult_99_n305), .CI(
        DP_mult_99_n294), .CO(DP_mult_99_n202), .S(DP_mult_99_n203) );
  FA_X1 DP_mult_99_U86 ( .A(DP_mult_99_n214), .B(DP_mult_99_n316), .CI(
        DP_mult_99_n205), .CO(DP_mult_99_n200), .S(DP_mult_99_n201) );
  FA_X1 DP_mult_99_U85 ( .A(DP_mult_99_n203), .B(DP_mult_99_n212), .CI(
        DP_mult_99_n210), .CO(DP_mult_99_n198), .S(DP_mult_99_n199) );
  FA_X1 DP_mult_99_U84 ( .A(DP_mult_99_n208), .B(DP_mult_99_n201), .CI(
        DP_mult_99_n199), .CO(DP_mult_99_n196), .S(DP_mult_99_n197) );
  FA_X1 DP_mult_99_U81 ( .A(DP_mult_99_n271), .B(DP_mult_99_n293), .CI(
        DP_mult_99_n327), .CO(DP_mult_99_n192), .S(DP_mult_99_n193) );
  FA_X1 DP_mult_99_U80 ( .A(DP_mult_99_n204), .B(DP_mult_99_n315), .CI(
        DP_mult_99_n195), .CO(DP_mult_99_n190), .S(DP_mult_99_n191) );
  FA_X1 DP_mult_99_U79 ( .A(DP_mult_99_n193), .B(DP_mult_99_n202), .CI(
        DP_mult_99_n200), .CO(DP_mult_99_n188), .S(DP_mult_99_n189) );
  FA_X1 DP_mult_99_U78 ( .A(DP_mult_99_n198), .B(DP_mult_99_n191), .CI(
        DP_mult_99_n189), .CO(DP_mult_99_n186), .S(DP_mult_99_n187) );
  FA_X1 DP_mult_99_U76 ( .A(DP_mult_99_n303), .B(DP_mult_99_n281), .CI(
        DP_mult_99_n185), .CO(DP_mult_99_n182), .S(DP_mult_99_n183) );
  FA_X1 DP_mult_99_U75 ( .A(DP_mult_99_n270), .B(DP_mult_99_n292), .CI(
        DP_mult_99_n194), .CO(DP_mult_99_n180), .S(DP_mult_99_n181) );
  FA_X1 DP_mult_99_U74 ( .A(DP_mult_99_n190), .B(DP_mult_99_n192), .CI(
        DP_mult_99_n183), .CO(DP_mult_99_n178), .S(DP_mult_99_n179) );
  FA_X1 DP_mult_99_U73 ( .A(DP_mult_99_n188), .B(DP_mult_99_n181), .CI(
        DP_mult_99_n179), .CO(DP_mult_99_n176), .S(DP_mult_99_n177) );
  FA_X1 DP_mult_99_U72 ( .A(DP_mult_99_n184), .B(DP_mult_99_n269), .CI(
        DP_mult_99_n314), .CO(DP_mult_99_n174), .S(DP_mult_99_n175) );
  FA_X1 DP_mult_99_U71 ( .A(DP_mult_99_n280), .B(DP_mult_99_n302), .CI(
        DP_mult_99_n291), .CO(DP_mult_99_n172), .S(DP_mult_99_n173) );
  FA_X1 DP_mult_99_U70 ( .A(DP_mult_99_n180), .B(DP_mult_99_n182), .CI(
        DP_mult_99_n173), .CO(DP_mult_99_n170), .S(DP_mult_99_n171) );
  FA_X1 DP_mult_99_U69 ( .A(DP_mult_99_n178), .B(DP_mult_99_n175), .CI(
        DP_mult_99_n171), .CO(DP_mult_99_n168), .S(DP_mult_99_n169) );
  FA_X1 DP_mult_99_U67 ( .A(DP_mult_99_n268), .B(DP_mult_99_n279), .CI(
        DP_mult_99_n167), .CO(DP_mult_99_n164), .S(DP_mult_99_n165) );
  FA_X1 DP_mult_99_U66 ( .A(DP_mult_99_n174), .B(DP_mult_99_n290), .CI(
        DP_mult_99_n172), .CO(DP_mult_99_n162), .S(DP_mult_99_n163) );
  FA_X1 DP_mult_99_U65 ( .A(DP_mult_99_n170), .B(DP_mult_99_n165), .CI(
        DP_mult_99_n163), .CO(DP_mult_99_n160), .S(DP_mult_99_n161) );
  FA_X1 DP_mult_99_U64 ( .A(DP_mult_99_n166), .B(DP_mult_99_n267), .CI(
        DP_mult_99_n301), .CO(DP_mult_99_n158), .S(DP_mult_99_n159) );
  FA_X1 DP_mult_99_U63 ( .A(DP_mult_99_n278), .B(DP_mult_99_n289), .CI(
        DP_mult_99_n164), .CO(DP_mult_99_n156), .S(DP_mult_99_n157) );
  FA_X1 DP_mult_99_U62 ( .A(DP_mult_99_n162), .B(DP_mult_99_n159), .CI(
        DP_mult_99_n157), .CO(DP_mult_99_n154), .S(DP_mult_99_n155) );
  FA_X1 DP_mult_99_U60 ( .A(DP_mult_99_n266), .B(DP_mult_99_n277), .CI(
        DP_mult_99_n153), .CO(DP_mult_99_n150), .S(DP_mult_99_n151) );
  FA_X1 DP_mult_99_U59 ( .A(DP_mult_99_n151), .B(DP_mult_99_n158), .CI(
        DP_mult_99_n156), .CO(DP_mult_99_n148), .S(DP_mult_99_n149) );
  FA_X1 DP_mult_99_U58 ( .A(DP_mult_99_n265), .B(DP_mult_99_n152), .CI(
        DP_mult_99_n288), .CO(DP_mult_99_n146), .S(DP_mult_99_n147) );
  FA_X1 DP_mult_99_U57 ( .A(DP_mult_99_n150), .B(DP_mult_99_n276), .CI(
        DP_mult_99_n147), .CO(DP_mult_99_n144), .S(DP_mult_99_n145) );
  FA_X1 DP_mult_99_U55 ( .A(DP_mult_99_n143), .B(DP_mult_99_n264), .CI(
        DP_mult_99_n146), .CO(DP_mult_99_n140), .S(DP_mult_99_n141) );
  FA_X1 DP_mult_99_U54 ( .A(DP_mult_99_n263), .B(DP_mult_99_n142), .CI(
        DP_mult_99_n275), .CO(DP_mult_99_n138), .S(DP_mult_99_n139) );
  FA_X1 DP_mult_99_U42 ( .A(DP_mult_99_n207), .B(DP_mult_99_n216), .CI(
        DP_mult_99_n126), .CO(DP_mult_99_n125), .S(DP_sw1_b2_0_) );
  FA_X1 DP_mult_99_U41 ( .A(DP_mult_99_n197), .B(DP_mult_99_n206), .CI(
        DP_mult_99_n125), .CO(DP_mult_99_n124), .S(DP_sw1_b2_1_) );
  FA_X1 DP_mult_99_U40 ( .A(DP_mult_99_n187), .B(DP_mult_99_n196), .CI(
        DP_mult_99_n124), .CO(DP_mult_99_n123), .S(DP_sw1_b2_2_) );
  FA_X1 DP_mult_99_U39 ( .A(DP_mult_99_n177), .B(DP_mult_99_n186), .CI(
        DP_mult_99_n123), .CO(DP_mult_99_n122), .S(DP_sw1_b2_3_) );
  FA_X1 DP_mult_99_U38 ( .A(DP_mult_99_n169), .B(DP_mult_99_n176), .CI(
        DP_mult_99_n122), .CO(DP_mult_99_n121), .S(DP_sw1_b2_4_) );
  FA_X1 DP_mult_99_U37 ( .A(DP_mult_99_n161), .B(DP_mult_99_n168), .CI(
        DP_mult_99_n121), .CO(DP_mult_99_n120), .S(DP_sw1_b2_5_) );
  FA_X1 DP_mult_99_U36 ( .A(DP_mult_99_n155), .B(DP_mult_99_n160), .CI(
        DP_mult_99_n120), .CO(DP_mult_99_n119), .S(DP_sw1_b2_6_) );
  FA_X1 DP_mult_99_U30 ( .A(DP_mult_99_n149), .B(DP_mult_99_n154), .CI(
        DP_mult_99_n119), .CO(DP_mult_99_n118), .S(DP_sw1_b2_7_) );
  FA_X1 DP_mult_99_U20 ( .A(DP_mult_99_n145), .B(DP_mult_99_n148), .CI(
        DP_mult_99_n118), .CO(DP_mult_99_n117), .S(DP_sw1_b2_8_) );
  FA_X1 DP_mult_99_U10 ( .A(DP_mult_99_n141), .B(DP_mult_99_n144), .CI(
        DP_mult_99_n117), .CO(DP_mult_99_n116), .S(DP_sw1_b2_9_) );
  FA_X1 DP_mult_99_U9 ( .A(DP_mult_99_n140), .B(DP_mult_99_n139), .CI(
        DP_mult_99_n116), .CO(DP_mult_99_n115), .S(DP_sw1_b2_10_) );
  XOR2_X1 DP_mult_98_U564 ( .A(DP_b_int[21]), .B(DP_b_int[22]), .Z(
        DP_mult_98_n654) );
  INV_X1 DP_mult_98_U563 ( .A(DP_b_int[22]), .ZN(DP_mult_98_n544) );
  NOR2_X1 DP_mult_98_U562 ( .A1(DP_mult_98_n544), .A2(DP_n1), .ZN(
        DP_mult_98_n659) );
  INV_X1 DP_mult_98_U561 ( .A(DP_mult_98_n659), .ZN(DP_mult_98_n661) );
  NAND2_X1 DP_mult_98_U560 ( .A1(DP_b_int[22]), .A2(DP_mult_98_n533), .ZN(
        DP_mult_98_n531) );
  XNOR2_X1 DP_mult_98_U559 ( .A(DP_sw0_2_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n530) );
  OAI22_X1 DP_mult_98_U558 ( .A1(DP_mult_98_n661), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n530), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n660) );
  NAND2_X1 DP_mult_98_U557 ( .A1(DP_mult_98_n654), .A2(DP_mult_98_n660), .ZN(
        DP_mult_98_n657) );
  NAND2_X1 DP_mult_98_U556 ( .A1(DP_mult_98_n659), .A2(DP_mult_98_n660), .ZN(
        DP_mult_98_n658) );
  INV_X1 DP_mult_98_U555 ( .A(DP_mult_98_n519), .ZN(DP_mult_98_n561) );
  MUX2_X1 DP_mult_98_U554 ( .A(DP_mult_98_n657), .B(DP_mult_98_n658), .S(
        DP_mult_98_n561), .Z(DP_mult_98_n656) );
  INV_X1 DP_mult_98_U553 ( .A(DP_mult_98_n656), .ZN(DP_mult_98_n651) );
  INV_X1 DP_mult_98_U552 ( .A(DP_b_int[20]), .ZN(DP_mult_98_n633) );
  XNOR2_X1 DP_mult_98_U551 ( .A(DP_mult_98_n633), .B(DP_b_int[21]), .ZN(
        DP_mult_98_n655) );
  NAND2_X1 DP_mult_98_U550 ( .A1(DP_mult_98_n547), .A2(DP_mult_98_n655), .ZN(
        DP_mult_98_n546) );
  NAND3_X1 DP_mult_98_U549 ( .A1(DP_mult_98_n654), .A2(DP_mult_98_n561), .A3(
        DP_b_int[20]), .ZN(DP_mult_98_n653) );
  OAI21_X1 DP_mult_98_U548 ( .B1(DP_mult_98_n633), .B2(DP_mult_98_n546), .A(
        DP_mult_98_n653), .ZN(DP_mult_98_n652) );
  AOI222_X1 DP_mult_98_U547 ( .A1(DP_mult_98_n651), .A2(DP_mult_98_n255), .B1(
        DP_mult_98_n652), .B2(DP_mult_98_n651), .C1(DP_mult_98_n652), .C2(
        DP_mult_98_n255), .ZN(DP_mult_98_n650) );
  INV_X1 DP_mult_98_U546 ( .A(DP_mult_98_n650), .ZN(DP_mult_98_n649) );
  AOI222_X1 DP_mult_98_U545 ( .A1(DP_mult_98_n649), .A2(DP_mult_98_n253), .B1(
        DP_mult_98_n649), .B2(DP_mult_98_n254), .C1(DP_mult_98_n254), .C2(
        DP_mult_98_n253), .ZN(DP_mult_98_n648) );
  INV_X1 DP_mult_98_U544 ( .A(DP_mult_98_n648), .ZN(DP_mult_98_n647) );
  AOI222_X1 DP_mult_98_U543 ( .A1(DP_mult_98_n647), .A2(DP_mult_98_n249), .B1(
        DP_mult_98_n647), .B2(DP_mult_98_n252), .C1(DP_mult_98_n252), .C2(
        DP_mult_98_n249), .ZN(DP_mult_98_n646) );
  INV_X1 DP_mult_98_U542 ( .A(DP_mult_98_n646), .ZN(DP_mult_98_n645) );
  AOI222_X1 DP_mult_98_U541 ( .A1(DP_mult_98_n645), .A2(DP_mult_98_n245), .B1(
        DP_mult_98_n645), .B2(DP_mult_98_n248), .C1(DP_mult_98_n248), .C2(
        DP_mult_98_n245), .ZN(DP_mult_98_n644) );
  INV_X1 DP_mult_98_U540 ( .A(DP_mult_98_n644), .ZN(DP_mult_98_n643) );
  AOI222_X1 DP_mult_98_U539 ( .A1(DP_mult_98_n643), .A2(DP_mult_98_n239), .B1(
        DP_mult_98_n643), .B2(DP_mult_98_n244), .C1(DP_mult_98_n244), .C2(
        DP_mult_98_n239), .ZN(DP_mult_98_n640) );
  INV_X1 DP_mult_98_U538 ( .A(DP_mult_98_n233), .ZN(DP_mult_98_n641) );
  INV_X1 DP_mult_98_U537 ( .A(DP_mult_98_n238), .ZN(DP_mult_98_n642) );
  OAI222_X1 DP_mult_98_U536 ( .A1(DP_mult_98_n640), .A2(DP_mult_98_n641), .B1(
        DP_mult_98_n640), .B2(DP_mult_98_n642), .C1(DP_mult_98_n642), .C2(
        DP_mult_98_n641), .ZN(DP_mult_98_n639) );
  AOI222_X1 DP_mult_98_U535 ( .A1(DP_mult_98_n639), .A2(DP_mult_98_n225), .B1(
        DP_mult_98_n639), .B2(DP_mult_98_n232), .C1(DP_mult_98_n232), .C2(
        DP_mult_98_n225), .ZN(DP_mult_98_n636) );
  INV_X1 DP_mult_98_U534 ( .A(DP_mult_98_n217), .ZN(DP_mult_98_n637) );
  INV_X1 DP_mult_98_U533 ( .A(DP_mult_98_n224), .ZN(DP_mult_98_n638) );
  OAI222_X1 DP_mult_98_U532 ( .A1(DP_mult_98_n636), .A2(DP_mult_98_n637), .B1(
        DP_mult_98_n636), .B2(DP_mult_98_n638), .C1(DP_mult_98_n638), .C2(
        DP_mult_98_n637), .ZN(DP_mult_98_n126) );
  XNOR2_X1 DP_mult_98_U531 ( .A(DP_sw0_11_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n607) );
  INV_X1 DP_mult_98_U530 ( .A(DP_b_int[16]), .ZN(DP_mult_98_n623) );
  INV_X1 DP_mult_98_U529 ( .A(DP_b_int[14]), .ZN(DP_mult_98_n625) );
  XNOR2_X1 DP_mult_98_U528 ( .A(DP_mult_98_n625), .B(DP_b_int[15]), .ZN(
        DP_mult_98_n635) );
  NAND2_X1 DP_mult_98_U527 ( .A1(DP_mult_98_n594), .A2(DP_mult_98_n635), .ZN(
        DP_mult_98_n596) );
  XNOR2_X1 DP_mult_98_U526 ( .A(DP_sw0_12_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n609) );
  OAI22_X1 DP_mult_98_U525 ( .A1(DP_mult_98_n607), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n609), .ZN(DP_mult_98_n142) );
  INV_X1 DP_mult_98_U524 ( .A(DP_mult_98_n142), .ZN(DP_mult_98_n143) );
  XNOR2_X1 DP_mult_98_U523 ( .A(DP_sw0_11_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n591) );
  INV_X1 DP_mult_98_U522 ( .A(DP_b_int[18]), .ZN(DP_mult_98_n621) );
  XNOR2_X1 DP_mult_98_U521 ( .A(DP_mult_98_n623), .B(DP_b_int[17]), .ZN(
        DP_mult_98_n634) );
  NAND2_X1 DP_mult_98_U520 ( .A1(DP_mult_98_n578), .A2(DP_mult_98_n634), .ZN(
        DP_mult_98_n580) );
  XNOR2_X1 DP_mult_98_U519 ( .A(DP_sw0_12_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n593) );
  OAI22_X1 DP_mult_98_U518 ( .A1(DP_mult_98_n591), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n593), .ZN(DP_mult_98_n152) );
  INV_X1 DP_mult_98_U517 ( .A(DP_mult_98_n152), .ZN(DP_mult_98_n153) );
  XNOR2_X1 DP_mult_98_U516 ( .A(DP_sw0_11_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n575) );
  XNOR2_X1 DP_mult_98_U515 ( .A(DP_mult_98_n621), .B(DP_b_int[19]), .ZN(
        DP_mult_98_n632) );
  NAND2_X1 DP_mult_98_U514 ( .A1(DP_mult_98_n562), .A2(DP_mult_98_n632), .ZN(
        DP_mult_98_n564) );
  XNOR2_X1 DP_mult_98_U513 ( .A(DP_sw0_12_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n577) );
  OAI22_X1 DP_mult_98_U512 ( .A1(DP_mult_98_n575), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n577), .ZN(DP_mult_98_n166) );
  INV_X1 DP_mult_98_U511 ( .A(DP_mult_98_n166), .ZN(DP_mult_98_n167) );
  XNOR2_X1 DP_mult_98_U510 ( .A(DP_sw0_11_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n558) );
  XNOR2_X1 DP_mult_98_U509 ( .A(DP_sw0_12_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n560) );
  OAI22_X1 DP_mult_98_U508 ( .A1(DP_mult_98_n558), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n560), .ZN(DP_mult_98_n184) );
  INV_X1 DP_mult_98_U507 ( .A(DP_mult_98_n184), .ZN(DP_mult_98_n185) );
  XNOR2_X1 DP_mult_98_U506 ( .A(DP_sw0_4_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n600) );
  XNOR2_X1 DP_mult_98_U505 ( .A(DP_sw0_5_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n601) );
  OAI22_X1 DP_mult_98_U504 ( .A1(DP_mult_98_n600), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n601), .ZN(DP_mult_98_n630) );
  XNOR2_X1 DP_mult_98_U503 ( .A(DP_sw0_8_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n572) );
  XNOR2_X1 DP_mult_98_U502 ( .A(DP_sw0_9_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n573) );
  OAI22_X1 DP_mult_98_U501 ( .A1(DP_mult_98_n572), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n573), .ZN(DP_mult_98_n631) );
  OR2_X1 DP_mult_98_U500 ( .A1(DP_mult_98_n630), .A2(DP_mult_98_n631), .ZN(
        DP_mult_98_n194) );
  XNOR2_X1 DP_mult_98_U499 ( .A(DP_mult_98_n630), .B(DP_mult_98_n631), .ZN(
        DP_mult_98_n195) );
  INV_X1 DP_mult_98_U498 ( .A(DP_b_int[12]), .ZN(DP_mult_98_n627) );
  XNOR2_X1 DP_mult_98_U497 ( .A(DP_mult_98_n627), .B(DP_b_int[13]), .ZN(
        DP_mult_98_n629) );
  NAND2_X1 DP_mult_98_U496 ( .A1(DP_mult_98_n527), .A2(DP_mult_98_n629), .ZN(
        DP_mult_98_n526) );
  OR3_X1 DP_mult_98_U495 ( .A1(DP_mult_98_n527), .A2(DP_mult_98_n519), .A3(
        DP_mult_98_n627), .ZN(DP_mult_98_n628) );
  OAI21_X1 DP_mult_98_U494 ( .B1(DP_mult_98_n627), .B2(DP_mult_98_n526), .A(
        DP_mult_98_n628), .ZN(DP_mult_98_n256) );
  OR3_X1 DP_mult_98_U493 ( .A1(DP_mult_98_n594), .A2(DP_mult_98_n519), .A3(
        DP_mult_98_n625), .ZN(DP_mult_98_n626) );
  OAI21_X1 DP_mult_98_U492 ( .B1(DP_mult_98_n625), .B2(DP_mult_98_n596), .A(
        DP_mult_98_n626), .ZN(DP_mult_98_n257) );
  OR3_X1 DP_mult_98_U491 ( .A1(DP_mult_98_n578), .A2(DP_mult_98_n519), .A3(
        DP_mult_98_n623), .ZN(DP_mult_98_n624) );
  OAI21_X1 DP_mult_98_U490 ( .B1(DP_mult_98_n623), .B2(DP_mult_98_n580), .A(
        DP_mult_98_n624), .ZN(DP_mult_98_n258) );
  OR3_X1 DP_mult_98_U489 ( .A1(DP_mult_98_n562), .A2(DP_mult_98_n519), .A3(
        DP_mult_98_n621), .ZN(DP_mult_98_n622) );
  OAI21_X1 DP_mult_98_U488 ( .B1(DP_mult_98_n621), .B2(DP_mult_98_n564), .A(
        DP_mult_98_n622), .ZN(DP_mult_98_n259) );
  XNOR2_X1 DP_mult_98_U487 ( .A(DP_sw0_10_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n620) );
  XNOR2_X1 DP_mult_98_U486 ( .A(DP_sw0_11_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n529) );
  OAI22_X1 DP_mult_98_U485 ( .A1(DP_mult_98_n620), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n529), .ZN(DP_mult_98_n263) );
  XNOR2_X1 DP_mult_98_U484 ( .A(DP_sw0_9_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n619) );
  OAI22_X1 DP_mult_98_U483 ( .A1(DP_mult_98_n619), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n620), .ZN(DP_mult_98_n264) );
  XNOR2_X1 DP_mult_98_U482 ( .A(DP_sw0_8_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n618) );
  OAI22_X1 DP_mult_98_U481 ( .A1(DP_mult_98_n618), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n619), .ZN(DP_mult_98_n265) );
  XNOR2_X1 DP_mult_98_U480 ( .A(DP_sw0_7_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n617) );
  OAI22_X1 DP_mult_98_U479 ( .A1(DP_mult_98_n617), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n618), .ZN(DP_mult_98_n266) );
  XNOR2_X1 DP_mult_98_U478 ( .A(DP_sw0_6_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n616) );
  OAI22_X1 DP_mult_98_U477 ( .A1(DP_mult_98_n616), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n617), .ZN(DP_mult_98_n267) );
  XNOR2_X1 DP_mult_98_U476 ( .A(DP_sw0_5_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n615) );
  OAI22_X1 DP_mult_98_U475 ( .A1(DP_mult_98_n615), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n616), .ZN(DP_mult_98_n268) );
  XNOR2_X1 DP_mult_98_U474 ( .A(DP_sw0_4_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n614) );
  OAI22_X1 DP_mult_98_U473 ( .A1(DP_mult_98_n614), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n615), .ZN(DP_mult_98_n269) );
  XNOR2_X1 DP_mult_98_U472 ( .A(DP_sw0_3_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n613) );
  OAI22_X1 DP_mult_98_U471 ( .A1(DP_mult_98_n613), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n614), .ZN(DP_mult_98_n270) );
  XNOR2_X1 DP_mult_98_U470 ( .A(DP_sw0_2_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n612) );
  OAI22_X1 DP_mult_98_U469 ( .A1(DP_mult_98_n612), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n613), .ZN(DP_mult_98_n271) );
  XNOR2_X1 DP_mult_98_U468 ( .A(DP_n1), .B(DP_b_int[12]), .ZN(DP_mult_98_n611)
         );
  OAI22_X1 DP_mult_98_U467 ( .A1(DP_mult_98_n611), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n612), .ZN(DP_mult_98_n272) );
  XNOR2_X1 DP_mult_98_U466 ( .A(DP_mult_98_n519), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n610) );
  OAI22_X1 DP_mult_98_U465 ( .A1(DP_mult_98_n610), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n611), .ZN(DP_mult_98_n273) );
  NOR2_X1 DP_mult_98_U464 ( .A1(DP_mult_98_n561), .A2(DP_mult_98_n527), .ZN(
        DP_mult_98_n274) );
  AOI21_X1 DP_mult_98_U463 ( .B1(DP_mult_98_n596), .B2(DP_mult_98_n594), .A(
        DP_mult_98_n609), .ZN(DP_mult_98_n608) );
  INV_X1 DP_mult_98_U462 ( .A(DP_mult_98_n608), .ZN(DP_mult_98_n275) );
  XNOR2_X1 DP_mult_98_U461 ( .A(DP_sw0_10_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n606) );
  OAI22_X1 DP_mult_98_U460 ( .A1(DP_mult_98_n606), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n607), .ZN(DP_mult_98_n276) );
  XNOR2_X1 DP_mult_98_U459 ( .A(DP_sw0_9_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n605) );
  OAI22_X1 DP_mult_98_U458 ( .A1(DP_mult_98_n605), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n606), .ZN(DP_mult_98_n277) );
  XNOR2_X1 DP_mult_98_U457 ( .A(DP_sw0_8_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n604) );
  OAI22_X1 DP_mult_98_U456 ( .A1(DP_mult_98_n604), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n605), .ZN(DP_mult_98_n278) );
  XNOR2_X1 DP_mult_98_U455 ( .A(DP_sw0_7_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n603) );
  OAI22_X1 DP_mult_98_U454 ( .A1(DP_mult_98_n603), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n604), .ZN(DP_mult_98_n279) );
  XNOR2_X1 DP_mult_98_U453 ( .A(DP_sw0_6_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n602) );
  OAI22_X1 DP_mult_98_U452 ( .A1(DP_mult_98_n602), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n603), .ZN(DP_mult_98_n280) );
  OAI22_X1 DP_mult_98_U451 ( .A1(DP_mult_98_n601), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n602), .ZN(DP_mult_98_n281) );
  XNOR2_X1 DP_mult_98_U450 ( .A(DP_sw0_3_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n599) );
  OAI22_X1 DP_mult_98_U449 ( .A1(DP_mult_98_n599), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n600), .ZN(DP_mult_98_n283) );
  XNOR2_X1 DP_mult_98_U448 ( .A(DP_sw0_2_), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n598) );
  OAI22_X1 DP_mult_98_U447 ( .A1(DP_mult_98_n598), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n599), .ZN(DP_mult_98_n284) );
  XNOR2_X1 DP_mult_98_U446 ( .A(DP_n1), .B(DP_b_int[14]), .ZN(DP_mult_98_n597)
         );
  OAI22_X1 DP_mult_98_U445 ( .A1(DP_mult_98_n597), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n598), .ZN(DP_mult_98_n285) );
  XNOR2_X1 DP_mult_98_U444 ( .A(DP_mult_98_n519), .B(DP_b_int[14]), .ZN(
        DP_mult_98_n595) );
  OAI22_X1 DP_mult_98_U443 ( .A1(DP_mult_98_n595), .A2(DP_mult_98_n596), .B1(
        DP_mult_98_n594), .B2(DP_mult_98_n597), .ZN(DP_mult_98_n286) );
  NOR2_X1 DP_mult_98_U442 ( .A1(DP_mult_98_n561), .A2(DP_mult_98_n594), .ZN(
        DP_mult_98_n287) );
  AOI21_X1 DP_mult_98_U441 ( .B1(DP_mult_98_n580), .B2(DP_mult_98_n578), .A(
        DP_mult_98_n593), .ZN(DP_mult_98_n592) );
  INV_X1 DP_mult_98_U440 ( .A(DP_mult_98_n592), .ZN(DP_mult_98_n288) );
  XNOR2_X1 DP_mult_98_U439 ( .A(DP_sw0_10_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n590) );
  OAI22_X1 DP_mult_98_U438 ( .A1(DP_mult_98_n590), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n591), .ZN(DP_mult_98_n289) );
  XNOR2_X1 DP_mult_98_U437 ( .A(DP_sw0_9_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n589) );
  OAI22_X1 DP_mult_98_U436 ( .A1(DP_mult_98_n589), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n590), .ZN(DP_mult_98_n290) );
  XNOR2_X1 DP_mult_98_U435 ( .A(DP_sw0_8_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n588) );
  OAI22_X1 DP_mult_98_U434 ( .A1(DP_mult_98_n588), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n589), .ZN(DP_mult_98_n291) );
  XNOR2_X1 DP_mult_98_U433 ( .A(DP_sw0_7_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n587) );
  OAI22_X1 DP_mult_98_U432 ( .A1(DP_mult_98_n587), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n588), .ZN(DP_mult_98_n292) );
  XNOR2_X1 DP_mult_98_U431 ( .A(DP_sw0_6_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n586) );
  OAI22_X1 DP_mult_98_U430 ( .A1(DP_mult_98_n586), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n587), .ZN(DP_mult_98_n293) );
  XNOR2_X1 DP_mult_98_U429 ( .A(DP_sw0_5_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n585) );
  OAI22_X1 DP_mult_98_U428 ( .A1(DP_mult_98_n585), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n586), .ZN(DP_mult_98_n294) );
  XNOR2_X1 DP_mult_98_U427 ( .A(DP_sw0_4_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n584) );
  OAI22_X1 DP_mult_98_U426 ( .A1(DP_mult_98_n584), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n585), .ZN(DP_mult_98_n295) );
  XNOR2_X1 DP_mult_98_U425 ( .A(DP_sw0_3_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n583) );
  OAI22_X1 DP_mult_98_U424 ( .A1(DP_mult_98_n583), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n584), .ZN(DP_mult_98_n296) );
  XNOR2_X1 DP_mult_98_U423 ( .A(DP_sw0_2_), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n582) );
  OAI22_X1 DP_mult_98_U422 ( .A1(DP_mult_98_n582), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n583), .ZN(DP_mult_98_n297) );
  XNOR2_X1 DP_mult_98_U421 ( .A(DP_n1), .B(DP_b_int[16]), .ZN(DP_mult_98_n581)
         );
  OAI22_X1 DP_mult_98_U420 ( .A1(DP_mult_98_n581), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n582), .ZN(DP_mult_98_n298) );
  XNOR2_X1 DP_mult_98_U419 ( .A(DP_mult_98_n519), .B(DP_b_int[16]), .ZN(
        DP_mult_98_n579) );
  OAI22_X1 DP_mult_98_U418 ( .A1(DP_mult_98_n579), .A2(DP_mult_98_n580), .B1(
        DP_mult_98_n578), .B2(DP_mult_98_n581), .ZN(DP_mult_98_n299) );
  NOR2_X1 DP_mult_98_U417 ( .A1(DP_mult_98_n561), .A2(DP_mult_98_n578), .ZN(
        DP_mult_98_n300) );
  AOI21_X1 DP_mult_98_U416 ( .B1(DP_mult_98_n564), .B2(DP_mult_98_n562), .A(
        DP_mult_98_n577), .ZN(DP_mult_98_n576) );
  INV_X1 DP_mult_98_U415 ( .A(DP_mult_98_n576), .ZN(DP_mult_98_n301) );
  XNOR2_X1 DP_mult_98_U414 ( .A(DP_sw0_10_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n574) );
  OAI22_X1 DP_mult_98_U413 ( .A1(DP_mult_98_n574), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n575), .ZN(DP_mult_98_n302) );
  OAI22_X1 DP_mult_98_U412 ( .A1(DP_mult_98_n573), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n574), .ZN(DP_mult_98_n303) );
  XNOR2_X1 DP_mult_98_U411 ( .A(DP_sw0_7_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n571) );
  OAI22_X1 DP_mult_98_U410 ( .A1(DP_mult_98_n571), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n572), .ZN(DP_mult_98_n305) );
  XNOR2_X1 DP_mult_98_U409 ( .A(DP_sw0_6_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n570) );
  OAI22_X1 DP_mult_98_U408 ( .A1(DP_mult_98_n570), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n571), .ZN(DP_mult_98_n306) );
  XNOR2_X1 DP_mult_98_U407 ( .A(DP_sw0_5_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n569) );
  OAI22_X1 DP_mult_98_U406 ( .A1(DP_mult_98_n569), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n570), .ZN(DP_mult_98_n307) );
  XNOR2_X1 DP_mult_98_U405 ( .A(DP_sw0_4_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n568) );
  OAI22_X1 DP_mult_98_U404 ( .A1(DP_mult_98_n568), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n569), .ZN(DP_mult_98_n308) );
  XNOR2_X1 DP_mult_98_U403 ( .A(DP_sw0_3_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n567) );
  OAI22_X1 DP_mult_98_U402 ( .A1(DP_mult_98_n567), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n568), .ZN(DP_mult_98_n309) );
  XNOR2_X1 DP_mult_98_U401 ( .A(DP_sw0_2_), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n566) );
  OAI22_X1 DP_mult_98_U400 ( .A1(DP_mult_98_n566), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n567), .ZN(DP_mult_98_n310) );
  XNOR2_X1 DP_mult_98_U399 ( .A(DP_n1), .B(DP_b_int[18]), .ZN(DP_mult_98_n565)
         );
  OAI22_X1 DP_mult_98_U398 ( .A1(DP_mult_98_n565), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n566), .ZN(DP_mult_98_n311) );
  XNOR2_X1 DP_mult_98_U397 ( .A(DP_mult_98_n519), .B(DP_b_int[18]), .ZN(
        DP_mult_98_n563) );
  OAI22_X1 DP_mult_98_U396 ( .A1(DP_mult_98_n563), .A2(DP_mult_98_n564), .B1(
        DP_mult_98_n562), .B2(DP_mult_98_n565), .ZN(DP_mult_98_n312) );
  NOR2_X1 DP_mult_98_U395 ( .A1(DP_mult_98_n561), .A2(DP_mult_98_n562), .ZN(
        DP_mult_98_n313) );
  AOI21_X1 DP_mult_98_U394 ( .B1(DP_mult_98_n546), .B2(DP_mult_98_n547), .A(
        DP_mult_98_n560), .ZN(DP_mult_98_n559) );
  INV_X1 DP_mult_98_U393 ( .A(DP_mult_98_n559), .ZN(DP_mult_98_n314) );
  XNOR2_X1 DP_mult_98_U392 ( .A(DP_sw0_10_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n557) );
  OAI22_X1 DP_mult_98_U391 ( .A1(DP_mult_98_n557), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n558), .ZN(DP_mult_98_n315) );
  XNOR2_X1 DP_mult_98_U390 ( .A(DP_sw0_9_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n556) );
  OAI22_X1 DP_mult_98_U389 ( .A1(DP_mult_98_n556), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n557), .ZN(DP_mult_98_n316) );
  XNOR2_X1 DP_mult_98_U388 ( .A(DP_sw0_8_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n555) );
  OAI22_X1 DP_mult_98_U387 ( .A1(DP_mult_98_n555), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n556), .ZN(DP_mult_98_n317) );
  XNOR2_X1 DP_mult_98_U386 ( .A(DP_sw0_7_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n554) );
  OAI22_X1 DP_mult_98_U385 ( .A1(DP_mult_98_n554), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n555), .ZN(DP_mult_98_n318) );
  XNOR2_X1 DP_mult_98_U384 ( .A(DP_sw0_6_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n553) );
  OAI22_X1 DP_mult_98_U383 ( .A1(DP_mult_98_n553), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n554), .ZN(DP_mult_98_n319) );
  XNOR2_X1 DP_mult_98_U382 ( .A(DP_sw0_5_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n552) );
  OAI22_X1 DP_mult_98_U381 ( .A1(DP_mult_98_n552), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n553), .ZN(DP_mult_98_n320) );
  XNOR2_X1 DP_mult_98_U380 ( .A(DP_sw0_4_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n551) );
  OAI22_X1 DP_mult_98_U379 ( .A1(DP_mult_98_n551), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n552), .ZN(DP_mult_98_n321) );
  XNOR2_X1 DP_mult_98_U378 ( .A(DP_sw0_3_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n550) );
  OAI22_X1 DP_mult_98_U377 ( .A1(DP_mult_98_n550), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n551), .ZN(DP_mult_98_n322) );
  XNOR2_X1 DP_mult_98_U376 ( .A(DP_sw0_2_), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n549) );
  OAI22_X1 DP_mult_98_U375 ( .A1(DP_mult_98_n549), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n550), .ZN(DP_mult_98_n323) );
  XNOR2_X1 DP_mult_98_U374 ( .A(DP_n1), .B(DP_b_int[20]), .ZN(DP_mult_98_n548)
         );
  OAI22_X1 DP_mult_98_U373 ( .A1(DP_mult_98_n548), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n549), .ZN(DP_mult_98_n324) );
  XNOR2_X1 DP_mult_98_U372 ( .A(DP_mult_98_n519), .B(DP_b_int[20]), .ZN(
        DP_mult_98_n545) );
  OAI22_X1 DP_mult_98_U371 ( .A1(DP_mult_98_n545), .A2(DP_mult_98_n546), .B1(
        DP_mult_98_n547), .B2(DP_mult_98_n548), .ZN(DP_mult_98_n325) );
  XOR2_X1 DP_mult_98_U370 ( .A(DP_sw0_12_), .B(DP_mult_98_n544), .Z(
        DP_mult_98_n542) );
  AOI21_X1 DP_mult_98_U369 ( .B1(DP_mult_98_n531), .B2(DP_mult_98_n533), .A(
        DP_mult_98_n542), .ZN(DP_mult_98_n543) );
  INV_X1 DP_mult_98_U368 ( .A(DP_mult_98_n543), .ZN(DP_mult_98_n327) );
  XNOR2_X1 DP_mult_98_U367 ( .A(DP_sw0_11_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n541) );
  OAI22_X1 DP_mult_98_U366 ( .A1(DP_mult_98_n541), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n542), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n328) );
  XNOR2_X1 DP_mult_98_U365 ( .A(DP_sw0_10_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n540) );
  OAI22_X1 DP_mult_98_U364 ( .A1(DP_mult_98_n540), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n541), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n329) );
  XNOR2_X1 DP_mult_98_U363 ( .A(DP_sw0_9_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n539) );
  OAI22_X1 DP_mult_98_U362 ( .A1(DP_mult_98_n539), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n540), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n330) );
  XNOR2_X1 DP_mult_98_U361 ( .A(DP_sw0_8_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n538) );
  OAI22_X1 DP_mult_98_U360 ( .A1(DP_mult_98_n538), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n539), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n331) );
  XNOR2_X1 DP_mult_98_U359 ( .A(DP_sw0_7_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n537) );
  OAI22_X1 DP_mult_98_U358 ( .A1(DP_mult_98_n537), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n538), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n332) );
  XNOR2_X1 DP_mult_98_U357 ( .A(DP_sw0_6_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n536) );
  OAI22_X1 DP_mult_98_U356 ( .A1(DP_mult_98_n536), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n537), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n333) );
  XNOR2_X1 DP_mult_98_U355 ( .A(DP_sw0_5_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n535) );
  OAI22_X1 DP_mult_98_U354 ( .A1(DP_mult_98_n535), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n536), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n334) );
  XNOR2_X1 DP_mult_98_U353 ( .A(DP_sw0_4_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n534) );
  OAI22_X1 DP_mult_98_U352 ( .A1(DP_mult_98_n534), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n535), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n335) );
  XNOR2_X1 DP_mult_98_U351 ( .A(DP_sw0_3_), .B(DP_b_int[22]), .ZN(
        DP_mult_98_n532) );
  OAI22_X1 DP_mult_98_U350 ( .A1(DP_mult_98_n532), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n534), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n336) );
  OAI22_X1 DP_mult_98_U349 ( .A1(DP_mult_98_n530), .A2(DP_mult_98_n531), .B1(
        DP_mult_98_n532), .B2(DP_mult_98_n533), .ZN(DP_mult_98_n337) );
  XNOR2_X1 DP_mult_98_U348 ( .A(DP_sw0_12_), .B(DP_b_int[12]), .ZN(
        DP_mult_98_n528) );
  OAI22_X1 DP_mult_98_U347 ( .A1(DP_mult_98_n529), .A2(DP_mult_98_n526), .B1(
        DP_mult_98_n527), .B2(DP_mult_98_n528), .ZN(DP_mult_98_n520) );
  AOI21_X1 DP_mult_98_U346 ( .B1(DP_mult_98_n526), .B2(DP_mult_98_n527), .A(
        DP_mult_98_n528), .ZN(DP_mult_98_n523) );
  INV_X1 DP_mult_98_U345 ( .A(DP_mult_98_n523), .ZN(DP_mult_98_n521) );
  INV_X1 DP_mult_98_U344 ( .A(DP_mult_98_n520), .ZN(DP_mult_98_n525) );
  AOI222_X1 DP_mult_98_U343 ( .A1(DP_mult_98_n115), .A2(DP_mult_98_n138), .B1(
        DP_mult_98_n525), .B2(DP_mult_98_n115), .C1(DP_mult_98_n525), .C2(
        DP_mult_98_n138), .ZN(DP_mult_98_n524) );
  OAI22_X1 DP_mult_98_U342 ( .A1(DP_mult_98_n523), .A2(DP_mult_98_n524), .B1(
        DP_mult_98_n525), .B2(DP_mult_98_n524), .ZN(DP_mult_98_n522) );
  AOI21_X1 DP_mult_98_U341 ( .B1(DP_mult_98_n520), .B2(DP_mult_98_n521), .A(
        DP_mult_98_n522), .ZN(DP_sw0_b1_11_) );
  XOR2_X2 DP_mult_98_U340 ( .A(DP_b_int[15]), .B(DP_mult_98_n623), .Z(
        DP_mult_98_n594) );
  XOR2_X2 DP_mult_98_U339 ( .A(DP_b_int[17]), .B(DP_mult_98_n621), .Z(
        DP_mult_98_n578) );
  XOR2_X2 DP_mult_98_U338 ( .A(DP_b_int[19]), .B(DP_mult_98_n633), .Z(
        DP_mult_98_n562) );
  XOR2_X2 DP_mult_98_U337 ( .A(DP_b_int[13]), .B(DP_mult_98_n625), .Z(
        DP_mult_98_n527) );
  CLKBUF_X1 DP_mult_98_U336 ( .A(DP_sw0_0_), .Z(DP_mult_98_n519) );
  INV_X1 DP_mult_98_U335 ( .A(DP_b_int[23]), .ZN(DP_mult_98_n533) );
  INV_X1 DP_mult_98_U334 ( .A(DP_mult_98_n654), .ZN(DP_mult_98_n547) );
  HA_X1 DP_mult_98_U120 ( .A(DP_mult_98_n325), .B(DP_mult_98_n337), .CO(
        DP_mult_98_n254), .S(DP_mult_98_n255) );
  FA_X1 DP_mult_98_U119 ( .A(DP_mult_98_n336), .B(DP_mult_98_n313), .CI(
        DP_mult_98_n324), .CO(DP_mult_98_n252), .S(DP_mult_98_n253) );
  HA_X1 DP_mult_98_U118 ( .A(DP_mult_98_n259), .B(DP_mult_98_n312), .CO(
        DP_mult_98_n250), .S(DP_mult_98_n251) );
  FA_X1 DP_mult_98_U117 ( .A(DP_mult_98_n323), .B(DP_mult_98_n335), .CI(
        DP_mult_98_n251), .CO(DP_mult_98_n248), .S(DP_mult_98_n249) );
  FA_X1 DP_mult_98_U109 ( .A(DP_mult_98_n334), .B(DP_mult_98_n300), .CI(
        DP_mult_98_n322), .CO(DP_mult_98_n246), .S(DP_mult_98_n247) );
  FA_X1 DP_mult_98_U108 ( .A(DP_mult_98_n250), .B(DP_mult_98_n311), .CI(
        DP_mult_98_n247), .CO(DP_mult_98_n244), .S(DP_mult_98_n245) );
  HA_X1 DP_mult_98_U107 ( .A(DP_mult_98_n258), .B(DP_mult_98_n299), .CO(
        DP_mult_98_n242), .S(DP_mult_98_n243) );
  FA_X1 DP_mult_98_U106 ( .A(DP_mult_98_n310), .B(DP_mult_98_n333), .CI(
        DP_mult_98_n321), .CO(DP_mult_98_n240), .S(DP_mult_98_n241) );
  FA_X1 DP_mult_98_U105 ( .A(DP_mult_98_n246), .B(DP_mult_98_n243), .CI(
        DP_mult_98_n241), .CO(DP_mult_98_n238), .S(DP_mult_98_n239) );
  FA_X1 DP_mult_98_U104 ( .A(DP_mult_98_n309), .B(DP_mult_98_n287), .CI(
        DP_mult_98_n332), .CO(DP_mult_98_n236), .S(DP_mult_98_n237) );
  FA_X1 DP_mult_98_U103 ( .A(DP_mult_98_n298), .B(DP_mult_98_n320), .CI(
        DP_mult_98_n242), .CO(DP_mult_98_n234), .S(DP_mult_98_n235) );
  FA_X1 DP_mult_98_U102 ( .A(DP_mult_98_n237), .B(DP_mult_98_n240), .CI(
        DP_mult_98_n235), .CO(DP_mult_98_n232), .S(DP_mult_98_n233) );
  HA_X1 DP_mult_98_U101 ( .A(DP_mult_98_n257), .B(DP_mult_98_n286), .CO(
        DP_mult_98_n230), .S(DP_mult_98_n231) );
  FA_X1 DP_mult_98_U100 ( .A(DP_mult_98_n297), .B(DP_mult_98_n308), .CI(
        DP_mult_98_n319), .CO(DP_mult_98_n228), .S(DP_mult_98_n229) );
  FA_X1 DP_mult_98_U99 ( .A(DP_mult_98_n231), .B(DP_mult_98_n331), .CI(
        DP_mult_98_n236), .CO(DP_mult_98_n226), .S(DP_mult_98_n227) );
  FA_X1 DP_mult_98_U98 ( .A(DP_mult_98_n229), .B(DP_mult_98_n234), .CI(
        DP_mult_98_n227), .CO(DP_mult_98_n224), .S(DP_mult_98_n225) );
  FA_X1 DP_mult_98_U97 ( .A(DP_mult_98_n296), .B(DP_mult_98_n274), .CI(
        DP_mult_98_n330), .CO(DP_mult_98_n222), .S(DP_mult_98_n223) );
  FA_X1 DP_mult_98_U96 ( .A(DP_mult_98_n285), .B(DP_mult_98_n318), .CI(
        DP_mult_98_n307), .CO(DP_mult_98_n220), .S(DP_mult_98_n221) );
  FA_X1 DP_mult_98_U95 ( .A(DP_mult_98_n228), .B(DP_mult_98_n230), .CI(
        DP_mult_98_n223), .CO(DP_mult_98_n218), .S(DP_mult_98_n219) );
  FA_X1 DP_mult_98_U94 ( .A(DP_mult_98_n226), .B(DP_mult_98_n221), .CI(
        DP_mult_98_n219), .CO(DP_mult_98_n216), .S(DP_mult_98_n217) );
  HA_X1 DP_mult_98_U93 ( .A(DP_mult_98_n256), .B(DP_mult_98_n273), .CO(
        DP_mult_98_n214), .S(DP_mult_98_n215) );
  FA_X1 DP_mult_98_U92 ( .A(DP_mult_98_n284), .B(DP_mult_98_n306), .CI(
        DP_mult_98_n329), .CO(DP_mult_98_n212), .S(DP_mult_98_n213) );
  FA_X1 DP_mult_98_U91 ( .A(DP_mult_98_n295), .B(DP_mult_98_n317), .CI(
        DP_mult_98_n215), .CO(DP_mult_98_n210), .S(DP_mult_98_n211) );
  FA_X1 DP_mult_98_U90 ( .A(DP_mult_98_n220), .B(DP_mult_98_n222), .CI(
        DP_mult_98_n213), .CO(DP_mult_98_n208), .S(DP_mult_98_n209) );
  FA_X1 DP_mult_98_U89 ( .A(DP_mult_98_n218), .B(DP_mult_98_n211), .CI(
        DP_mult_98_n209), .CO(DP_mult_98_n206), .S(DP_mult_98_n207) );
  HA_X1 DP_mult_98_U88 ( .A(DP_mult_98_n272), .B(DP_mult_98_n283), .CO(
        DP_mult_98_n204), .S(DP_mult_98_n205) );
  FA_X1 DP_mult_98_U87 ( .A(DP_mult_98_n328), .B(DP_mult_98_n305), .CI(
        DP_mult_98_n294), .CO(DP_mult_98_n202), .S(DP_mult_98_n203) );
  FA_X1 DP_mult_98_U86 ( .A(DP_mult_98_n214), .B(DP_mult_98_n316), .CI(
        DP_mult_98_n205), .CO(DP_mult_98_n200), .S(DP_mult_98_n201) );
  FA_X1 DP_mult_98_U85 ( .A(DP_mult_98_n203), .B(DP_mult_98_n212), .CI(
        DP_mult_98_n210), .CO(DP_mult_98_n198), .S(DP_mult_98_n199) );
  FA_X1 DP_mult_98_U84 ( .A(DP_mult_98_n208), .B(DP_mult_98_n201), .CI(
        DP_mult_98_n199), .CO(DP_mult_98_n196), .S(DP_mult_98_n197) );
  FA_X1 DP_mult_98_U81 ( .A(DP_mult_98_n271), .B(DP_mult_98_n293), .CI(
        DP_mult_98_n327), .CO(DP_mult_98_n192), .S(DP_mult_98_n193) );
  FA_X1 DP_mult_98_U80 ( .A(DP_mult_98_n204), .B(DP_mult_98_n315), .CI(
        DP_mult_98_n195), .CO(DP_mult_98_n190), .S(DP_mult_98_n191) );
  FA_X1 DP_mult_98_U79 ( .A(DP_mult_98_n193), .B(DP_mult_98_n202), .CI(
        DP_mult_98_n200), .CO(DP_mult_98_n188), .S(DP_mult_98_n189) );
  FA_X1 DP_mult_98_U78 ( .A(DP_mult_98_n198), .B(DP_mult_98_n191), .CI(
        DP_mult_98_n189), .CO(DP_mult_98_n186), .S(DP_mult_98_n187) );
  FA_X1 DP_mult_98_U76 ( .A(DP_mult_98_n303), .B(DP_mult_98_n281), .CI(
        DP_mult_98_n185), .CO(DP_mult_98_n182), .S(DP_mult_98_n183) );
  FA_X1 DP_mult_98_U75 ( .A(DP_mult_98_n270), .B(DP_mult_98_n292), .CI(
        DP_mult_98_n194), .CO(DP_mult_98_n180), .S(DP_mult_98_n181) );
  FA_X1 DP_mult_98_U74 ( .A(DP_mult_98_n190), .B(DP_mult_98_n192), .CI(
        DP_mult_98_n183), .CO(DP_mult_98_n178), .S(DP_mult_98_n179) );
  FA_X1 DP_mult_98_U73 ( .A(DP_mult_98_n188), .B(DP_mult_98_n181), .CI(
        DP_mult_98_n179), .CO(DP_mult_98_n176), .S(DP_mult_98_n177) );
  FA_X1 DP_mult_98_U72 ( .A(DP_mult_98_n184), .B(DP_mult_98_n269), .CI(
        DP_mult_98_n314), .CO(DP_mult_98_n174), .S(DP_mult_98_n175) );
  FA_X1 DP_mult_98_U71 ( .A(DP_mult_98_n280), .B(DP_mult_98_n302), .CI(
        DP_mult_98_n291), .CO(DP_mult_98_n172), .S(DP_mult_98_n173) );
  FA_X1 DP_mult_98_U70 ( .A(DP_mult_98_n180), .B(DP_mult_98_n182), .CI(
        DP_mult_98_n173), .CO(DP_mult_98_n170), .S(DP_mult_98_n171) );
  FA_X1 DP_mult_98_U69 ( .A(DP_mult_98_n178), .B(DP_mult_98_n175), .CI(
        DP_mult_98_n171), .CO(DP_mult_98_n168), .S(DP_mult_98_n169) );
  FA_X1 DP_mult_98_U67 ( .A(DP_mult_98_n268), .B(DP_mult_98_n279), .CI(
        DP_mult_98_n167), .CO(DP_mult_98_n164), .S(DP_mult_98_n165) );
  FA_X1 DP_mult_98_U66 ( .A(DP_mult_98_n174), .B(DP_mult_98_n290), .CI(
        DP_mult_98_n172), .CO(DP_mult_98_n162), .S(DP_mult_98_n163) );
  FA_X1 DP_mult_98_U65 ( .A(DP_mult_98_n170), .B(DP_mult_98_n165), .CI(
        DP_mult_98_n163), .CO(DP_mult_98_n160), .S(DP_mult_98_n161) );
  FA_X1 DP_mult_98_U64 ( .A(DP_mult_98_n166), .B(DP_mult_98_n267), .CI(
        DP_mult_98_n301), .CO(DP_mult_98_n158), .S(DP_mult_98_n159) );
  FA_X1 DP_mult_98_U63 ( .A(DP_mult_98_n278), .B(DP_mult_98_n289), .CI(
        DP_mult_98_n164), .CO(DP_mult_98_n156), .S(DP_mult_98_n157) );
  FA_X1 DP_mult_98_U62 ( .A(DP_mult_98_n162), .B(DP_mult_98_n159), .CI(
        DP_mult_98_n157), .CO(DP_mult_98_n154), .S(DP_mult_98_n155) );
  FA_X1 DP_mult_98_U60 ( .A(DP_mult_98_n266), .B(DP_mult_98_n277), .CI(
        DP_mult_98_n153), .CO(DP_mult_98_n150), .S(DP_mult_98_n151) );
  FA_X1 DP_mult_98_U59 ( .A(DP_mult_98_n151), .B(DP_mult_98_n158), .CI(
        DP_mult_98_n156), .CO(DP_mult_98_n148), .S(DP_mult_98_n149) );
  FA_X1 DP_mult_98_U58 ( .A(DP_mult_98_n265), .B(DP_mult_98_n152), .CI(
        DP_mult_98_n288), .CO(DP_mult_98_n146), .S(DP_mult_98_n147) );
  FA_X1 DP_mult_98_U57 ( .A(DP_mult_98_n150), .B(DP_mult_98_n276), .CI(
        DP_mult_98_n147), .CO(DP_mult_98_n144), .S(DP_mult_98_n145) );
  FA_X1 DP_mult_98_U55 ( .A(DP_mult_98_n143), .B(DP_mult_98_n264), .CI(
        DP_mult_98_n146), .CO(DP_mult_98_n140), .S(DP_mult_98_n141) );
  FA_X1 DP_mult_98_U54 ( .A(DP_mult_98_n263), .B(DP_mult_98_n142), .CI(
        DP_mult_98_n275), .CO(DP_mult_98_n138), .S(DP_mult_98_n139) );
  FA_X1 DP_mult_98_U42 ( .A(DP_mult_98_n207), .B(DP_mult_98_n216), .CI(
        DP_mult_98_n126), .CO(DP_mult_98_n125), .S(DP_sw0_b1_0_) );
  FA_X1 DP_mult_98_U41 ( .A(DP_mult_98_n197), .B(DP_mult_98_n206), .CI(
        DP_mult_98_n125), .CO(DP_mult_98_n124), .S(DP_sw0_b1_1_) );
  FA_X1 DP_mult_98_U40 ( .A(DP_mult_98_n187), .B(DP_mult_98_n196), .CI(
        DP_mult_98_n124), .CO(DP_mult_98_n123), .S(DP_sw0_b1_2_) );
  FA_X1 DP_mult_98_U39 ( .A(DP_mult_98_n177), .B(DP_mult_98_n186), .CI(
        DP_mult_98_n123), .CO(DP_mult_98_n122), .S(DP_sw0_b1_3_) );
  FA_X1 DP_mult_98_U38 ( .A(DP_mult_98_n169), .B(DP_mult_98_n176), .CI(
        DP_mult_98_n122), .CO(DP_mult_98_n121), .S(DP_sw0_b1_4_) );
  FA_X1 DP_mult_98_U37 ( .A(DP_mult_98_n161), .B(DP_mult_98_n168), .CI(
        DP_mult_98_n121), .CO(DP_mult_98_n120), .S(DP_sw0_b1_5_) );
  FA_X1 DP_mult_98_U36 ( .A(DP_mult_98_n155), .B(DP_mult_98_n160), .CI(
        DP_mult_98_n120), .CO(DP_mult_98_n119), .S(DP_sw0_b1_6_) );
  FA_X1 DP_mult_98_U30 ( .A(DP_mult_98_n149), .B(DP_mult_98_n154), .CI(
        DP_mult_98_n119), .CO(DP_mult_98_n118), .S(DP_sw0_b1_7_) );
  FA_X1 DP_mult_98_U20 ( .A(DP_mult_98_n145), .B(DP_mult_98_n148), .CI(
        DP_mult_98_n118), .CO(DP_mult_98_n117), .S(DP_sw0_b1_8_) );
  FA_X1 DP_mult_98_U10 ( .A(DP_mult_98_n141), .B(DP_mult_98_n144), .CI(
        DP_mult_98_n117), .CO(DP_mult_98_n116), .S(DP_sw0_b1_9_) );
  FA_X1 DP_mult_98_U9 ( .A(DP_mult_98_n140), .B(DP_mult_98_n139), .CI(
        DP_mult_98_n116), .CO(DP_mult_98_n115), .S(DP_sw0_b1_10_) );
  NAND2_X1 DP_mult_97_U971 ( .A1(DP_mult_97_n391), .A2(DP_mult_97_n394), .ZN(
        DP_mult_97_n254) );
  NOR2_X1 DP_mult_97_U970 ( .A1(DP_mult_97_n205), .A2(DP_mult_97_n198), .ZN(
        DP_mult_97_n196) );
  XNOR2_X1 DP_mult_97_U969 ( .A(DP_mult_97_n605), .B(DP_mult_97_n575), .ZN(
        DP_mult_97_n519) );
  XNOR2_X1 DP_mult_97_U968 ( .A(DP_mult_97_n605), .B(DP_mult_97_n576), .ZN(
        DP_mult_97_n520) );
  XNOR2_X1 DP_mult_97_U967 ( .A(DP_mult_97_n605), .B(DP_sw1_1_), .ZN(
        DP_mult_97_n521) );
  XNOR2_X1 DP_mult_97_U966 ( .A(DP_mult_97_n756), .B(DP_mult_97_n670), .ZN(
        DP_mult_97_n515) );
  XNOR2_X1 DP_mult_97_U965 ( .A(DP_mult_97_n756), .B(DP_mult_97_n572), .ZN(
        DP_mult_97_n516) );
  XNOR2_X1 DP_mult_97_U964 ( .A(DP_mult_97_n756), .B(DP_mult_97_n574), .ZN(
        DP_mult_97_n518) );
  NAND2_X1 DP_mult_97_U963 ( .A1(DP_mult_97_n64), .A2(DP_mult_97_n756), .ZN(
        DP_mult_97_n523) );
  XNOR2_X1 DP_mult_97_U962 ( .A(DP_mult_97_n756), .B(DP_sw1_5_), .ZN(
        DP_mult_97_n517) );
  XNOR2_X1 DP_mult_97_U961 ( .A(DP_mult_97_n756), .B(DP_sw1_0_), .ZN(
        DP_mult_97_n522) );
  XNOR2_X1 DP_mult_97_U960 ( .A(DP_mult_97_n756), .B(DP_sw1_8_), .ZN(
        DP_mult_97_n514) );
  XNOR2_X1 DP_mult_97_U959 ( .A(DP_mult_97_n756), .B(DP_sw1_9_), .ZN(
        DP_mult_97_n513) );
  XNOR2_X1 DP_mult_97_U958 ( .A(DP_mult_97_n756), .B(DP_mult_97_n566), .ZN(
        DP_mult_97_n510) );
  XNOR2_X1 DP_mult_97_U957 ( .A(DP_mult_97_n756), .B(DP_mult_97_n567), .ZN(
        DP_mult_97_n511) );
  XNOR2_X1 DP_mult_97_U956 ( .A(DP_mult_97_n756), .B(DP_mult_97_n568), .ZN(
        DP_mult_97_n512) );
  NOR2_X1 DP_mult_97_U955 ( .A1(DP_mult_97_n696), .A2(DP_mult_97_n255), .ZN(
        DP_mult_97_n251) );
  NAND2_X1 DP_mult_97_U954 ( .A1(DP_mult_97_n584), .A2(DP_mult_97_n620), .ZN(
        DP_mult_97_n614) );
  AOI21_X1 DP_mult_97_U953 ( .B1(DP_mult_97_n221), .B2(DP_mult_97_n721), .A(
        DP_mult_97_n218), .ZN(DP_mult_97_n216) );
  XNOR2_X1 DP_mult_97_U952 ( .A(DP_mult_97_n603), .B(DP_sw1_1_), .ZN(
        DP_mult_97_n493) );
  OAI21_X1 DP_mult_97_U951 ( .B1(DP_mult_97_n759), .B2(DP_mult_97_n229), .A(
        DP_mult_97_n226), .ZN(DP_mult_97_n224) );
  NOR2_X1 DP_mult_97_U950 ( .A1(DP_mult_97_n228), .A2(DP_mult_97_n225), .ZN(
        DP_mult_97_n223) );
  NOR2_X1 DP_mult_97_U949 ( .A1(DP_mult_97_n191), .A2(DP_mult_97_n169), .ZN(
        DP_mult_97_n167) );
  XOR2_X1 DP_mult_97_U948 ( .A(DP_a_int[22]), .B(DP_a_int[23]), .Z(
        DP_mult_97_n584) );
  OAI22_X1 DP_mult_97_U947 ( .A1(DP_mult_97_n557), .A2(DP_mult_97_n590), .B1(
        DP_mult_97_n728), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n474) );
  OAI22_X1 DP_mult_97_U946 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n562), .B1(
        DP_mult_97_n561), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n479) );
  OAI22_X1 DP_mult_97_U945 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n560), .B1(
        DP_mult_97_n559), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n477) );
  OAI22_X1 DP_mult_97_U944 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n558), .B1(
        DP_mult_97_n596), .B2(DP_mult_97_n557), .ZN(DP_mult_97_n475) );
  OAI22_X1 DP_mult_97_U943 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n559), .B1(
        DP_mult_97_n558), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n476) );
  OAI22_X1 DP_mult_97_U942 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n553), .B1(
        DP_mult_97_n552), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n470) );
  OAI22_X1 DP_mult_97_U941 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n561), .B1(
        DP_mult_97_n560), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n478) );
  OAI22_X1 DP_mult_97_U940 ( .A1(DP_mult_97_n590), .A2(DP_mult_97_n554), .B1(
        DP_mult_97_n553), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n471) );
  OAI22_X1 DP_mult_97_U939 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n563), .B1(
        DP_mult_97_n562), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n480) );
  OAI22_X1 DP_mult_97_U938 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n555), .B1(
        DP_mult_97_n554), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n472) );
  OAI22_X1 DP_mult_97_U937 ( .A1(DP_mult_97_n762), .A2(DP_mult_97_n728), .B1(
        DP_mult_97_n555), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n473) );
  OAI22_X1 DP_mult_97_U936 ( .A1(DP_mult_97_n677), .A2(DP_mult_97_n564), .B1(
        DP_mult_97_n563), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n481) );
  OAI22_X1 DP_mult_97_U935 ( .A1(DP_mult_97_n677), .A2(DP_mult_97_n602), .B1(
        DP_mult_97_n565), .B2(DP_mult_97_n596), .ZN(DP_mult_97_n403) );
  AOI21_X1 DP_mult_97_U934 ( .B1(DP_mult_97_n193), .B2(DP_mult_97_n185), .A(
        DP_mult_97_n190), .ZN(DP_mult_97_n184) );
  AOI21_X1 DP_mult_97_U933 ( .B1(DP_mult_97_n193), .B2(DP_mult_97_n176), .A(
        DP_mult_97_n177), .ZN(DP_mult_97_n175) );
  AOI21_X1 DP_mult_97_U932 ( .B1(DP_mult_97_n193), .B2(DP_mult_97_n167), .A(
        DP_mult_97_n168), .ZN(DP_mult_97_n166) );
  XNOR2_X1 DP_mult_97_U931 ( .A(DP_mult_97_n193), .B(DP_mult_97_n119), .ZN(
        DP_sw1_a2_5_) );
  AOI21_X1 DP_mult_97_U930 ( .B1(DP_mult_97_n193), .B2(DP_mult_97_n156), .A(
        DP_mult_97_n157), .ZN(DP_mult_97_n155) );
  AOI21_X1 DP_mult_97_U929 ( .B1(DP_mult_97_n193), .B2(DP_mult_97_n147), .A(
        DP_mult_97_n148), .ZN(DP_mult_97_n146) );
  AOI21_X1 DP_mult_97_U928 ( .B1(DP_mult_97_n193), .B2(DP_mult_97_n126), .A(
        DP_mult_97_n127), .ZN(DP_sw1_a2_11_) );
  XNOR2_X1 DP_mult_97_U927 ( .A(DP_mult_97_n606), .B(DP_sw1_9_), .ZN(
        DP_mult_97_n527) );
  XNOR2_X1 DP_mult_97_U926 ( .A(DP_mult_97_n606), .B(DP_sw1_1_), .ZN(
        DP_mult_97_n535) );
  XOR2_X1 DP_mult_97_U925 ( .A(DP_a_int[18]), .B(DP_a_int[19]), .Z(
        DP_mult_97_n582) );
  XNOR2_X1 DP_mult_97_U924 ( .A(DP_a_int[18]), .B(DP_a_int[17]), .ZN(
        DP_mult_97_n617) );
  XNOR2_X1 DP_mult_97_U923 ( .A(DP_mult_97_n603), .B(DP_sw1_5_), .ZN(
        DP_mult_97_n489) );
  XNOR2_X1 DP_mult_97_U922 ( .A(DP_mult_97_n603), .B(DP_mult_97_n575), .ZN(
        DP_mult_97_n491) );
  XNOR2_X1 DP_mult_97_U921 ( .A(DP_mult_97_n603), .B(DP_sw1_0_), .ZN(
        DP_mult_97_n494) );
  XNOR2_X1 DP_mult_97_U920 ( .A(DP_mult_97_n603), .B(DP_mult_97_n576), .ZN(
        DP_mult_97_n492) );
  XNOR2_X1 DP_mult_97_U919 ( .A(DP_mult_97_n753), .B(DP_mult_97_n576), .ZN(
        DP_mult_97_n562) );
  XNOR2_X1 DP_mult_97_U918 ( .A(DP_mult_97_n753), .B(DP_mult_97_n575), .ZN(
        DP_mult_97_n561) );
  XNOR2_X1 DP_mult_97_U917 ( .A(DP_mult_97_n753), .B(DP_mult_97_n566), .ZN(
        DP_mult_97_n552) );
  XNOR2_X1 DP_mult_97_U916 ( .A(DP_mult_97_n608), .B(DP_mult_97_n571), .ZN(
        DP_mult_97_n557) );
  XNOR2_X1 DP_mult_97_U915 ( .A(DP_mult_97_n608), .B(DP_mult_97_n574), .ZN(
        DP_mult_97_n560) );
  XNOR2_X1 DP_mult_97_U914 ( .A(DP_mult_97_n753), .B(DP_sw1_5_), .ZN(
        DP_mult_97_n559) );
  XNOR2_X1 DP_mult_97_U913 ( .A(DP_mult_97_n753), .B(DP_mult_97_n567), .ZN(
        DP_mult_97_n553) );
  XNOR2_X1 DP_mult_97_U912 ( .A(DP_mult_97_n753), .B(DP_mult_97_n572), .ZN(
        DP_mult_97_n558) );
  XNOR2_X1 DP_mult_97_U911 ( .A(DP_mult_97_n753), .B(DP_sw1_1_), .ZN(
        DP_mult_97_n563) );
  XNOR2_X1 DP_mult_97_U910 ( .A(DP_mult_97_n753), .B(DP_mult_97_n568), .ZN(
        DP_mult_97_n554) );
  XNOR2_X1 DP_mult_97_U909 ( .A(DP_mult_97_n753), .B(DP_sw1_9_), .ZN(
        DP_mult_97_n555) );
  XNOR2_X1 DP_mult_97_U908 ( .A(DP_mult_97_n753), .B(DP_mult_97_n733), .ZN(
        DP_mult_97_n564) );
  NAND2_X1 DP_mult_97_U907 ( .A1(DP_mult_97_n82), .A2(DP_mult_97_n753), .ZN(
        DP_mult_97_n565) );
  XOR2_X1 DP_mult_97_U906 ( .A(DP_a_int[15]), .B(DP_a_int[14]), .Z(
        DP_mult_97_n580) );
  XNOR2_X1 DP_mult_97_U905 ( .A(DP_a_int[13]), .B(DP_a_int[14]), .ZN(
        DP_mult_97_n615) );
  XNOR2_X1 DP_mult_97_U904 ( .A(DP_mult_97_n732), .B(DP_mult_97_n574), .ZN(
        DP_mult_97_n504) );
  XNOR2_X1 DP_mult_97_U903 ( .A(DP_mult_97_n604), .B(DP_mult_97_n575), .ZN(
        DP_mult_97_n505) );
  XNOR2_X1 DP_mult_97_U902 ( .A(DP_mult_97_n732), .B(DP_mult_97_n576), .ZN(
        DP_mult_97_n506) );
  XNOR2_X1 DP_mult_97_U901 ( .A(DP_mult_97_n604), .B(DP_sw1_1_), .ZN(
        DP_mult_97_n507) );
  XNOR2_X1 DP_mult_97_U900 ( .A(DP_mult_97_n732), .B(DP_sw1_5_), .ZN(
        DP_mult_97_n503) );
  XNOR2_X1 DP_mult_97_U899 ( .A(DP_mult_97_n732), .B(DP_mult_97_n572), .ZN(
        DP_mult_97_n502) );
  XNOR2_X1 DP_mult_97_U898 ( .A(DP_mult_97_n732), .B(DP_sw1_8_), .ZN(
        DP_mult_97_n500) );
  NAND2_X1 DP_mult_97_U897 ( .A1(DP_mult_97_n35), .A2(DP_mult_97_n732), .ZN(
        DP_mult_97_n509) );
  XNOR2_X1 DP_mult_97_U896 ( .A(DP_mult_97_n732), .B(DP_mult_97_n670), .ZN(
        DP_mult_97_n501) );
  XNOR2_X1 DP_mult_97_U895 ( .A(DP_mult_97_n732), .B(DP_mult_97_n568), .ZN(
        DP_mult_97_n498) );
  XNOR2_X1 DP_mult_97_U894 ( .A(DP_mult_97_n732), .B(DP_sw1_9_), .ZN(
        DP_mult_97_n499) );
  XNOR2_X1 DP_mult_97_U893 ( .A(DP_mult_97_n732), .B(DP_mult_97_n567), .ZN(
        DP_mult_97_n497) );
  XNOR2_X1 DP_mult_97_U892 ( .A(DP_mult_97_n732), .B(DP_mult_97_n566), .ZN(
        DP_mult_97_n496) );
  XNOR2_X1 DP_mult_97_U891 ( .A(DP_mult_97_n603), .B(DP_mult_97_n574), .ZN(
        DP_mult_97_n490) );
  NAND2_X1 DP_mult_97_U890 ( .A1(DP_mult_97_n35), .A2(DP_mult_97_n603), .ZN(
        DP_mult_97_n495) );
  XNOR2_X1 DP_mult_97_U889 ( .A(DP_mult_97_n603), .B(DP_mult_97_n572), .ZN(
        DP_mult_97_n488) );
  XNOR2_X1 DP_mult_97_U888 ( .A(DP_mult_97_n603), .B(DP_sw1_8_), .ZN(
        DP_mult_97_n486) );
  XNOR2_X1 DP_mult_97_U887 ( .A(DP_mult_97_n603), .B(DP_mult_97_n670), .ZN(
        DP_mult_97_n487) );
  XNOR2_X1 DP_mult_97_U886 ( .A(DP_mult_97_n603), .B(DP_sw1_9_), .ZN(
        DP_mult_97_n485) );
  XNOR2_X1 DP_mult_97_U885 ( .A(DP_mult_97_n603), .B(DP_mult_97_n568), .ZN(
        DP_mult_97_n484) );
  XNOR2_X1 DP_mult_97_U884 ( .A(DP_mult_97_n671), .B(DP_mult_97_n567), .ZN(
        DP_mult_97_n483) );
  XNOR2_X1 DP_mult_97_U883 ( .A(DP_mult_97_n671), .B(DP_mult_97_n566), .ZN(
        DP_mult_97_n482) );
  NAND2_X1 DP_mult_97_U882 ( .A1(DP_mult_97_n296), .A2(DP_mult_97_n291), .ZN(
        DP_mult_97_n174) );
  XNOR2_X1 DP_mult_97_U881 ( .A(DP_mult_97_n606), .B(DP_sw1_0_), .ZN(
        DP_mult_97_n536) );
  XNOR2_X1 DP_mult_97_U880 ( .A(DP_mult_97_n606), .B(DP_mult_97_n576), .ZN(
        DP_mult_97_n534) );
  XNOR2_X1 DP_mult_97_U879 ( .A(DP_mult_97_n606), .B(DP_mult_97_n575), .ZN(
        DP_mult_97_n533) );
  XNOR2_X1 DP_mult_97_U878 ( .A(DP_mult_97_n606), .B(DP_sw1_8_), .ZN(
        DP_mult_97_n528) );
  XNOR2_X1 DP_mult_97_U877 ( .A(DP_mult_97_n606), .B(DP_mult_97_n571), .ZN(
        DP_mult_97_n529) );
  XNOR2_X1 DP_mult_97_U876 ( .A(DP_mult_97_n606), .B(DP_sw1_5_), .ZN(
        DP_mult_97_n531) );
  XNOR2_X1 DP_mult_97_U875 ( .A(DP_mult_97_n606), .B(DP_mult_97_n572), .ZN(
        DP_mult_97_n530) );
  XNOR2_X1 DP_mult_97_U874 ( .A(DP_mult_97_n606), .B(DP_mult_97_n568), .ZN(
        DP_mult_97_n526) );
  XNOR2_X1 DP_mult_97_U873 ( .A(DP_mult_97_n606), .B(DP_mult_97_n574), .ZN(
        DP_mult_97_n532) );
  XNOR2_X1 DP_mult_97_U872 ( .A(DP_mult_97_n692), .B(DP_mult_97_n567), .ZN(
        DP_mult_97_n525) );
  XNOR2_X1 DP_mult_97_U871 ( .A(DP_mult_97_n700), .B(DP_mult_97_n566), .ZN(
        DP_mult_97_n524) );
  NAND2_X1 DP_mult_97_U870 ( .A1(DP_mult_97_n692), .A2(DP_mult_97_n82), .ZN(
        DP_mult_97_n537) );
  XNOR2_X1 DP_mult_97_U869 ( .A(DP_mult_97_n709), .B(DP_sw1_0_), .ZN(
        DP_mult_97_n550) );
  XNOR2_X1 DP_mult_97_U868 ( .A(DP_mult_97_n607), .B(DP_mult_97_n572), .ZN(
        DP_mult_97_n544) );
  XNOR2_X1 DP_mult_97_U867 ( .A(DP_mult_97_n607), .B(DP_sw1_5_), .ZN(
        DP_mult_97_n545) );
  XNOR2_X1 DP_mult_97_U866 ( .A(DP_mult_97_n709), .B(DP_sw1_1_), .ZN(
        DP_mult_97_n549) );
  XNOR2_X1 DP_mult_97_U865 ( .A(DP_mult_97_n709), .B(DP_mult_97_n566), .ZN(
        DP_mult_97_n538) );
  XNOR2_X1 DP_mult_97_U864 ( .A(DP_mult_97_n607), .B(DP_mult_97_n574), .ZN(
        DP_mult_97_n546) );
  XNOR2_X1 DP_mult_97_U863 ( .A(DP_mult_97_n709), .B(DP_mult_97_n567), .ZN(
        DP_mult_97_n539) );
  XNOR2_X1 DP_mult_97_U862 ( .A(DP_mult_97_n709), .B(DP_mult_97_n575), .ZN(
        DP_mult_97_n547) );
  XNOR2_X1 DP_mult_97_U861 ( .A(DP_mult_97_n709), .B(DP_mult_97_n576), .ZN(
        DP_mult_97_n548) );
  XNOR2_X1 DP_mult_97_U860 ( .A(DP_mult_97_n709), .B(DP_mult_97_n568), .ZN(
        DP_mult_97_n540) );
  XNOR2_X1 DP_mult_97_U859 ( .A(DP_mult_97_n709), .B(DP_mult_97_n670), .ZN(
        DP_mult_97_n543) );
  XNOR2_X1 DP_mult_97_U858 ( .A(DP_mult_97_n607), .B(DP_sw1_8_), .ZN(
        DP_mult_97_n542) );
  XNOR2_X1 DP_mult_97_U857 ( .A(DP_mult_97_n709), .B(DP_sw1_9_), .ZN(
        DP_mult_97_n541) );
  NAND2_X1 DP_mult_97_U856 ( .A1(DP_mult_97_n98), .A2(DP_mult_97_n709), .ZN(
        DP_mult_97_n551) );
  NOR2_X1 DP_mult_97_U855 ( .A1(DP_mult_97_n397), .A2(DP_mult_97_n402), .ZN(
        DP_mult_97_n258) );
  NAND2_X1 DP_mult_97_U854 ( .A1(DP_mult_97_n397), .A2(DP_mult_97_n402), .ZN(
        DP_mult_97_n259) );
  INV_X1 DP_mult_97_U853 ( .A(DP_mult_97_n222), .ZN(DP_mult_97_n221) );
  AOI21_X1 DP_mult_97_U852 ( .B1(DP_mult_97_n768), .B2(DP_mult_97_n208), .A(
        DP_mult_97_n209), .ZN(DP_mult_97_n207) );
  AOI21_X1 DP_mult_97_U851 ( .B1(DP_mult_97_n201), .B2(DP_mult_97_n661), .A(
        DP_mult_97_n202), .ZN(DP_mult_97_n200) );
  NAND2_X1 DP_mult_97_U850 ( .A1(DP_mult_97_n583), .A2(DP_mult_97_n619), .ZN(
        DP_mult_97_n613) );
  OAI22_X1 DP_mult_97_U849 ( .A1(DP_mult_97_n589), .A2(DP_mult_97_n545), .B1(
        DP_mult_97_n544), .B2(DP_mult_97_n595), .ZN(DP_mult_97_n462) );
  OAI22_X1 DP_mult_97_U848 ( .A1(DP_mult_97_n698), .A2(DP_mult_97_n550), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n549), .ZN(DP_mult_97_n467) );
  OAI22_X1 DP_mult_97_U847 ( .A1(DP_mult_97_n699), .A2(DP_mult_97_n539), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n538), .ZN(DP_mult_97_n326) );
  OAI22_X1 DP_mult_97_U846 ( .A1(DP_mult_97_n546), .A2(DP_mult_97_n589), .B1(
        DP_mult_97_n595), .B2(DP_mult_97_n545), .ZN(DP_mult_97_n463) );
  OAI22_X1 DP_mult_97_U845 ( .A1(DP_mult_97_n698), .A2(DP_mult_97_n547), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n546), .ZN(DP_mult_97_n464) );
  OAI22_X1 DP_mult_97_U844 ( .A1(DP_mult_97_n699), .A2(DP_mult_97_n549), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n548), .ZN(DP_mult_97_n466) );
  OAI22_X1 DP_mult_97_U843 ( .A1(DP_mult_97_n698), .A2(DP_mult_97_n548), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n547), .ZN(DP_mult_97_n465) );
  OAI22_X1 DP_mult_97_U842 ( .A1(DP_mult_97_n699), .A2(DP_mult_97_n540), .B1(
        DP_mult_97_n595), .B2(DP_mult_97_n539), .ZN(DP_mult_97_n457) );
  OAI22_X1 DP_mult_97_U841 ( .A1(DP_mult_97_n699), .A2(DP_mult_97_n544), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n543), .ZN(DP_mult_97_n461) );
  OAI22_X1 DP_mult_97_U840 ( .A1(DP_mult_97_n698), .A2(DP_mult_97_n543), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n542), .ZN(DP_mult_97_n460) );
  OAI22_X1 DP_mult_97_U839 ( .A1(DP_mult_97_n699), .A2(DP_mult_97_n541), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n540), .ZN(DP_mult_97_n458) );
  OAI22_X1 DP_mult_97_U838 ( .A1(DP_mult_97_n698), .A2(DP_mult_97_n542), .B1(
        DP_mult_97_n693), .B2(DP_mult_97_n541), .ZN(DP_mult_97_n459) );
  OAI22_X1 DP_mult_97_U837 ( .A1(DP_mult_97_n699), .A2(DP_mult_97_n601), .B1(
        DP_mult_97_n551), .B2(DP_mult_97_n693), .ZN(DP_mult_97_n402) );
  OAI22_X1 DP_mult_97_U836 ( .A1(DP_mult_97_n508), .A2(DP_mult_97_n610), .B1(
        DP_mult_97_n507), .B2(DP_mult_97_n592), .ZN(DP_mult_97_n428) );
  NAND2_X1 DP_mult_97_U835 ( .A1(DP_mult_97_n580), .A2(DP_mult_97_n616), .ZN(
        DP_mult_97_n610) );
  NAND2_X1 DP_mult_97_U834 ( .A1(DP_mult_97_n581), .A2(DP_mult_97_n617), .ZN(
        DP_mult_97_n611) );
  INV_X1 DP_mult_97_U833 ( .A(DP_mult_97_n688), .ZN(DP_mult_97_n230) );
  OAI21_X1 DP_mult_97_U832 ( .B1(DP_mult_97_n230), .B2(DP_mult_97_n228), .A(
        DP_mult_97_n722), .ZN(DP_mult_97_n227) );
  XOR2_X1 DP_mult_97_U831 ( .A(DP_a_int[20]), .B(DP_a_int[21]), .Z(
        DP_mult_97_n583) );
  XNOR2_X1 DP_mult_97_U830 ( .A(DP_a_int[20]), .B(DP_a_int[19]), .ZN(
        DP_mult_97_n618) );
  NAND2_X1 DP_mult_97_U829 ( .A1(DP_mult_97_n579), .A2(DP_mult_97_n615), .ZN(
        DP_mult_97_n609) );
  NAND2_X1 DP_mult_97_U828 ( .A1(DP_mult_97_n196), .A2(DP_mult_97_n212), .ZN(
        DP_mult_97_n194) );
  AOI21_X1 DP_mult_97_U827 ( .B1(DP_mult_97_n213), .B2(DP_mult_97_n196), .A(
        DP_mult_97_n197), .ZN(DP_mult_97_n195) );
  XOR2_X1 DP_mult_97_U826 ( .A(DP_mult_97_n184), .B(DP_mult_97_n118), .Z(
        DP_sw1_a2_6_) );
  XNOR2_X1 DP_mult_97_U825 ( .A(DP_a_int[21]), .B(DP_a_int[22]), .ZN(
        DP_mult_97_n619) );
  OAI22_X1 DP_mult_97_U824 ( .A1(DP_mult_97_n520), .A2(DP_mult_97_n587), .B1(
        DP_mult_97_n519), .B2(DP_mult_97_n593), .ZN(DP_mult_97_n439) );
  NOR2_X1 DP_mult_97_U823 ( .A1(DP_mult_97_n391), .A2(DP_mult_97_n394), .ZN(
        DP_mult_97_n253) );
  NOR2_X1 DP_mult_97_U822 ( .A1(DP_mult_97_n395), .A2(DP_mult_97_n743), .ZN(
        DP_mult_97_n255) );
  INV_X1 DP_mult_97_U821 ( .A(DP_mult_97_n726), .ZN(DP_mult_97_n769) );
  OR2_X1 DP_mult_97_U820 ( .A1(DP_mult_97_n413), .A2(DP_mult_97_n669), .ZN(
        DP_mult_97_n336) );
  XNOR2_X1 DP_mult_97_U819 ( .A(DP_mult_97_n413), .B(DP_mult_97_n669), .ZN(
        DP_mult_97_n337) );
  OAI21_X1 DP_mult_97_U818 ( .B1(DP_mult_97_n198), .B2(DP_mult_97_n206), .A(
        DP_mult_97_n199), .ZN(DP_mult_97_n197) );
  NOR2_X1 DP_mult_97_U817 ( .A1(DP_mult_97_n219), .A2(DP_mult_97_n214), .ZN(
        DP_mult_97_n212) );
  OAI22_X1 DP_mult_97_U816 ( .A1(DP_mult_97_n587), .A2(DP_mult_97_n521), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n520), .ZN(DP_mult_97_n440) );
  OAI22_X1 DP_mult_97_U815 ( .A1(DP_mult_97_n758), .A2(DP_mult_97_n599), .B1(
        DP_mult_97_n523), .B2(DP_mult_97_n754), .ZN(DP_mult_97_n400) );
  OAI22_X1 DP_mult_97_U814 ( .A1(DP_mult_97_n758), .A2(DP_mult_97_n522), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n521), .ZN(DP_mult_97_n441) );
  OAI22_X1 DP_mult_97_U813 ( .A1(DP_mult_97_n757), .A2(DP_mult_97_n519), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n518), .ZN(DP_mult_97_n438) );
  OAI22_X1 DP_mult_97_U812 ( .A1(DP_mult_97_n758), .A2(DP_mult_97_n517), .B1(
        DP_mult_97_n593), .B2(DP_mult_97_n516), .ZN(DP_mult_97_n436) );
  OAI22_X1 DP_mult_97_U811 ( .A1(DP_mult_97_n757), .A2(DP_mult_97_n516), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n515), .ZN(DP_mult_97_n435) );
  OAI22_X1 DP_mult_97_U810 ( .A1(DP_mult_97_n511), .A2(DP_mult_97_n758), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n510), .ZN(DP_mult_97_n294) );
  OAI22_X1 DP_mult_97_U809 ( .A1(DP_mult_97_n757), .A2(DP_mult_97_n518), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n517), .ZN(DP_mult_97_n437) );
  OAI22_X1 DP_mult_97_U808 ( .A1(DP_mult_97_n757), .A2(DP_mult_97_n515), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n514), .ZN(DP_mult_97_n434) );
  OAI22_X1 DP_mult_97_U807 ( .A1(DP_mult_97_n758), .A2(DP_mult_97_n512), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n511), .ZN(DP_mult_97_n431) );
  OAI22_X1 DP_mult_97_U806 ( .A1(DP_mult_97_n758), .A2(DP_mult_97_n513), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n512), .ZN(DP_mult_97_n432) );
  OAI22_X1 DP_mult_97_U805 ( .A1(DP_mult_97_n757), .A2(DP_mult_97_n514), .B1(
        DP_mult_97_n754), .B2(DP_mult_97_n513), .ZN(DP_mult_97_n433) );
  NAND2_X1 DP_mult_97_U804 ( .A1(DP_mult_97_n760), .A2(DP_mult_97_n746), .ZN(
        DP_mult_97_n232) );
  AOI21_X1 DP_mult_97_U803 ( .B1(DP_mult_97_n695), .B2(DP_mult_97_n744), .A(
        DP_mult_97_n741), .ZN(DP_mult_97_n233) );
  NAND2_X1 DP_mult_97_U802 ( .A1(DP_mult_97_n349), .A2(DP_mult_97_n358), .ZN(
        DP_mult_97_n226) );
  XOR2_X1 DP_mult_97_U801 ( .A(DP_mult_97_n200), .B(DP_mult_97_n120), .Z(
        DP_sw1_a2_4_) );
  OAI21_X1 DP_mult_97_U800 ( .B1(DP_mult_97_n250), .B2(DP_mult_97_n248), .A(
        DP_mult_97_n249), .ZN(DP_mult_97_n247) );
  AOI21_X1 DP_mult_97_U799 ( .B1(DP_mult_97_n251), .B2(DP_mult_97_n257), .A(
        DP_mult_97_n252), .ZN(DP_mult_97_n250) );
  XNOR2_X1 DP_mult_97_U798 ( .A(DP_a_int[16]), .B(DP_a_int[15]), .ZN(
        DP_mult_97_n616) );
  XOR2_X1 DP_mult_97_U797 ( .A(DP_a_int[16]), .B(DP_a_int[17]), .Z(
        DP_mult_97_n581) );
  OAI22_X1 DP_mult_97_U796 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n503), .B1(
        DP_mult_97_n690), .B2(DP_mult_97_n502), .ZN(DP_mult_97_n423) );
  OAI22_X1 DP_mult_97_U795 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n501), .B1(
        DP_mult_97_n678), .B2(DP_mult_97_n500), .ZN(DP_mult_97_n421) );
  OAI22_X1 DP_mult_97_U794 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n499), .B1(
        DP_mult_97_n678), .B2(DP_mult_97_n498), .ZN(DP_mult_97_n419) );
  OAI22_X1 DP_mult_97_U793 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n500), .B1(
        DP_mult_97_n690), .B2(DP_mult_97_n499), .ZN(DP_mult_97_n420) );
  OAI22_X1 DP_mult_97_U792 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n498), .B1(
        DP_mult_97_n690), .B2(DP_mult_97_n497), .ZN(DP_mult_97_n418) );
  OAI22_X1 DP_mult_97_U791 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n497), .B1(
        DP_mult_97_n690), .B2(DP_mult_97_n496), .ZN(DP_mult_97_n284) );
  OAI22_X1 DP_mult_97_U790 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n502), .B1(
        DP_mult_97_n690), .B2(DP_mult_97_n501), .ZN(DP_mult_97_n422) );
  INV_X1 DP_mult_97_U789 ( .A(DP_sw1_0_), .ZN(DP_mult_97_n64) );
  INV_X1 DP_mult_97_U788 ( .A(DP_sw1_0_), .ZN(DP_mult_97_n35) );
  INV_X1 DP_mult_97_U787 ( .A(DP_sw1_0_), .ZN(DP_mult_97_n82) );
  INV_X1 DP_mult_97_U786 ( .A(DP_sw1_0_), .ZN(DP_mult_97_n98) );
  OAI21_X1 DP_mult_97_U785 ( .B1(DP_mult_97_n214), .B2(DP_mult_97_n220), .A(
        DP_mult_97_n215), .ZN(DP_mult_97_n213) );
  INV_X1 DP_mult_97_U784 ( .A(DP_mult_97_n98), .ZN(DP_mult_97_n767) );
  OAI22_X1 DP_mult_97_U783 ( .A1(DP_mult_97_n506), .A2(DP_mult_97_n755), .B1(
        DP_mult_97_n592), .B2(DP_mult_97_n505), .ZN(DP_mult_97_n426) );
  OAI22_X1 DP_mult_97_U782 ( .A1(DP_mult_97_n755), .A2(DP_mult_97_n507), .B1(
        DP_mult_97_n689), .B2(DP_mult_97_n506), .ZN(DP_mult_97_n427) );
  BUF_X2 DP_mult_97_U781 ( .A(DP_sw1_2_), .Z(DP_mult_97_n576) );
  NOR2_X1 DP_mult_97_U780 ( .A1(DP_mult_97_n319), .A2(DP_mult_97_n328), .ZN(
        DP_mult_97_n205) );
  OAI22_X1 DP_mult_97_U779 ( .A1(DP_mult_97_n710), .A2(DP_mult_97_n530), .B1(
        DP_mult_97_n529), .B2(DP_mult_97_n594), .ZN(DP_mult_97_n448) );
  OAI22_X1 DP_mult_97_U778 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n532), .B1(
        DP_mult_97_n681), .B2(DP_mult_97_n531), .ZN(DP_mult_97_n450) );
  OAI22_X1 DP_mult_97_U777 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n535), .B1(
        DP_mult_97_n682), .B2(DP_mult_97_n534), .ZN(DP_mult_97_n453) );
  OAI22_X1 DP_mult_97_U776 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n531), .B1(
        DP_mult_97_n682), .B2(DP_mult_97_n530), .ZN(DP_mult_97_n449) );
  OAI22_X1 DP_mult_97_U775 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n536), .B1(
        DP_mult_97_n682), .B2(DP_mult_97_n535), .ZN(DP_mult_97_n454) );
  OAI22_X1 DP_mult_97_U774 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n528), .B1(
        DP_mult_97_n681), .B2(DP_mult_97_n527), .ZN(DP_mult_97_n446) );
  OAI22_X1 DP_mult_97_U773 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n534), .B1(
        DP_mult_97_n681), .B2(DP_mult_97_n533), .ZN(DP_mult_97_n452) );
  OAI22_X1 DP_mult_97_U772 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n704), .B1(
        DP_mult_97_n682), .B2(DP_mult_97_n528), .ZN(DP_mult_97_n447) );
  OAI22_X1 DP_mult_97_U771 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n527), .B1(
        DP_mult_97_n681), .B2(DP_mult_97_n526), .ZN(DP_mult_97_n445) );
  OAI22_X1 DP_mult_97_U770 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n525), .B1(
        DP_mult_97_n524), .B2(DP_mult_97_n681), .ZN(DP_mult_97_n308) );
  OAI22_X1 DP_mult_97_U769 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n526), .B1(
        DP_mult_97_n681), .B2(DP_mult_97_n525), .ZN(DP_mult_97_n444) );
  OAI22_X1 DP_mult_97_U768 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n533), .B1(
        DP_mult_97_n682), .B2(DP_mult_97_n532), .ZN(DP_mult_97_n451) );
  OAI22_X1 DP_mult_97_U767 ( .A1(DP_mult_97_n711), .A2(DP_mult_97_n600), .B1(
        DP_mult_97_n537), .B2(DP_mult_97_n682), .ZN(DP_mult_97_n401) );
  BUF_X2 DP_mult_97_U766 ( .A(DP_sw1_3_), .Z(DP_mult_97_n575) );
  XNOR2_X1 DP_mult_97_U765 ( .A(DP_mult_97_n227), .B(DP_mult_97_n124), .ZN(
        DP_sw1_a2_0_) );
  INV_X1 DP_mult_97_U764 ( .A(DP_mult_97_n213), .ZN(DP_mult_97_n211) );
  OAI21_X1 DP_mult_97_U763 ( .B1(DP_mult_97_n211), .B2(DP_mult_97_n203), .A(
        DP_mult_97_n206), .ZN(DP_mult_97_n202) );
  INV_X1 DP_mult_97_U762 ( .A(DP_mult_97_n211), .ZN(DP_mult_97_n209) );
  NOR2_X1 DP_mult_97_U761 ( .A1(DP_mult_97_n359), .A2(DP_mult_97_n366), .ZN(
        DP_mult_97_n228) );
  NAND2_X1 DP_mult_97_U760 ( .A1(DP_mult_97_n359), .A2(DP_mult_97_n366), .ZN(
        DP_mult_97_n229) );
  OAI22_X1 DP_mult_97_U759 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n492), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n491), .ZN(DP_mult_97_n413) );
  OAI22_X1 DP_mult_97_U758 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n493), .B1(
        DP_mult_97_n492), .B2(DP_mult_97_n591), .ZN(DP_mult_97_n414) );
  OAI22_X1 DP_mult_97_U757 ( .A1(DP_mult_97_n585), .A2(DP_mult_97_n597), .B1(
        DP_mult_97_n495), .B2(DP_mult_97_n591), .ZN(DP_mult_97_n398) );
  OAI22_X1 DP_mult_97_U756 ( .A1(DP_mult_97_n585), .A2(DP_mult_97_n494), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n493), .ZN(DP_mult_97_n415) );
  NAND2_X1 DP_mult_97_U755 ( .A1(DP_mult_97_n387), .A2(DP_mult_97_n390), .ZN(
        DP_mult_97_n249) );
  NOR2_X1 DP_mult_97_U754 ( .A1(DP_mult_97_n387), .A2(DP_mult_97_n390), .ZN(
        DP_mult_97_n248) );
  INV_X1 DP_mult_97_U753 ( .A(DP_mult_97_n212), .ZN(DP_mult_97_n210) );
  OAI22_X1 DP_mult_97_U752 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n486), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n485), .ZN(DP_mult_97_n407) );
  OAI22_X1 DP_mult_97_U751 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n485), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n484), .ZN(DP_mult_97_n406) );
  OAI22_X1 DP_mult_97_U750 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n484), .B1(
        DP_mult_97_n676), .B2(DP_mult_97_n483), .ZN(DP_mult_97_n405) );
  OAI22_X1 DP_mult_97_U749 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n483), .B1(
        DP_mult_97_n687), .B2(DP_mult_97_n482), .ZN(DP_mult_97_n278) );
  NAND3_X1 DP_mult_97_U748 ( .A1(DP_mult_97_n764), .A2(DP_mult_97_n765), .A3(
        DP_mult_97_n766), .ZN(DP_mult_97_n374) );
  NAND2_X1 DP_mult_97_U747 ( .A1(DP_mult_97_n379), .A2(DP_mult_97_n742), .ZN(
        DP_mult_97_n766) );
  NAND2_X1 DP_mult_97_U746 ( .A1(DP_mult_97_n380), .A2(DP_mult_97_n742), .ZN(
        DP_mult_97_n765) );
  NAND2_X1 DP_mult_97_U745 ( .A1(DP_mult_97_n380), .A2(DP_mult_97_n379), .ZN(
        DP_mult_97_n764) );
  XOR2_X1 DP_mult_97_U744 ( .A(DP_mult_97_n380), .B(DP_mult_97_n763), .Z(
        DP_mult_97_n375) );
  XOR2_X1 DP_mult_97_U743 ( .A(DP_mult_97_n379), .B(DP_mult_97_n742), .Z(
        DP_mult_97_n763) );
  INV_X1 DP_mult_97_U742 ( .A(DP_mult_97_n762), .ZN(DP_mult_97_n103) );
  INV_X1 DP_mult_97_U741 ( .A(DP_mult_97_n308), .ZN(DP_mult_97_n309) );
  INV_X1 DP_mult_97_U740 ( .A(DP_mult_97_n754), .ZN(DP_mult_97_n47) );
  BUF_X2 DP_mult_97_U739 ( .A(DP_sw1_6_), .Z(DP_mult_97_n572) );
  OAI22_X1 DP_mult_97_U738 ( .A1(DP_mult_97_n755), .A2(DP_mult_97_n505), .B1(
        DP_mult_97_n689), .B2(DP_mult_97_n504), .ZN(DP_mult_97_n425) );
  OAI22_X1 DP_mult_97_U737 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n712), .B1(
        DP_mult_97_n509), .B2(DP_mult_97_n678), .ZN(DP_mult_97_n399) );
  INV_X1 DP_mult_97_U736 ( .A(DP_mult_97_n691), .ZN(DP_mult_97_n24) );
  OR2_X1 DP_mult_97_U735 ( .A1(DP_mult_97_n358), .A2(DP_mult_97_n697), .ZN(
        DP_mult_97_n761) );
  INV_X1 DP_mult_97_U734 ( .A(DP_mult_97_n690), .ZN(DP_mult_97_n30) );
  OR2_X1 DP_mult_97_U733 ( .A1(DP_mult_97_n374), .A2(DP_mult_97_n367), .ZN(
        DP_mult_97_n760) );
  NOR2_X1 DP_mult_97_U732 ( .A1(DP_mult_97_n358), .A2(DP_mult_97_n349), .ZN(
        DP_mult_97_n225) );
  NAND2_X1 DP_mult_97_U731 ( .A1(DP_mult_97_n226), .A2(DP_mult_97_n761), .ZN(
        DP_mult_97_n124) );
  NOR2_X1 DP_mult_97_U730 ( .A1(DP_mult_97_n349), .A2(DP_mult_97_n358), .ZN(
        DP_mult_97_n759) );
  INV_X1 DP_mult_97_U729 ( .A(DP_mult_97_n710), .ZN(DP_mult_97_n69) );
  OAI21_X1 DP_mult_97_U728 ( .B1(DP_mult_97_n253), .B2(DP_mult_97_n256), .A(
        DP_mult_97_n254), .ZN(DP_mult_97_n252) );
  INV_X1 DP_mult_97_U727 ( .A(DP_mult_97_n757), .ZN(DP_mult_97_n40) );
  INV_X1 DP_mult_97_U726 ( .A(DP_mult_97_n756), .ZN(DP_mult_97_n599) );
  INV_X1 DP_mult_97_U725 ( .A(DP_mult_97_n682), .ZN(DP_mult_97_n77) );
  AOI21_X1 DP_mult_97_U724 ( .B1(DP_mult_97_n247), .B2(DP_mult_97_n745), .A(
        DP_mult_97_n747), .ZN(DP_mult_97_n242) );
  OAI22_X1 DP_mult_97_U723 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n490), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n489), .ZN(DP_mult_97_n411) );
  OAI22_X1 DP_mult_97_U722 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n489), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n488), .ZN(DP_mult_97_n410) );
  OAI22_X1 DP_mult_97_U721 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n491), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n490), .ZN(DP_mult_97_n412) );
  OAI22_X1 DP_mult_97_U720 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n487), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n486), .ZN(DP_mult_97_n408) );
  OAI22_X1 DP_mult_97_U719 ( .A1(DP_mult_97_n727), .A2(DP_mult_97_n488), .B1(
        DP_mult_97_n591), .B2(DP_mult_97_n487), .ZN(DP_mult_97_n409) );
  INV_X1 DP_mult_97_U718 ( .A(DP_mult_97_n727), .ZN(DP_mult_97_n8) );
  INV_X1 DP_mult_97_U717 ( .A(DP_mult_97_n693), .ZN(DP_mult_97_n88) );
  BUF_X1 DP_mult_97_U716 ( .A(DP_mult_97_n614), .Z(DP_mult_97_n590) );
  INV_X1 DP_mult_97_U715 ( .A(DP_mult_97_n326), .ZN(DP_mult_97_n327) );
  NAND2_X1 DP_mult_97_U714 ( .A1(DP_mult_97_n311), .A2(DP_mult_97_n318), .ZN(
        DP_mult_97_n199) );
  INV_X1 DP_mult_97_U713 ( .A(DP_a_int[23]), .ZN(DP_mult_97_n620) );
  BUF_X2 DP_mult_97_U712 ( .A(DP_sw1_11_), .Z(DP_mult_97_n567) );
  BUF_X2 DP_mult_97_U711 ( .A(DP_sw1_10_), .Z(DP_mult_97_n568) );
  BUF_X2 DP_mult_97_U710 ( .A(DP_sw1_12_), .Z(DP_mult_97_n566) );
  BUF_X2 DP_mult_97_U709 ( .A(DP_sw1_4_), .Z(DP_mult_97_n574) );
  XOR2_X1 DP_mult_97_U708 ( .A(DP_a_int[13]), .B(DP_a_int[12]), .Z(
        DP_mult_97_n579) );
  CLKBUF_X3 DP_mult_97_U707 ( .A(DP_a_int[12]), .Z(DP_mult_97_n603) );
  AND2_X1 DP_mult_97_U706 ( .A1(DP_mult_97_n733), .A2(DP_mult_97_n88), .ZN(
        DP_mult_97_n752) );
  INV_X1 DP_mult_97_U705 ( .A(DP_mult_97_n687), .ZN(DP_mult_97_n9) );
  INV_X1 DP_mult_97_U704 ( .A(DP_mult_97_n482), .ZN(DP_mult_97_n10) );
  INV_X1 DP_mult_97_U703 ( .A(DP_mult_97_n603), .ZN(DP_mult_97_n597) );
  INV_X1 DP_mult_97_U702 ( .A(DP_mult_97_n606), .ZN(DP_mult_97_n600) );
  INV_X1 DP_mult_97_U701 ( .A(DP_mult_97_n698), .ZN(DP_mult_97_n87) );
  AND2_X1 DP_mult_97_U700 ( .A1(DP_mult_97_n752), .A2(DP_mult_97_n480), .ZN(
        DP_mult_97_n751) );
  OR2_X1 DP_mult_97_U699 ( .A1(DP_mult_97_n752), .A2(DP_mult_97_n480), .ZN(
        DP_mult_97_n750) );
  AND2_X1 DP_mult_97_U698 ( .A1(DP_mult_97_n403), .A2(DP_mult_97_n481), .ZN(
        DP_mult_97_n749) );
  INV_X1 DP_mult_97_U697 ( .A(DP_mult_97_n608), .ZN(DP_mult_97_n602) );
  AOI21_X1 DP_mult_97_U696 ( .B1(DP_mult_97_n750), .B2(DP_mult_97_n749), .A(
        DP_mult_97_n751), .ZN(DP_mult_97_n260) );
  OAI21_X1 DP_mult_97_U695 ( .B1(DP_mult_97_n260), .B2(DP_mult_97_n258), .A(
        DP_mult_97_n259), .ZN(DP_mult_97_n257) );
  AND2_X1 DP_mult_97_U694 ( .A1(DP_mult_97_n767), .A2(DP_mult_97_n47), .ZN(
        DP_mult_97_n748) );
  BUF_X1 DP_mult_97_U693 ( .A(DP_mult_97_n611), .Z(DP_mult_97_n758) );
  INV_X1 DP_mult_97_U692 ( .A(DP_mult_97_n294), .ZN(DP_mult_97_n295) );
  INV_X1 DP_mult_97_U691 ( .A(DP_mult_97_n284), .ZN(DP_mult_97_n285) );
  OAI21_X1 DP_mult_97_U690 ( .B1(DP_mult_97_n24), .B2(DP_mult_97_n30), .A(
        DP_mult_97_n26), .ZN(DP_mult_97_n417) );
  INV_X1 DP_mult_97_U689 ( .A(DP_mult_97_n709), .ZN(DP_mult_97_n601) );
  INV_X1 DP_mult_97_U688 ( .A(DP_mult_97_n496), .ZN(DP_mult_97_n26) );
  NAND2_X1 DP_mult_97_U687 ( .A1(DP_mult_97_n404), .A2(DP_mult_97_n278), .ZN(
        DP_mult_97_n129) );
  INV_X1 DP_mult_97_U686 ( .A(DP_mult_97_n278), .ZN(DP_mult_97_n279) );
  AND2_X1 DP_mult_97_U685 ( .A1(DP_mult_97_n381), .A2(DP_mult_97_n386), .ZN(
        DP_mult_97_n747) );
  INV_X1 DP_mult_97_U684 ( .A(DP_mult_97_n596), .ZN(DP_mult_97_n104) );
  OR2_X1 DP_mult_97_U683 ( .A1(DP_mult_97_n375), .A2(DP_mult_97_n377), .ZN(
        DP_mult_97_n746) );
  OR2_X1 DP_mult_97_U682 ( .A1(DP_mult_97_n381), .A2(DP_mult_97_n386), .ZN(
        DP_mult_97_n745) );
  AND2_X1 DP_mult_97_U681 ( .A1(DP_mult_97_n375), .A2(DP_mult_97_n377), .ZN(
        DP_mult_97_n744) );
  AND2_X1 DP_mult_97_U680 ( .A1(DP_mult_97_n767), .A2(DP_mult_97_n77), .ZN(
        DP_mult_97_n743) );
  INV_X1 DP_mult_97_U679 ( .A(DP_mult_97_n538), .ZN(DP_mult_97_n89) );
  INV_X1 DP_mult_97_U678 ( .A(DP_mult_97_n524), .ZN(DP_mult_97_n73) );
  INV_X1 DP_mult_97_U677 ( .A(DP_mult_97_n552), .ZN(DP_mult_97_n105) );
  OAI21_X1 DP_mult_97_U676 ( .B1(DP_mult_97_n103), .B2(DP_mult_97_n104), .A(
        DP_mult_97_n105), .ZN(DP_mult_97_n469) );
  NAND2_X1 DP_mult_97_U675 ( .A1(DP_mult_97_n283), .A2(DP_mult_97_n286), .ZN(
        DP_mult_97_n154) );
  NAND2_X1 DP_mult_97_U674 ( .A1(DP_mult_97_n281), .A2(DP_mult_97_n282), .ZN(
        DP_mult_97_n145) );
  INV_X1 DP_mult_97_U673 ( .A(DP_mult_97_n591), .ZN(DP_mult_97_n14) );
  OAI21_X1 DP_mult_97_U672 ( .B1(DP_mult_97_n69), .B2(DP_mult_97_n77), .A(
        DP_mult_97_n73), .ZN(DP_mult_97_n443) );
  OAI21_X1 DP_mult_97_U671 ( .B1(DP_mult_97_n87), .B2(DP_mult_97_n88), .A(
        DP_mult_97_n89), .ZN(DP_mult_97_n456) );
  AOI21_X1 DP_mult_97_U670 ( .B1(DP_mult_97_n740), .B2(DP_mult_97_n163), .A(
        DP_mult_97_n139), .ZN(DP_mult_97_n137) );
  NAND2_X1 DP_mult_97_U669 ( .A1(DP_mult_97_n280), .A2(DP_mult_97_n279), .ZN(
        DP_mult_97_n135) );
  OAI21_X1 DP_mult_97_U668 ( .B1(DP_mult_97_n137), .B2(DP_mult_97_n134), .A(
        DP_mult_97_n135), .ZN(DP_mult_97_n133) );
  AOI21_X1 DP_mult_97_U667 ( .B1(DP_mult_97_n168), .B2(DP_mult_97_n132), .A(
        DP_mult_97_n133), .ZN(DP_mult_97_n131) );
  AND2_X1 DP_mult_97_U666 ( .A1(DP_mult_97_n767), .A2(DP_mult_97_n30), .ZN(
        DP_mult_97_n742) );
  NAND2_X1 DP_mult_97_U665 ( .A1(DP_mult_97_n395), .A2(DP_mult_97_n743), .ZN(
        DP_mult_97_n256) );
  INV_X1 DP_mult_97_U664 ( .A(DP_mult_97_n510), .ZN(DP_mult_97_n48) );
  OAI21_X1 DP_mult_97_U663 ( .B1(DP_mult_97_n40), .B2(DP_mult_97_n47), .A(
        DP_mult_97_n48), .ZN(DP_mult_97_n430) );
  INV_X1 DP_mult_97_U662 ( .A(DP_mult_97_n145), .ZN(DP_mult_97_n143) );
  AOI21_X1 DP_mult_97_U661 ( .B1(DP_mult_97_n663), .B2(DP_mult_97_n152), .A(
        DP_mult_97_n143), .ZN(DP_mult_97_n141) );
  INV_X1 DP_mult_97_U660 ( .A(DP_mult_97_n141), .ZN(DP_mult_97_n139) );
  AND2_X1 DP_mult_97_U659 ( .A1(DP_mult_97_n367), .A2(DP_mult_97_n374), .ZN(
        DP_mult_97_n741) );
  OAI21_X1 DP_mult_97_U658 ( .B1(DP_mult_97_n131), .B2(DP_mult_97_n128), .A(
        DP_mult_97_n129), .ZN(DP_mult_97_n127) );
  NOR2_X1 DP_mult_97_U657 ( .A1(DP_mult_97_n130), .A2(DP_mult_97_n128), .ZN(
        DP_mult_97_n126) );
  INV_X1 DP_mult_97_U656 ( .A(DP_mult_97_n154), .ZN(DP_mult_97_n152) );
  NAND2_X1 DP_mult_97_U655 ( .A1(DP_mult_97_n329), .A2(DP_mult_97_n338), .ZN(
        DP_mult_97_n215) );
  NAND2_X1 DP_mult_97_U654 ( .A1(DP_mult_97_n297), .A2(DP_mult_97_n302), .ZN(
        DP_mult_97_n183) );
  NAND2_X1 DP_mult_97_U653 ( .A1(DP_mult_97_n287), .A2(DP_mult_97_n290), .ZN(
        DP_mult_97_n165) );
  NAND2_X1 DP_mult_97_U652 ( .A1(DP_mult_97_n319), .A2(DP_mult_97_n328), .ZN(
        DP_mult_97_n206) );
  NAND2_X1 DP_mult_97_U651 ( .A1(DP_mult_97_n339), .A2(DP_mult_97_n348), .ZN(
        DP_mult_97_n220) );
  NAND2_X1 DP_mult_97_U650 ( .A1(DP_mult_97_n666), .A2(DP_mult_97_n740), .ZN(
        DP_mult_97_n136) );
  INV_X1 DP_mult_97_U649 ( .A(DP_mult_97_n220), .ZN(DP_mult_97_n218) );
  INV_X1 DP_mult_97_U648 ( .A(DP_mult_97_n198), .ZN(DP_mult_97_n273) );
  INV_X1 DP_mult_97_U647 ( .A(DP_mult_97_n668), .ZN(DP_mult_97_n203) );
  AND2_X1 DP_mult_97_U646 ( .A1(DP_mult_97_n665), .A2(DP_mult_97_n663), .ZN(
        DP_mult_97_n740) );
  INV_X1 DP_mult_97_U645 ( .A(DP_mult_97_n214), .ZN(DP_mult_97_n275) );
  INV_X1 DP_mult_97_U644 ( .A(DP_mult_97_n183), .ZN(DP_mult_97_n181) );
  INV_X1 DP_mult_97_U643 ( .A(DP_mult_97_n665), .ZN(DP_mult_97_n149) );
  INV_X1 DP_mult_97_U642 ( .A(DP_mult_97_n165), .ZN(DP_mult_97_n163) );
  INV_X1 DP_mult_97_U641 ( .A(DP_mult_97_n152), .ZN(DP_mult_97_n150) );
  OAI21_X1 DP_mult_97_U640 ( .B1(DP_mult_97_n159), .B2(DP_mult_97_n149), .A(
        DP_mult_97_n150), .ZN(DP_mult_97_n148) );
  AND2_X1 DP_mult_97_U639 ( .A1(DP_mult_97_n668), .A2(DP_mult_97_n206), .ZN(
        DP_mult_97_n739) );
  XNOR2_X1 DP_mult_97_U638 ( .A(DP_mult_97_n207), .B(DP_mult_97_n739), .ZN(
        DP_sw1_a2_3_) );
  NAND2_X1 DP_mult_97_U637 ( .A1(DP_mult_97_n273), .A2(DP_mult_97_n199), .ZN(
        DP_mult_97_n120) );
  NAND2_X1 DP_mult_97_U636 ( .A1(DP_mult_97_n167), .A2(DP_mult_97_n132), .ZN(
        DP_mult_97_n130) );
  NAND2_X1 DP_mult_97_U635 ( .A1(DP_mult_97_n662), .A2(DP_mult_97_n183), .ZN(
        DP_mult_97_n118) );
  INV_X1 DP_mult_97_U634 ( .A(DP_mult_97_n174), .ZN(DP_mult_97_n172) );
  AOI21_X1 DP_mult_97_U633 ( .B1(DP_mult_97_n181), .B2(DP_mult_97_n664), .A(
        DP_mult_97_n172), .ZN(DP_mult_97_n170) );
  OAI21_X1 DP_mult_97_U632 ( .B1(DP_mult_97_n169), .B2(DP_mult_97_n192), .A(
        DP_mult_97_n170), .ZN(DP_mult_97_n168) );
  INV_X1 DP_mult_97_U631 ( .A(DP_mult_97_n192), .ZN(DP_mult_97_n190) );
  INV_X1 DP_mult_97_U630 ( .A(DP_mult_97_n662), .ZN(DP_mult_97_n178) );
  NOR2_X1 DP_mult_97_U629 ( .A1(DP_mult_97_n210), .A2(DP_mult_97_n203), .ZN(
        DP_mult_97_n201) );
  NAND2_X1 DP_mult_97_U628 ( .A1(DP_mult_97_n662), .A2(DP_mult_97_n664), .ZN(
        DP_mult_97_n169) );
  NOR2_X1 DP_mult_97_U627 ( .A1(DP_mult_97_n158), .A2(DP_mult_97_n149), .ZN(
        DP_mult_97_n147) );
  NAND2_X1 DP_mult_97_U626 ( .A1(DP_mult_97_n185), .A2(DP_mult_97_n192), .ZN(
        DP_mult_97_n119) );
  INV_X1 DP_mult_97_U625 ( .A(DP_mult_97_n181), .ZN(DP_mult_97_n179) );
  OAI21_X1 DP_mult_97_U624 ( .B1(DP_mult_97_n192), .B2(DP_mult_97_n178), .A(
        DP_mult_97_n179), .ZN(DP_mult_97_n177) );
  AOI21_X1 DP_mult_97_U623 ( .B1(DP_mult_97_n168), .B2(DP_mult_97_n666), .A(
        DP_mult_97_n163), .ZN(DP_mult_97_n159) );
  INV_X1 DP_mult_97_U622 ( .A(DP_mult_97_n191), .ZN(DP_mult_97_n185) );
  INV_X1 DP_mult_97_U621 ( .A(DP_mult_97_n159), .ZN(DP_mult_97_n157) );
  INV_X1 DP_mult_97_U620 ( .A(DP_mult_97_n210), .ZN(DP_mult_97_n208) );
  NOR2_X1 DP_mult_97_U619 ( .A1(DP_mult_97_n191), .A2(DP_mult_97_n178), .ZN(
        DP_mult_97_n176) );
  NAND2_X1 DP_mult_97_U618 ( .A1(DP_mult_97_n167), .A2(DP_mult_97_n666), .ZN(
        DP_mult_97_n158) );
  INV_X1 DP_mult_97_U617 ( .A(DP_mult_97_n158), .ZN(DP_mult_97_n156) );
  NOR2_X1 DP_mult_97_U616 ( .A1(DP_mult_97_n404), .A2(DP_mult_97_n278), .ZN(
        DP_mult_97_n128) );
  NOR2_X1 DP_mult_97_U615 ( .A1(DP_mult_97_n280), .A2(DP_mult_97_n279), .ZN(
        DP_mult_97_n134) );
  NOR2_X1 DP_mult_97_U614 ( .A1(DP_mult_97_n136), .A2(DP_mult_97_n134), .ZN(
        DP_mult_97_n132) );
  AND2_X1 DP_mult_97_U613 ( .A1(DP_mult_97_n665), .A2(DP_mult_97_n154), .ZN(
        DP_mult_97_n738) );
  XNOR2_X1 DP_mult_97_U612 ( .A(DP_mult_97_n155), .B(DP_mult_97_n738), .ZN(
        DP_sw1_a2_9_) );
  AND2_X1 DP_mult_97_U611 ( .A1(DP_mult_97_n663), .A2(DP_mult_97_n145), .ZN(
        DP_mult_97_n737) );
  XNOR2_X1 DP_mult_97_U610 ( .A(DP_mult_97_n146), .B(DP_mult_97_n737), .ZN(
        DP_sw1_a2_10_) );
  AND2_X1 DP_mult_97_U609 ( .A1(DP_mult_97_n666), .A2(DP_mult_97_n165), .ZN(
        DP_mult_97_n736) );
  XNOR2_X1 DP_mult_97_U608 ( .A(DP_mult_97_n166), .B(DP_mult_97_n736), .ZN(
        DP_sw1_a2_8_) );
  NAND2_X1 DP_mult_97_U607 ( .A1(DP_mult_97_n303), .A2(DP_mult_97_n310), .ZN(
        DP_mult_97_n192) );
  AND2_X1 DP_mult_97_U606 ( .A1(DP_mult_97_n664), .A2(DP_mult_97_n174), .ZN(
        DP_mult_97_n735) );
  XNOR2_X1 DP_mult_97_U605 ( .A(DP_mult_97_n175), .B(DP_mult_97_n735), .ZN(
        DP_sw1_a2_7_) );
  AND2_X1 DP_mult_97_U604 ( .A1(DP_mult_97_n721), .A2(DP_mult_97_n220), .ZN(
        DP_mult_97_n734) );
  XNOR2_X1 DP_mult_97_U603 ( .A(DP_mult_97_n730), .B(DP_mult_97_n734), .ZN(
        DP_sw1_a2_1_) );
  INV_X1 DP_mult_97_U602 ( .A(DP_mult_97_n64), .ZN(DP_mult_97_n733) );
  CLKBUF_X3 DP_mult_97_U601 ( .A(DP_a_int[14]), .Z(DP_mult_97_n732) );
  AND2_X1 DP_mult_97_U600 ( .A1(DP_mult_97_n275), .A2(DP_mult_97_n215), .ZN(
        DP_mult_97_n731) );
  XNOR2_X1 DP_mult_97_U599 ( .A(DP_mult_97_n216), .B(DP_mult_97_n731), .ZN(
        DP_sw1_a2_2_) );
  AOI21_X1 DP_mult_97_U598 ( .B1(DP_mult_97_n688), .B2(DP_mult_97_n716), .A(
        DP_mult_97_n224), .ZN(DP_mult_97_n222) );
  AOI21_X1 DP_mult_97_U597 ( .B1(DP_mult_97_n688), .B2(DP_mult_97_n223), .A(
        DP_mult_97_n224), .ZN(DP_mult_97_n730) );
  XNOR2_X1 DP_mult_97_U596 ( .A(DP_mult_97_n608), .B(DP_sw1_8_), .ZN(
        DP_mult_97_n728) );
  INV_X1 DP_mult_97_U595 ( .A(DP_mult_97_n730), .ZN(DP_mult_97_n726) );
  NAND3_X1 DP_mult_97_U594 ( .A1(DP_mult_97_n723), .A2(DP_mult_97_n724), .A3(
        DP_mult_97_n725), .ZN(DP_mult_97_n358) );
  NAND2_X1 DP_mult_97_U593 ( .A1(DP_mult_97_n363), .A2(DP_mult_97_n368), .ZN(
        DP_mult_97_n725) );
  NAND2_X1 DP_mult_97_U592 ( .A1(DP_mult_97_n361), .A2(DP_mult_97_n368), .ZN(
        DP_mult_97_n724) );
  NAND2_X1 DP_mult_97_U591 ( .A1(DP_mult_97_n361), .A2(DP_mult_97_n363), .ZN(
        DP_mult_97_n723) );
  CLKBUF_X1 DP_mult_97_U590 ( .A(DP_mult_97_n229), .Z(DP_mult_97_n722) );
  OR2_X2 DP_mult_97_U589 ( .A1(DP_mult_97_n339), .A2(DP_mult_97_n348), .ZN(
        DP_mult_97_n721) );
  NAND3_X1 DP_mult_97_U588 ( .A1(DP_mult_97_n718), .A2(DP_mult_97_n719), .A3(
        DP_mult_97_n720), .ZN(DP_mult_97_n338) );
  NAND2_X1 DP_mult_97_U587 ( .A1(DP_mult_97_n350), .A2(DP_mult_97_n343), .ZN(
        DP_mult_97_n720) );
  NAND2_X1 DP_mult_97_U586 ( .A1(DP_mult_97_n341), .A2(DP_mult_97_n343), .ZN(
        DP_mult_97_n719) );
  NAND2_X1 DP_mult_97_U585 ( .A1(DP_mult_97_n341), .A2(DP_mult_97_n350), .ZN(
        DP_mult_97_n718) );
  XOR2_X1 DP_mult_97_U584 ( .A(DP_mult_97_n341), .B(DP_mult_97_n717), .Z(
        DP_mult_97_n339) );
  XOR2_X1 DP_mult_97_U583 ( .A(DP_mult_97_n350), .B(DP_mult_97_n343), .Z(
        DP_mult_97_n717) );
  NOR2_X1 DP_mult_97_U582 ( .A1(DP_mult_97_n228), .A2(DP_mult_97_n225), .ZN(
        DP_mult_97_n716) );
  BUF_X1 DP_mult_97_U581 ( .A(DP_a_int[14]), .Z(DP_mult_97_n604) );
  INV_X1 DP_mult_97_U580 ( .A(DP_sw1_0_), .ZN(DP_mult_97_n713) );
  INV_X1 DP_mult_97_U579 ( .A(DP_mult_97_n604), .ZN(DP_mult_97_n712) );
  NAND2_X1 DP_mult_97_U578 ( .A1(DP_mult_97_n714), .A2(DP_mult_97_n715), .ZN(
        DP_mult_97_n508) );
  NAND2_X1 DP_mult_97_U577 ( .A1(DP_mult_97_n712), .A2(DP_mult_97_n713), .ZN(
        DP_mult_97_n715) );
  NAND2_X1 DP_mult_97_U576 ( .A1(DP_mult_97_n604), .A2(DP_sw1_0_), .ZN(
        DP_mult_97_n714) );
  NAND2_X1 DP_mult_97_U575 ( .A1(DP_mult_97_n694), .A2(DP_mult_97_n582), .ZN(
        DP_mult_97_n612) );
  BUF_X1 DP_mult_97_U574 ( .A(DP_mult_97_n611), .Z(DP_mult_97_n587) );
  NAND3_X1 DP_mult_97_U573 ( .A1(DP_mult_97_n706), .A2(DP_mult_97_n707), .A3(
        DP_mult_97_n708), .ZN(DP_mult_97_n376) );
  NAND2_X1 DP_mult_97_U572 ( .A1(DP_mult_97_n384), .A2(DP_mult_97_n451), .ZN(
        DP_mult_97_n708) );
  NAND2_X1 DP_mult_97_U571 ( .A1(DP_mult_97_n382), .A2(DP_mult_97_n451), .ZN(
        DP_mult_97_n707) );
  NAND2_X1 DP_mult_97_U570 ( .A1(DP_mult_97_n382), .A2(DP_mult_97_n384), .ZN(
        DP_mult_97_n706) );
  XOR2_X1 DP_mult_97_U569 ( .A(DP_mult_97_n382), .B(DP_mult_97_n705), .Z(
        DP_mult_97_n377) );
  XOR2_X1 DP_mult_97_U568 ( .A(DP_mult_97_n384), .B(DP_mult_97_n451), .Z(
        DP_mult_97_n705) );
  NAND3_X1 DP_mult_97_U567 ( .A1(DP_mult_97_n701), .A2(DP_mult_97_n702), .A3(
        DP_mult_97_n703), .ZN(DP_mult_97_n360) );
  NAND2_X1 DP_mult_97_U566 ( .A1(DP_mult_97_n370), .A2(DP_mult_97_n667), .ZN(
        DP_mult_97_n703) );
  NAND2_X1 DP_mult_97_U565 ( .A1(DP_mult_97_n365), .A2(DP_mult_97_n667), .ZN(
        DP_mult_97_n702) );
  NAND2_X1 DP_mult_97_U564 ( .A1(DP_mult_97_n365), .A2(DP_mult_97_n370), .ZN(
        DP_mult_97_n701) );
  INV_X1 DP_mult_97_U563 ( .A(DP_mult_97_n600), .ZN(DP_mult_97_n700) );
  BUF_X1 DP_mult_97_U562 ( .A(DP_mult_97_n726), .Z(DP_mult_97_n768) );
  BUF_X1 DP_mult_97_U561 ( .A(DP_mult_97_n613), .Z(DP_mult_97_n698) );
  BUF_X1 DP_mult_97_U560 ( .A(DP_mult_97_n613), .Z(DP_mult_97_n699) );
  CLKBUF_X2 DP_mult_97_U559 ( .A(DP_a_int[16]), .Z(DP_mult_97_n756) );
  CLKBUF_X1 DP_mult_97_U558 ( .A(DP_mult_97_n349), .Z(DP_mult_97_n697) );
  NOR2_X1 DP_mult_97_U557 ( .A1(DP_mult_97_n391), .A2(DP_mult_97_n394), .ZN(
        DP_mult_97_n696) );
  NOR2_X2 DP_mult_97_U556 ( .A1(DP_mult_97_n329), .A2(DP_mult_97_n338), .ZN(
        DP_mult_97_n214) );
  OR2_X1 DP_mult_97_U555 ( .A1(DP_mult_97_n367), .A2(DP_mult_97_n374), .ZN(
        DP_mult_97_n695) );
  XNOR2_X1 DP_mult_97_U554 ( .A(DP_a_int[20]), .B(DP_a_int[19]), .ZN(
        DP_mult_97_n694) );
  BUF_X1 DP_mult_97_U553 ( .A(DP_mult_97_n612), .Z(DP_mult_97_n710) );
  CLKBUF_X1 DP_mult_97_U552 ( .A(DP_mult_97_n529), .Z(DP_mult_97_n704) );
  INV_X1 DP_mult_97_U551 ( .A(DP_mult_97_n600), .ZN(DP_mult_97_n692) );
  BUF_X1 DP_mult_97_U550 ( .A(DP_mult_97_n616), .Z(DP_mult_97_n729) );
  CLKBUF_X3 DP_mult_97_U549 ( .A(DP_mult_97_n729), .Z(DP_mult_97_n690) );
  OAI21_X1 DP_mult_97_U548 ( .B1(DP_mult_97_n242), .B2(DP_mult_97_n232), .A(
        DP_mult_97_n233), .ZN(DP_mult_97_n688) );
  BUF_X1 DP_mult_97_U547 ( .A(DP_mult_97_n613), .Z(DP_mult_97_n589) );
  BUF_X1 DP_mult_97_U546 ( .A(DP_a_int[20]), .Z(DP_mult_97_n607) );
  CLKBUF_X3 DP_mult_97_U545 ( .A(DP_a_int[20]), .Z(DP_mult_97_n709) );
  BUF_X2 DP_mult_97_U544 ( .A(DP_mult_97_n615), .Z(DP_mult_97_n591) );
  BUF_X2 DP_mult_97_U543 ( .A(DP_mult_97_n610), .Z(DP_mult_97_n691) );
  CLKBUF_X1 DP_mult_97_U542 ( .A(DP_mult_97_n676), .Z(DP_mult_97_n687) );
  NAND3_X1 DP_mult_97_U541 ( .A1(DP_mult_97_n686), .A2(DP_mult_97_n684), .A3(
        DP_mult_97_n685), .ZN(DP_mult_97_n362) );
  NAND2_X1 DP_mult_97_U540 ( .A1(DP_mult_97_n372), .A2(DP_mult_97_n449), .ZN(
        DP_mult_97_n686) );
  NAND2_X1 DP_mult_97_U539 ( .A1(DP_mult_97_n460), .A2(DP_mult_97_n449), .ZN(
        DP_mult_97_n685) );
  NAND2_X1 DP_mult_97_U538 ( .A1(DP_mult_97_n372), .A2(DP_mult_97_n460), .ZN(
        DP_mult_97_n684) );
  XOR2_X1 DP_mult_97_U537 ( .A(DP_mult_97_n683), .B(DP_mult_97_n460), .Z(
        DP_mult_97_n363) );
  XOR2_X1 DP_mult_97_U536 ( .A(DP_mult_97_n372), .B(DP_mult_97_n449), .Z(
        DP_mult_97_n683) );
  CLKBUF_X1 DP_mult_97_U535 ( .A(DP_mult_97_n618), .Z(DP_mult_97_n594) );
  BUF_X2 DP_mult_97_U534 ( .A(DP_mult_97_n618), .Z(DP_mult_97_n682) );
  XNOR2_X1 DP_mult_97_U533 ( .A(DP_mult_97_n363), .B(DP_mult_97_n368), .ZN(
        DP_mult_97_n680) );
  XNOR2_X1 DP_mult_97_U532 ( .A(DP_mult_97_n361), .B(DP_mult_97_n680), .ZN(
        DP_mult_97_n359) );
  XNOR2_X1 DP_mult_97_U531 ( .A(DP_mult_97_n370), .B(DP_mult_97_n667), .ZN(
        DP_mult_97_n679) );
  XNOR2_X1 DP_mult_97_U530 ( .A(DP_mult_97_n365), .B(DP_mult_97_n679), .ZN(
        DP_mult_97_n361) );
  BUF_X1 DP_mult_97_U529 ( .A(DP_mult_97_n610), .Z(DP_mult_97_n755) );
  CLKBUF_X3 DP_mult_97_U528 ( .A(DP_mult_97_n609), .Z(DP_mult_97_n727) );
  BUF_X1 DP_mult_97_U527 ( .A(DP_mult_97_n609), .Z(DP_mult_97_n585) );
  BUF_X2 DP_mult_97_U526 ( .A(DP_a_int[22]), .Z(DP_mult_97_n753) );
  BUF_X1 DP_mult_97_U525 ( .A(DP_mult_97_n617), .Z(DP_mult_97_n754) );
  CLKBUF_X1 DP_mult_97_U524 ( .A(DP_mult_97_n617), .Z(DP_mult_97_n593) );
  BUF_X2 DP_mult_97_U523 ( .A(DP_a_int[18]), .Z(DP_mult_97_n606) );
  CLKBUF_X1 DP_mult_97_U522 ( .A(DP_a_int[16]), .Z(DP_mult_97_n605) );
  CLKBUF_X1 DP_mult_97_U521 ( .A(DP_a_int[22]), .Z(DP_mult_97_n608) );
  BUF_X1 DP_mult_97_U520 ( .A(DP_mult_97_n729), .Z(DP_mult_97_n689) );
  CLKBUF_X1 DP_mult_97_U519 ( .A(DP_mult_97_n762), .Z(DP_mult_97_n677) );
  CLKBUF_X1 DP_mult_97_U518 ( .A(DP_mult_97_n611), .Z(DP_mult_97_n757) );
  BUF_X2 DP_mult_97_U517 ( .A(DP_mult_97_n619), .Z(DP_mult_97_n693) );
  CLKBUF_X1 DP_mult_97_U516 ( .A(DP_mult_97_n619), .Z(DP_mult_97_n595) );
  CLKBUF_X1 DP_mult_97_U515 ( .A(DP_mult_97_n591), .Z(DP_mult_97_n676) );
  BUF_X1 DP_mult_97_U514 ( .A(DP_mult_97_n616), .Z(DP_mult_97_n592) );
  CLKBUF_X3 DP_mult_97_U513 ( .A(DP_mult_97_n614), .Z(DP_mult_97_n762) );
  NAND3_X1 DP_mult_97_U512 ( .A1(DP_mult_97_n673), .A2(DP_mult_97_n674), .A3(
        DP_mult_97_n675), .ZN(DP_mult_97_n380) );
  NAND2_X1 DP_mult_97_U511 ( .A1(DP_mult_97_n388), .A2(DP_mult_97_n385), .ZN(
        DP_mult_97_n675) );
  NAND2_X1 DP_mult_97_U510 ( .A1(DP_mult_97_n383), .A2(DP_mult_97_n385), .ZN(
        DP_mult_97_n674) );
  NAND2_X1 DP_mult_97_U509 ( .A1(DP_mult_97_n383), .A2(DP_mult_97_n388), .ZN(
        DP_mult_97_n673) );
  XOR2_X1 DP_mult_97_U508 ( .A(DP_mult_97_n383), .B(DP_mult_97_n672), .Z(
        DP_mult_97_n381) );
  XOR2_X1 DP_mult_97_U507 ( .A(DP_mult_97_n388), .B(DP_mult_97_n385), .Z(
        DP_mult_97_n672) );
  INV_X1 DP_mult_97_U506 ( .A(DP_mult_97_n597), .ZN(DP_mult_97_n671) );
  CLKBUF_X1 DP_mult_97_U505 ( .A(DP_sw1_7_), .Z(DP_mult_97_n571) );
  BUF_X2 DP_mult_97_U504 ( .A(DP_sw1_7_), .Z(DP_mult_97_n670) );
  OAI22_X1 DP_mult_97_U503 ( .A1(DP_mult_97_n691), .A2(DP_mult_97_n504), .B1(
        DP_mult_97_n690), .B2(DP_mult_97_n503), .ZN(DP_mult_97_n669) );
  OR2_X1 DP_mult_97_U502 ( .A1(DP_mult_97_n319), .A2(DP_mult_97_n328), .ZN(
        DP_mult_97_n668) );
  BUF_X1 DP_mult_97_U501 ( .A(DP_mult_97_n618), .Z(DP_mult_97_n681) );
  BUF_X1 DP_mult_97_U500 ( .A(DP_mult_97_n592), .Z(DP_mult_97_n678) );
  AND2_X1 DP_mult_97_U499 ( .A1(DP_mult_97_n767), .A2(DP_mult_97_n14), .ZN(
        DP_mult_97_n667) );
  OR2_X1 DP_mult_97_U498 ( .A1(DP_mult_97_n287), .A2(DP_mult_97_n290), .ZN(
        DP_mult_97_n666) );
  OR2_X1 DP_mult_97_U497 ( .A1(DP_mult_97_n283), .A2(DP_mult_97_n286), .ZN(
        DP_mult_97_n665) );
  OR2_X1 DP_mult_97_U496 ( .A1(DP_mult_97_n296), .A2(DP_mult_97_n291), .ZN(
        DP_mult_97_n664) );
  OR2_X1 DP_mult_97_U495 ( .A1(DP_mult_97_n281), .A2(DP_mult_97_n282), .ZN(
        DP_mult_97_n663) );
  OR2_X1 DP_mult_97_U494 ( .A1(DP_mult_97_n297), .A2(DP_mult_97_n302), .ZN(
        DP_mult_97_n662) );
  OAI21_X1 DP_mult_97_U493 ( .B1(DP_mult_97_n8), .B2(DP_mult_97_n9), .A(
        DP_mult_97_n10), .ZN(DP_mult_97_n404) );
  NOR2_X1 DP_mult_97_U492 ( .A1(DP_mult_97_n311), .A2(DP_mult_97_n318), .ZN(
        DP_mult_97_n198) );
  INV_X1 DP_mult_97_U491 ( .A(DP_mult_97_n721), .ZN(DP_mult_97_n219) );
  BUF_X2 DP_mult_97_U490 ( .A(DP_mult_97_n612), .Z(DP_mult_97_n711) );
  BUF_X1 DP_mult_97_U489 ( .A(DP_mult_97_n726), .Z(DP_mult_97_n661) );
  OAI21_X2 DP_mult_97_U488 ( .B1(DP_mult_97_n194), .B2(DP_mult_97_n769), .A(
        DP_mult_97_n195), .ZN(DP_mult_97_n193) );
  NOR2_X2 DP_mult_97_U487 ( .A1(DP_mult_97_n303), .A2(DP_mult_97_n310), .ZN(
        DP_mult_97_n191) );
  BUF_X4 DP_mult_97_U464 ( .A(DP_mult_97_n620), .Z(DP_mult_97_n596) );
  HA_X1 DP_mult_97_U274 ( .A(DP_mult_97_n467), .B(DP_mult_97_n479), .CO(
        DP_mult_97_n396), .S(DP_mult_97_n397) );
  FA_X1 DP_mult_97_U273 ( .A(DP_mult_97_n466), .B(DP_mult_97_n478), .CI(
        DP_mult_97_n396), .CO(DP_mult_97_n394), .S(DP_mult_97_n395) );
  HA_X1 DP_mult_97_U272 ( .A(DP_mult_97_n454), .B(DP_mult_97_n477), .CO(
        DP_mult_97_n392), .S(DP_mult_97_n393) );
  FA_X1 DP_mult_97_U271 ( .A(DP_mult_97_n401), .B(DP_mult_97_n465), .CI(
        DP_mult_97_n393), .CO(DP_mult_97_n390), .S(DP_mult_97_n391) );
  FA_X1 DP_mult_97_U270 ( .A(DP_mult_97_n476), .B(DP_mult_97_n464), .CI(
        DP_mult_97_n453), .CO(DP_mult_97_n388), .S(DP_mult_97_n389) );
  FA_X1 DP_mult_97_U269 ( .A(DP_mult_97_n748), .B(DP_mult_97_n392), .CI(
        DP_mult_97_n389), .CO(DP_mult_97_n386), .S(DP_mult_97_n387) );
  HA_X1 DP_mult_97_U268 ( .A(DP_mult_97_n441), .B(DP_mult_97_n452), .CO(
        DP_mult_97_n384), .S(DP_mult_97_n385) );
  FA_X1 DP_mult_97_U267 ( .A(DP_mult_97_n400), .B(DP_mult_97_n463), .CI(
        DP_mult_97_n475), .CO(DP_mult_97_n382), .S(DP_mult_97_n383) );
  FA_X1 DP_mult_97_U265 ( .A(DP_mult_97_n440), .B(DP_mult_97_n474), .CI(
        DP_mult_97_n462), .CO(DP_mult_97_n378), .S(DP_mult_97_n379) );
  HA_X1 DP_mult_97_U262 ( .A(DP_mult_97_n439), .B(DP_mult_97_n428), .CO(
        DP_mult_97_n372), .S(DP_mult_97_n373) );
  FA_X1 DP_mult_97_U261 ( .A(DP_mult_97_n461), .B(DP_mult_97_n450), .CI(
        DP_mult_97_n399), .CO(DP_mult_97_n370), .S(DP_mult_97_n371) );
  FA_X1 DP_mult_97_U260 ( .A(DP_mult_97_n373), .B(DP_mult_97_n473), .CI(
        DP_mult_97_n378), .CO(DP_mult_97_n368), .S(DP_mult_97_n369) );
  FA_X1 DP_mult_97_U259 ( .A(DP_mult_97_n376), .B(DP_mult_97_n371), .CI(
        DP_mult_97_n369), .CO(DP_mult_97_n366), .S(DP_mult_97_n367) );
  FA_X1 DP_mult_97_U258 ( .A(DP_mult_97_n472), .B(DP_mult_97_n427), .CI(
        DP_mult_97_n438), .CO(DP_mult_97_n364), .S(DP_mult_97_n365) );
  HA_X1 DP_mult_97_U254 ( .A(DP_mult_97_n415), .B(DP_mult_97_n426), .CO(
        DP_mult_97_n356), .S(DP_mult_97_n357) );
  FA_X1 DP_mult_97_U253 ( .A(DP_mult_97_n448), .B(DP_mult_97_n471), .CI(
        DP_mult_97_n398), .CO(DP_mult_97_n354), .S(DP_mult_97_n355) );
  FA_X1 DP_mult_97_U252 ( .A(DP_mult_97_n437), .B(DP_mult_97_n459), .CI(
        DP_mult_97_n357), .CO(DP_mult_97_n352), .S(DP_mult_97_n353) );
  FA_X1 DP_mult_97_U251 ( .A(DP_mult_97_n362), .B(DP_mult_97_n364), .CI(
        DP_mult_97_n355), .CO(DP_mult_97_n350), .S(DP_mult_97_n351) );
  FA_X1 DP_mult_97_U250 ( .A(DP_mult_97_n360), .B(DP_mult_97_n353), .CI(
        DP_mult_97_n351), .CO(DP_mult_97_n348), .S(DP_mult_97_n349) );
  HA_X1 DP_mult_97_U249 ( .A(DP_mult_97_n414), .B(DP_mult_97_n425), .CO(
        DP_mult_97_n346), .S(DP_mult_97_n347) );
  FA_X1 DP_mult_97_U248 ( .A(DP_mult_97_n470), .B(DP_mult_97_n447), .CI(
        DP_mult_97_n436), .CO(DP_mult_97_n344), .S(DP_mult_97_n345) );
  FA_X1 DP_mult_97_U247 ( .A(DP_mult_97_n356), .B(DP_mult_97_n458), .CI(
        DP_mult_97_n347), .CO(DP_mult_97_n342), .S(DP_mult_97_n343) );
  FA_X1 DP_mult_97_U246 ( .A(DP_mult_97_n345), .B(DP_mult_97_n354), .CI(
        DP_mult_97_n352), .CO(DP_mult_97_n340), .S(DP_mult_97_n341) );
  FA_X1 DP_mult_97_U242 ( .A(DP_mult_97_n457), .B(DP_mult_97_n446), .CI(
        DP_mult_97_n435), .CO(DP_mult_97_n334), .S(DP_mult_97_n335) );
  FA_X1 DP_mult_97_U241 ( .A(DP_mult_97_n337), .B(DP_mult_97_n346), .CI(
        DP_mult_97_n469), .CO(DP_mult_97_n332), .S(DP_mult_97_n333) );
  FA_X1 DP_mult_97_U240 ( .A(DP_mult_97_n335), .B(DP_mult_97_n344), .CI(
        DP_mult_97_n342), .CO(DP_mult_97_n330), .S(DP_mult_97_n331) );
  FA_X1 DP_mult_97_U239 ( .A(DP_mult_97_n340), .B(DP_mult_97_n333), .CI(
        DP_mult_97_n331), .CO(DP_mult_97_n328), .S(DP_mult_97_n329) );
  FA_X1 DP_mult_97_U237 ( .A(DP_mult_97_n445), .B(DP_mult_97_n423), .CI(
        DP_mult_97_n327), .CO(DP_mult_97_n324), .S(DP_mult_97_n325) );
  FA_X1 DP_mult_97_U236 ( .A(DP_mult_97_n412), .B(DP_mult_97_n434), .CI(
        DP_mult_97_n336), .CO(DP_mult_97_n322), .S(DP_mult_97_n323) );
  FA_X1 DP_mult_97_U235 ( .A(DP_mult_97_n325), .B(DP_mult_97_n334), .CI(
        DP_mult_97_n332), .CO(DP_mult_97_n320), .S(DP_mult_97_n321) );
  FA_X1 DP_mult_97_U234 ( .A(DP_mult_97_n330), .B(DP_mult_97_n323), .CI(
        DP_mult_97_n321), .CO(DP_mult_97_n318), .S(DP_mult_97_n319) );
  FA_X1 DP_mult_97_U233 ( .A(DP_mult_97_n444), .B(DP_mult_97_n411), .CI(
        DP_mult_97_n326), .CO(DP_mult_97_n316), .S(DP_mult_97_n317) );
  FA_X1 DP_mult_97_U232 ( .A(DP_mult_97_n422), .B(DP_mult_97_n433), .CI(
        DP_mult_97_n456), .CO(DP_mult_97_n314), .S(DP_mult_97_n315) );
  FA_X1 DP_mult_97_U231 ( .A(DP_mult_97_n322), .B(DP_mult_97_n324), .CI(
        DP_mult_97_n317), .CO(DP_mult_97_n312), .S(DP_mult_97_n313) );
  FA_X1 DP_mult_97_U230 ( .A(DP_mult_97_n320), .B(DP_mult_97_n315), .CI(
        DP_mult_97_n313), .CO(DP_mult_97_n310), .S(DP_mult_97_n311) );
  FA_X1 DP_mult_97_U228 ( .A(DP_mult_97_n421), .B(DP_mult_97_n410), .CI(
        DP_mult_97_n309), .CO(DP_mult_97_n306), .S(DP_mult_97_n307) );
  FA_X1 DP_mult_97_U227 ( .A(DP_mult_97_n316), .B(DP_mult_97_n432), .CI(
        DP_mult_97_n307), .CO(DP_mult_97_n304), .S(DP_mult_97_n305) );
  FA_X1 DP_mult_97_U226 ( .A(DP_mult_97_n312), .B(DP_mult_97_n314), .CI(
        DP_mult_97_n305), .CO(DP_mult_97_n302), .S(DP_mult_97_n303) );
  FA_X1 DP_mult_97_U225 ( .A(DP_mult_97_n420), .B(DP_mult_97_n409), .CI(
        DP_mult_97_n308), .CO(DP_mult_97_n300), .S(DP_mult_97_n301) );
  FA_X1 DP_mult_97_U224 ( .A(DP_mult_97_n443), .B(DP_mult_97_n431), .CI(
        DP_mult_97_n306), .CO(DP_mult_97_n298), .S(DP_mult_97_n299) );
  FA_X1 DP_mult_97_U223 ( .A(DP_mult_97_n304), .B(DP_mult_97_n301), .CI(
        DP_mult_97_n299), .CO(DP_mult_97_n296), .S(DP_mult_97_n297) );
  FA_X1 DP_mult_97_U221 ( .A(DP_mult_97_n408), .B(DP_mult_97_n419), .CI(
        DP_mult_97_n295), .CO(DP_mult_97_n292), .S(DP_mult_97_n293) );
  FA_X1 DP_mult_97_U220 ( .A(DP_mult_97_n293), .B(DP_mult_97_n300), .CI(
        DP_mult_97_n298), .CO(DP_mult_97_n290), .S(DP_mult_97_n291) );
  FA_X1 DP_mult_97_U219 ( .A(DP_mult_97_n418), .B(DP_mult_97_n294), .CI(
        DP_mult_97_n407), .CO(DP_mult_97_n288), .S(DP_mult_97_n289) );
  FA_X1 DP_mult_97_U218 ( .A(DP_mult_97_n292), .B(DP_mult_97_n430), .CI(
        DP_mult_97_n289), .CO(DP_mult_97_n286), .S(DP_mult_97_n287) );
  FA_X1 DP_mult_97_U216 ( .A(DP_mult_97_n285), .B(DP_mult_97_n406), .CI(
        DP_mult_97_n288), .CO(DP_mult_97_n282), .S(DP_mult_97_n283) );
  FA_X1 DP_mult_97_U215 ( .A(DP_mult_97_n405), .B(DP_mult_97_n284), .CI(
        DP_mult_97_n417), .CO(DP_mult_97_n280), .S(DP_mult_97_n281) );
  OAI21_X1 DP_mult_96_U898 ( .B1(DP_mult_96_n225), .B2(DP_mult_96_n229), .A(
        DP_mult_96_n226), .ZN(DP_mult_96_n224) );
  NOR2_X1 DP_mult_96_U897 ( .A1(DP_mult_96_n228), .A2(DP_mult_96_n225), .ZN(
        DP_mult_96_n223) );
  NAND2_X1 DP_mult_96_U896 ( .A1(DP_mult_96_n391), .A2(DP_mult_96_n394), .ZN(
        DP_mult_96_n254) );
  INV_X1 DP_mult_96_U895 ( .A(DP_a_int[11]), .ZN(DP_mult_96_n620) );
  XOR2_X1 DP_mult_96_U894 ( .A(DP_a_int[11]), .B(DP_a_int[10]), .Z(
        DP_mult_96_n584) );
  NAND2_X1 DP_mult_96_U893 ( .A1(DP_mult_96_n681), .A2(DP_mult_96_n682), .ZN(
        DP_mult_96_n232) );
  AOI21_X1 DP_mult_96_U892 ( .B1(DP_mult_96_n681), .B2(DP_mult_96_n683), .A(
        DP_mult_96_n684), .ZN(DP_mult_96_n233) );
  INV_X1 DP_mult_96_U891 ( .A(DP_mult_96_n231), .ZN(DP_mult_96_n230) );
  OAI21_X1 DP_mult_96_U890 ( .B1(DP_mult_96_n230), .B2(DP_mult_96_n228), .A(
        DP_mult_96_n229), .ZN(DP_mult_96_n227) );
  XNOR2_X1 DP_mult_96_U889 ( .A(DP_mult_96_n605), .B(DP_mult_96_n572), .ZN(
        DP_mult_96_n516) );
  XNOR2_X1 DP_mult_96_U888 ( .A(DP_mult_96_n605), .B(DP_mult_96_n576), .ZN(
        DP_mult_96_n520) );
  XNOR2_X1 DP_mult_96_U887 ( .A(DP_mult_96_n605), .B(DP_mult_96_n573), .ZN(
        DP_mult_96_n517) );
  XNOR2_X1 DP_mult_96_U886 ( .A(DP_mult_96_n605), .B(DP_mult_96_n574), .ZN(
        DP_mult_96_n518) );
  XNOR2_X1 DP_mult_96_U885 ( .A(DP_mult_96_n605), .B(DP_mult_96_n577), .ZN(
        DP_mult_96_n521) );
  NAND2_X1 DP_mult_96_U884 ( .A1(DP_mult_96_n109), .A2(DP_mult_96_n605), .ZN(
        DP_mult_96_n523) );
  XNOR2_X1 DP_mult_96_U883 ( .A(DP_mult_96_n605), .B(DP_mult_96_n571), .ZN(
        DP_mult_96_n515) );
  XNOR2_X1 DP_mult_96_U882 ( .A(DP_mult_96_n605), .B(DP_mult_96_n111), .ZN(
        DP_mult_96_n522) );
  XNOR2_X1 DP_mult_96_U881 ( .A(DP_mult_96_n605), .B(DP_mult_96_n570), .ZN(
        DP_mult_96_n514) );
  XNOR2_X1 DP_mult_96_U880 ( .A(DP_mult_96_n605), .B(DP_mult_96_n569), .ZN(
        DP_mult_96_n513) );
  XNOR2_X1 DP_mult_96_U879 ( .A(DP_mult_96_n605), .B(DP_mult_96_n566), .ZN(
        DP_mult_96_n510) );
  XNOR2_X1 DP_mult_96_U878 ( .A(DP_mult_96_n605), .B(DP_mult_96_n567), .ZN(
        DP_mult_96_n511) );
  XNOR2_X1 DP_mult_96_U877 ( .A(DP_mult_96_n605), .B(DP_mult_96_n568), .ZN(
        DP_mult_96_n512) );
  XNOR2_X1 DP_mult_96_U876 ( .A(DP_mult_96_n227), .B(DP_mult_96_n124), .ZN(
        DP_sw0_a1_0_) );
  INV_X1 DP_mult_96_U875 ( .A(DP_mult_96_n219), .ZN(DP_mult_96_n217) );
  NOR2_X1 DP_mult_96_U874 ( .A1(DP_mult_96_n219), .A2(DP_mult_96_n214), .ZN(
        DP_mult_96_n212) );
  XNOR2_X1 DP_mult_96_U873 ( .A(DP_mult_96_n606), .B(DP_mult_96_n577), .ZN(
        DP_mult_96_n535) );
  XNOR2_X1 DP_mult_96_U872 ( .A(DP_mult_96_n606), .B(DP_mult_96_n111), .ZN(
        DP_mult_96_n536) );
  XNOR2_X1 DP_mult_96_U871 ( .A(DP_mult_96_n606), .B(DP_mult_96_n569), .ZN(
        DP_mult_96_n527) );
  XNOR2_X1 DP_mult_96_U870 ( .A(DP_mult_96_n606), .B(DP_mult_96_n575), .ZN(
        DP_mult_96_n533) );
  XNOR2_X1 DP_mult_96_U869 ( .A(DP_mult_96_n606), .B(DP_mult_96_n576), .ZN(
        DP_mult_96_n534) );
  XNOR2_X1 DP_mult_96_U868 ( .A(DP_mult_96_n606), .B(DP_mult_96_n570), .ZN(
        DP_mult_96_n528) );
  XNOR2_X1 DP_mult_96_U867 ( .A(DP_mult_96_n606), .B(DP_mult_96_n571), .ZN(
        DP_mult_96_n529) );
  XNOR2_X1 DP_mult_96_U866 ( .A(DP_mult_96_n606), .B(DP_mult_96_n572), .ZN(
        DP_mult_96_n530) );
  XNOR2_X1 DP_mult_96_U865 ( .A(DP_mult_96_n606), .B(DP_mult_96_n573), .ZN(
        DP_mult_96_n531) );
  XNOR2_X1 DP_mult_96_U864 ( .A(DP_mult_96_n606), .B(DP_mult_96_n574), .ZN(
        DP_mult_96_n532) );
  XNOR2_X1 DP_mult_96_U863 ( .A(DP_mult_96_n606), .B(DP_mult_96_n566), .ZN(
        DP_mult_96_n524) );
  NAND2_X1 DP_mult_96_U862 ( .A1(DP_mult_96_n109), .A2(DP_mult_96_n606), .ZN(
        DP_mult_96_n537) );
  XNOR2_X1 DP_mult_96_U861 ( .A(DP_mult_96_n606), .B(DP_mult_96_n567), .ZN(
        DP_mult_96_n525) );
  XNOR2_X1 DP_mult_96_U860 ( .A(DP_mult_96_n606), .B(DP_mult_96_n568), .ZN(
        DP_mult_96_n526) );
  OAI21_X1 DP_mult_96_U859 ( .B1(DP_mult_96_n253), .B2(DP_mult_96_n256), .A(
        DP_mult_96_n254), .ZN(DP_mult_96_n252) );
  NOR2_X1 DP_mult_96_U858 ( .A1(DP_mult_96_n253), .A2(DP_mult_96_n255), .ZN(
        DP_mult_96_n251) );
  XOR2_X1 DP_mult_96_U857 ( .A(DP_mult_96_n216), .B(DP_mult_96_n122), .Z(
        DP_sw0_a1_2_) );
  INV_X1 DP_mult_96_U856 ( .A(DP_mult_96_n205), .ZN(DP_mult_96_n204) );
  OAI22_X1 DP_mult_96_U855 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n539), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n538), .ZN(DP_mult_96_n326) );
  INV_X1 DP_mult_96_U854 ( .A(DP_mult_96_n326), .ZN(DP_mult_96_n327) );
  NAND2_X1 DP_mult_96_U853 ( .A1(DP_mult_96_n349), .A2(DP_mult_96_n358), .ZN(
        DP_mult_96_n226) );
  XNOR2_X1 DP_mult_96_U852 ( .A(DP_mult_96_n604), .B(DP_mult_96_n577), .ZN(
        DP_mult_96_n507) );
  XNOR2_X1 DP_mult_96_U851 ( .A(DP_mult_96_n604), .B(DP_mult_96_n574), .ZN(
        DP_mult_96_n504) );
  XNOR2_X1 DP_mult_96_U850 ( .A(DP_mult_96_n604), .B(DP_mult_96_n575), .ZN(
        DP_mult_96_n505) );
  XNOR2_X1 DP_mult_96_U849 ( .A(DP_mult_96_n604), .B(DP_mult_96_n111), .ZN(
        DP_mult_96_n508) );
  XNOR2_X1 DP_mult_96_U848 ( .A(DP_mult_96_n604), .B(DP_mult_96_n576), .ZN(
        DP_mult_96_n506) );
  XNOR2_X1 DP_mult_96_U847 ( .A(DP_mult_96_n604), .B(DP_mult_96_n573), .ZN(
        DP_mult_96_n503) );
  NAND2_X1 DP_mult_96_U846 ( .A1(DP_mult_96_n109), .A2(DP_mult_96_n604), .ZN(
        DP_mult_96_n509) );
  XNOR2_X1 DP_mult_96_U845 ( .A(DP_mult_96_n604), .B(DP_mult_96_n572), .ZN(
        DP_mult_96_n502) );
  XNOR2_X1 DP_mult_96_U844 ( .A(DP_mult_96_n604), .B(DP_mult_96_n570), .ZN(
        DP_mult_96_n500) );
  XNOR2_X1 DP_mult_96_U843 ( .A(DP_mult_96_n604), .B(DP_mult_96_n571), .ZN(
        DP_mult_96_n501) );
  XNOR2_X1 DP_mult_96_U842 ( .A(DP_mult_96_n604), .B(DP_mult_96_n569), .ZN(
        DP_mult_96_n499) );
  XNOR2_X1 DP_mult_96_U841 ( .A(DP_mult_96_n604), .B(DP_mult_96_n568), .ZN(
        DP_mult_96_n498) );
  XNOR2_X1 DP_mult_96_U840 ( .A(DP_mult_96_n604), .B(DP_mult_96_n566), .ZN(
        DP_mult_96_n496) );
  XNOR2_X1 DP_mult_96_U839 ( .A(DP_mult_96_n604), .B(DP_mult_96_n567), .ZN(
        DP_mult_96_n497) );
  XNOR2_X1 DP_mult_96_U838 ( .A(DP_mult_96_n608), .B(DP_mult_96_n576), .ZN(
        DP_mult_96_n562) );
  XNOR2_X1 DP_mult_96_U837 ( .A(DP_mult_96_n608), .B(DP_mult_96_n575), .ZN(
        DP_mult_96_n561) );
  XNOR2_X1 DP_mult_96_U836 ( .A(DP_mult_96_n608), .B(DP_mult_96_n574), .ZN(
        DP_mult_96_n560) );
  XNOR2_X1 DP_mult_96_U835 ( .A(DP_mult_96_n608), .B(DP_mult_96_n573), .ZN(
        DP_mult_96_n559) );
  XNOR2_X1 DP_mult_96_U834 ( .A(DP_mult_96_n608), .B(DP_mult_96_n572), .ZN(
        DP_mult_96_n558) );
  XNOR2_X1 DP_mult_96_U833 ( .A(DP_mult_96_n608), .B(DP_mult_96_n571), .ZN(
        DP_mult_96_n557) );
  XNOR2_X1 DP_mult_96_U832 ( .A(DP_mult_96_n608), .B(DP_mult_96_n570), .ZN(
        DP_mult_96_n556) );
  XNOR2_X1 DP_mult_96_U831 ( .A(DP_mult_96_n608), .B(DP_mult_96_n577), .ZN(
        DP_mult_96_n563) );
  XNOR2_X1 DP_mult_96_U830 ( .A(DP_mult_96_n608), .B(DP_mult_96_n566), .ZN(
        DP_mult_96_n552) );
  XNOR2_X1 DP_mult_96_U829 ( .A(DP_mult_96_n608), .B(DP_mult_96_n567), .ZN(
        DP_mult_96_n553) );
  XNOR2_X1 DP_mult_96_U828 ( .A(DP_mult_96_n608), .B(DP_mult_96_n569), .ZN(
        DP_mult_96_n555) );
  XNOR2_X1 DP_mult_96_U827 ( .A(DP_mult_96_n608), .B(DP_mult_96_n568), .ZN(
        DP_mult_96_n554) );
  XNOR2_X1 DP_mult_96_U826 ( .A(DP_mult_96_n608), .B(DP_mult_96_n111), .ZN(
        DP_mult_96_n564) );
  NAND2_X1 DP_mult_96_U825 ( .A1(DP_mult_96_n109), .A2(DP_mult_96_n608), .ZN(
        DP_mult_96_n565) );
  AOI21_X1 DP_mult_96_U824 ( .B1(DP_mult_96_n231), .B2(DP_mult_96_n223), .A(
        DP_mult_96_n224), .ZN(DP_mult_96_n222) );
  XNOR2_X1 DP_mult_96_U823 ( .A(DP_mult_96_n603), .B(DP_mult_96_n576), .ZN(
        DP_mult_96_n492) );
  XNOR2_X1 DP_mult_96_U822 ( .A(DP_mult_96_n603), .B(DP_mult_96_n577), .ZN(
        DP_mult_96_n493) );
  XNOR2_X1 DP_mult_96_U821 ( .A(DP_mult_96_n603), .B(DP_mult_96_n111), .ZN(
        DP_mult_96_n494) );
  XNOR2_X1 DP_mult_96_U820 ( .A(DP_mult_96_n603), .B(DP_mult_96_n575), .ZN(
        DP_mult_96_n491) );
  NAND2_X1 DP_mult_96_U819 ( .A1(DP_mult_96_n109), .A2(DP_mult_96_n603), .ZN(
        DP_mult_96_n495) );
  XNOR2_X1 DP_mult_96_U818 ( .A(DP_mult_96_n603), .B(DP_mult_96_n573), .ZN(
        DP_mult_96_n489) );
  XNOR2_X1 DP_mult_96_U817 ( .A(DP_mult_96_n603), .B(DP_mult_96_n574), .ZN(
        DP_mult_96_n490) );
  XNOR2_X1 DP_mult_96_U816 ( .A(DP_mult_96_n603), .B(DP_mult_96_n572), .ZN(
        DP_mult_96_n488) );
  XNOR2_X1 DP_mult_96_U815 ( .A(DP_mult_96_n603), .B(DP_mult_96_n571), .ZN(
        DP_mult_96_n487) );
  XNOR2_X1 DP_mult_96_U814 ( .A(DP_mult_96_n603), .B(DP_mult_96_n570), .ZN(
        DP_mult_96_n486) );
  XNOR2_X1 DP_mult_96_U813 ( .A(DP_mult_96_n603), .B(DP_mult_96_n569), .ZN(
        DP_mult_96_n485) );
  XNOR2_X1 DP_mult_96_U812 ( .A(DP_mult_96_n603), .B(DP_mult_96_n567), .ZN(
        DP_mult_96_n483) );
  XNOR2_X1 DP_mult_96_U811 ( .A(DP_mult_96_n603), .B(DP_mult_96_n568), .ZN(
        DP_mult_96_n484) );
  XNOR2_X1 DP_mult_96_U810 ( .A(DP_mult_96_n603), .B(DP_mult_96_n566), .ZN(
        DP_mult_96_n482) );
  XNOR2_X1 DP_mult_96_U809 ( .A(DP_mult_96_n607), .B(DP_mult_96_n111), .ZN(
        DP_mult_96_n550) );
  OAI22_X1 DP_mult_96_U808 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n601), .B1(
        DP_mult_96_n551), .B2(DP_mult_96_n595), .ZN(DP_mult_96_n402) );
  INV_X1 DP_mult_96_U807 ( .A(DP_mult_96_n607), .ZN(DP_mult_96_n601) );
  NAND2_X1 DP_mult_96_U806 ( .A1(DP_mult_96_n395), .A2(DP_mult_96_n667), .ZN(
        DP_mult_96_n256) );
  NOR2_X1 DP_mult_96_U805 ( .A1(DP_mult_96_n395), .A2(DP_mult_96_n667), .ZN(
        DP_mult_96_n255) );
  AOI21_X1 DP_mult_96_U804 ( .B1(DP_mult_96_n251), .B2(DP_mult_96_n257), .A(
        DP_mult_96_n252), .ZN(DP_mult_96_n250) );
  INV_X1 DP_mult_96_U803 ( .A(DP_mult_96_n222), .ZN(DP_mult_96_n221) );
  AOI21_X1 DP_mult_96_U802 ( .B1(DP_mult_96_n221), .B2(DP_mult_96_n217), .A(
        DP_mult_96_n218), .ZN(DP_mult_96_n216) );
  AOI21_X1 DP_mult_96_U801 ( .B1(DP_mult_96_n221), .B2(DP_mult_96_n208), .A(
        DP_mult_96_n209), .ZN(DP_mult_96_n207) );
  AOI21_X1 DP_mult_96_U800 ( .B1(DP_mult_96_n201), .B2(DP_mult_96_n221), .A(
        DP_mult_96_n202), .ZN(DP_mult_96_n200) );
  OAI21_X1 DP_mult_96_U799 ( .B1(DP_mult_96_n194), .B2(DP_mult_96_n676), .A(
        DP_mult_96_n195), .ZN(DP_mult_96_n193) );
  NAND2_X1 DP_mult_96_U798 ( .A1(DP_mult_96_n387), .A2(DP_mult_96_n390), .ZN(
        DP_mult_96_n249) );
  NOR2_X1 DP_mult_96_U797 ( .A1(DP_mult_96_n387), .A2(DP_mult_96_n390), .ZN(
        DP_mult_96_n248) );
  XNOR2_X1 DP_mult_96_U796 ( .A(DP_a_int[7]), .B(DP_a_int[8]), .ZN(
        DP_mult_96_n618) );
  XOR2_X1 DP_mult_96_U795 ( .A(DP_a_int[9]), .B(DP_a_int[8]), .Z(
        DP_mult_96_n583) );
  NAND2_X1 DP_mult_96_U794 ( .A1(DP_mult_96_n581), .A2(DP_mult_96_n617), .ZN(
        DP_mult_96_n611) );
  OAI22_X1 DP_mult_96_U793 ( .A1(DP_mult_96_n674), .A2(DP_mult_96_n599), .B1(
        DP_mult_96_n523), .B2(DP_mult_96_n593), .ZN(DP_mult_96_n400) );
  OAI22_X1 DP_mult_96_U792 ( .A1(DP_mult_96_n587), .A2(DP_mult_96_n520), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n519), .ZN(DP_mult_96_n439) );
  OAI22_X1 DP_mult_96_U791 ( .A1(DP_mult_96_n587), .A2(DP_mult_96_n521), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n675), .ZN(DP_mult_96_n440) );
  OAI22_X1 DP_mult_96_U790 ( .A1(DP_mult_96_n587), .A2(DP_mult_96_n522), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n521), .ZN(DP_mult_96_n441) );
  OAI22_X1 DP_mult_96_U789 ( .A1(DP_mult_96_n674), .A2(DP_mult_96_n519), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n518), .ZN(DP_mult_96_n438) );
  OAI22_X1 DP_mult_96_U788 ( .A1(DP_mult_96_n587), .A2(DP_mult_96_n516), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n515), .ZN(DP_mult_96_n435) );
  OAI22_X1 DP_mult_96_U787 ( .A1(DP_mult_96_n674), .A2(DP_mult_96_n517), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n516), .ZN(DP_mult_96_n436) );
  OAI22_X1 DP_mult_96_U786 ( .A1(DP_mult_96_n674), .A2(DP_mult_96_n518), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n517), .ZN(DP_mult_96_n437) );
  OAI22_X1 DP_mult_96_U785 ( .A1(DP_mult_96_n587), .A2(DP_mult_96_n515), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n514), .ZN(DP_mult_96_n434) );
  OAI22_X1 DP_mult_96_U784 ( .A1(DP_mult_96_n674), .A2(DP_mult_96_n514), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n513), .ZN(DP_mult_96_n433) );
  OAI22_X1 DP_mult_96_U783 ( .A1(DP_mult_96_n587), .A2(DP_mult_96_n511), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n510), .ZN(DP_mult_96_n294) );
  OAI22_X1 DP_mult_96_U782 ( .A1(DP_mult_96_n674), .A2(DP_mult_96_n513), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n512), .ZN(DP_mult_96_n432) );
  OAI22_X1 DP_mult_96_U781 ( .A1(DP_mult_96_n587), .A2(DP_mult_96_n512), .B1(
        DP_mult_96_n593), .B2(DP_mult_96_n511), .ZN(DP_mult_96_n431) );
  NAND2_X1 DP_mult_96_U780 ( .A1(DP_mult_96_n583), .A2(DP_mult_96_n619), .ZN(
        DP_mult_96_n613) );
  OAI22_X1 DP_mult_96_U779 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n545), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n544), .ZN(DP_mult_96_n462) );
  OAI22_X1 DP_mult_96_U778 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n546), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n545), .ZN(DP_mult_96_n463) );
  OAI22_X1 DP_mult_96_U777 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n547), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n546), .ZN(DP_mult_96_n464) );
  OAI22_X1 DP_mult_96_U776 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n550), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n549), .ZN(DP_mult_96_n467) );
  OAI22_X1 DP_mult_96_U775 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n543), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n542), .ZN(DP_mult_96_n460) );
  OAI22_X1 DP_mult_96_U774 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n544), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n543), .ZN(DP_mult_96_n461) );
  OAI22_X1 DP_mult_96_U773 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n548), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n547), .ZN(DP_mult_96_n465) );
  OAI22_X1 DP_mult_96_U772 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n549), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n548), .ZN(DP_mult_96_n466) );
  OAI22_X1 DP_mult_96_U771 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n540), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n539), .ZN(DP_mult_96_n457) );
  OAI22_X1 DP_mult_96_U770 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n541), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n540), .ZN(DP_mult_96_n458) );
  OAI22_X1 DP_mult_96_U769 ( .A1(DP_mult_96_n589), .A2(DP_mult_96_n542), .B1(
        DP_mult_96_n595), .B2(DP_mult_96_n541), .ZN(DP_mult_96_n459) );
  NAND2_X1 DP_mult_96_U768 ( .A1(DP_mult_96_n584), .A2(DP_mult_96_n620), .ZN(
        DP_mult_96_n614) );
  OAI22_X1 DP_mult_96_U767 ( .A1(DP_mult_96_n670), .A2(DP_mult_96_n557), .B1(
        DP_mult_96_n556), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n474) );
  OAI22_X1 DP_mult_96_U766 ( .A1(DP_mult_96_n590), .A2(DP_mult_96_n558), .B1(
        DP_mult_96_n557), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n475) );
  OAI22_X1 DP_mult_96_U765 ( .A1(DP_mult_96_n590), .A2(DP_mult_96_n559), .B1(
        DP_mult_96_n558), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n476) );
  OAI22_X1 DP_mult_96_U764 ( .A1(DP_mult_96_n670), .A2(DP_mult_96_n560), .B1(
        DP_mult_96_n559), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n477) );
  OAI22_X1 DP_mult_96_U763 ( .A1(DP_mult_96_n590), .A2(DP_mult_96_n562), .B1(
        DP_mult_96_n561), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n479) );
  OAI22_X1 DP_mult_96_U762 ( .A1(DP_mult_96_n590), .A2(DP_mult_96_n563), .B1(
        DP_mult_96_n562), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n480) );
  OAI22_X1 DP_mult_96_U761 ( .A1(DP_mult_96_n670), .A2(DP_mult_96_n554), .B1(
        DP_mult_96_n553), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n471) );
  OAI22_X1 DP_mult_96_U760 ( .A1(DP_mult_96_n590), .A2(DP_mult_96_n555), .B1(
        DP_mult_96_n554), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n472) );
  OAI22_X1 DP_mult_96_U759 ( .A1(DP_mult_96_n590), .A2(DP_mult_96_n556), .B1(
        DP_mult_96_n555), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n473) );
  OAI22_X1 DP_mult_96_U758 ( .A1(DP_mult_96_n670), .A2(DP_mult_96_n561), .B1(
        DP_mult_96_n560), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n478) );
  OAI22_X1 DP_mult_96_U757 ( .A1(DP_mult_96_n670), .A2(DP_mult_96_n564), .B1(
        DP_mult_96_n563), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n481) );
  OAI22_X1 DP_mult_96_U756 ( .A1(DP_mult_96_n590), .A2(DP_mult_96_n602), .B1(
        DP_mult_96_n565), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n403) );
  OAI22_X1 DP_mult_96_U755 ( .A1(DP_mult_96_n670), .A2(DP_mult_96_n553), .B1(
        DP_mult_96_n552), .B2(DP_mult_96_n596), .ZN(DP_mult_96_n470) );
  XNOR2_X1 DP_mult_96_U754 ( .A(DP_a_int[3]), .B(DP_a_int[4]), .ZN(
        DP_mult_96_n616) );
  XOR2_X1 DP_mult_96_U753 ( .A(DP_a_int[5]), .B(DP_a_int[4]), .Z(
        DP_mult_96_n581) );
  NAND2_X1 DP_mult_96_U752 ( .A1(DP_mult_96_n580), .A2(DP_mult_96_n616), .ZN(
        DP_mult_96_n610) );
  XNOR2_X1 DP_mult_96_U751 ( .A(DP_mult_96_n113), .B(DP_mult_96_n119), .ZN(
        DP_sw0_a1_5_) );
  INV_X1 DP_mult_96_U750 ( .A(DP_mult_96_n191), .ZN(DP_mult_96_n189) );
  OAI22_X1 DP_mult_96_U749 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n525), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n524), .ZN(DP_mult_96_n308) );
  INV_X1 DP_mult_96_U748 ( .A(DP_mult_96_n308), .ZN(DP_mult_96_n309) );
  NAND2_X1 DP_mult_96_U747 ( .A1(DP_mult_96_n582), .A2(DP_mult_96_n618), .ZN(
        DP_mult_96_n612) );
  XOR2_X1 DP_mult_96_U746 ( .A(DP_a_int[3]), .B(DP_a_int[2]), .Z(
        DP_mult_96_n580) );
  XNOR2_X1 DP_mult_96_U745 ( .A(DP_a_int[1]), .B(DP_a_int[2]), .ZN(
        DP_mult_96_n615) );
  OAI22_X1 DP_mult_96_U744 ( .A1(DP_mult_96_n586), .A2(DP_mult_96_n503), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n502), .ZN(DP_mult_96_n423) );
  OAI22_X1 DP_mult_96_U743 ( .A1(DP_mult_96_n673), .A2(DP_mult_96_n502), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n501), .ZN(DP_mult_96_n422) );
  OAI22_X1 DP_mult_96_U742 ( .A1(DP_mult_96_n586), .A2(DP_mult_96_n501), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n500), .ZN(DP_mult_96_n421) );
  OAI22_X1 DP_mult_96_U741 ( .A1(DP_mult_96_n586), .A2(DP_mult_96_n500), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n499), .ZN(DP_mult_96_n420) );
  OAI22_X1 DP_mult_96_U740 ( .A1(DP_mult_96_n673), .A2(DP_mult_96_n499), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n498), .ZN(DP_mult_96_n419) );
  OAI22_X1 DP_mult_96_U739 ( .A1(DP_mult_96_n586), .A2(DP_mult_96_n497), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n496), .ZN(DP_mult_96_n284) );
  OAI22_X1 DP_mult_96_U738 ( .A1(DP_mult_96_n673), .A2(DP_mult_96_n498), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n497), .ZN(DP_mult_96_n418) );
  XNOR2_X1 DP_mult_96_U737 ( .A(DP_a_int[9]), .B(DP_a_int[10]), .ZN(
        DP_mult_96_n619) );
  OAI21_X1 DP_mult_96_U736 ( .B1(DP_mult_96_n232), .B2(DP_mult_96_n242), .A(
        DP_mult_96_n233), .ZN(DP_mult_96_n231) );
  XNOR2_X1 DP_mult_96_U735 ( .A(DP_mult_96_n607), .B(DP_mult_96_n573), .ZN(
        DP_mult_96_n545) );
  XNOR2_X1 DP_mult_96_U734 ( .A(DP_mult_96_n607), .B(DP_mult_96_n574), .ZN(
        DP_mult_96_n546) );
  BUF_X2 DP_mult_96_U733 ( .A(DP_mult_96_n611), .Z(DP_mult_96_n587) );
  AOI21_X1 DP_mult_96_U732 ( .B1(DP_mult_96_n247), .B2(DP_mult_96_n686), .A(
        DP_mult_96_n685), .ZN(DP_mult_96_n242) );
  INV_X1 DP_mult_96_U731 ( .A(DP_mult_96_n674), .ZN(DP_mult_96_n40) );
  BUF_X2 DP_mult_96_U730 ( .A(DP_sw0_5_), .Z(DP_mult_96_n573) );
  BUF_X2 DP_mult_96_U729 ( .A(DP_sw0_4_), .Z(DP_mult_96_n574) );
  BUF_X2 DP_mult_96_U728 ( .A(DP_sw0_1_), .Z(DP_mult_96_n577) );
  BUF_X2 DP_mult_96_U727 ( .A(DP_sw0_3_), .Z(DP_mult_96_n575) );
  BUF_X2 DP_mult_96_U726 ( .A(DP_sw0_11_), .Z(DP_mult_96_n567) );
  BUF_X2 DP_mult_96_U725 ( .A(DP_sw0_7_), .Z(DP_mult_96_n571) );
  BUF_X2 DP_mult_96_U724 ( .A(DP_sw0_12_), .Z(DP_mult_96_n566) );
  BUF_X2 DP_mult_96_U723 ( .A(DP_sw0_10_), .Z(DP_mult_96_n568) );
  BUF_X2 DP_mult_96_U722 ( .A(DP_sw0_8_), .Z(DP_mult_96_n570) );
  BUF_X2 DP_mult_96_U721 ( .A(DP_sw0_9_), .Z(DP_mult_96_n569) );
  XOR2_X1 DP_mult_96_U720 ( .A(DP_a_int[7]), .B(DP_a_int[6]), .Z(
        DP_mult_96_n582) );
  BUF_X2 DP_mult_96_U719 ( .A(DP_mult_96_n614), .Z(DP_mult_96_n590) );
  BUF_X2 DP_mult_96_U718 ( .A(DP_mult_96_n613), .Z(DP_mult_96_n589) );
  XNOR2_X1 DP_mult_96_U717 ( .A(DP_a_int[5]), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n617) );
  CLKBUF_X3 DP_mult_96_U716 ( .A(DP_a_int[0]), .Z(DP_mult_96_n603) );
  CLKBUF_X3 DP_mult_96_U715 ( .A(DP_a_int[10]), .Z(DP_mult_96_n608) );
  CLKBUF_X3 DP_mult_96_U714 ( .A(DP_a_int[2]), .Z(DP_mult_96_n604) );
  CLKBUF_X3 DP_mult_96_U713 ( .A(DP_a_int[4]), .Z(DP_mult_96_n605) );
  CLKBUF_X3 DP_mult_96_U712 ( .A(DP_a_int[6]), .Z(DP_mult_96_n606) );
  XOR2_X1 DP_mult_96_U711 ( .A(DP_a_int[1]), .B(DP_a_int[0]), .Z(
        DP_mult_96_n579) );
  NAND2_X1 DP_mult_96_U710 ( .A1(DP_mult_96_n579), .A2(DP_mult_96_n615), .ZN(
        DP_mult_96_n609) );
  CLKBUF_X3 DP_mult_96_U709 ( .A(DP_a_int[8]), .Z(DP_mult_96_n607) );
  INV_X1 DP_mult_96_U708 ( .A(DP_mult_96_n588), .ZN(DP_mult_96_n69) );
  OAI22_X1 DP_mult_96_U707 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n486), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n485), .ZN(DP_mult_96_n407) );
  OAI22_X1 DP_mult_96_U706 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n488), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n487), .ZN(DP_mult_96_n409) );
  INV_X1 DP_mult_96_U705 ( .A(DP_mult_96_n284), .ZN(DP_mult_96_n285) );
  OAI22_X1 DP_mult_96_U704 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n485), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n484), .ZN(DP_mult_96_n406) );
  INV_X1 DP_mult_96_U703 ( .A(DP_mult_96_n673), .ZN(DP_mult_96_n24) );
  OAI22_X1 DP_mult_96_U702 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n484), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n483), .ZN(DP_mult_96_n405) );
  OAI21_X1 DP_mult_96_U701 ( .B1(DP_mult_96_n24), .B2(DP_mult_96_n30), .A(
        DP_mult_96_n26), .ZN(DP_mult_96_n417) );
  INV_X1 DP_mult_96_U700 ( .A(DP_mult_96_n585), .ZN(DP_mult_96_n8) );
  INV_X1 DP_mult_96_U699 ( .A(DP_mult_96_n482), .ZN(DP_mult_96_n10) );
  OAI21_X1 DP_mult_96_U698 ( .B1(DP_mult_96_n8), .B2(DP_mult_96_n14), .A(
        DP_mult_96_n10), .ZN(DP_mult_96_n404) );
  INV_X1 DP_mult_96_U697 ( .A(DP_mult_96_n608), .ZN(DP_mult_96_n602) );
  INV_X1 DP_mult_96_U696 ( .A(DP_mult_96_n605), .ZN(DP_mult_96_n599) );
  INV_X1 DP_mult_96_U695 ( .A(DP_mult_96_n603), .ZN(DP_mult_96_n597) );
  INV_X1 DP_mult_96_U694 ( .A(DP_mult_96_n604), .ZN(DP_mult_96_n598) );
  INV_X1 DP_mult_96_U693 ( .A(DP_mult_96_n606), .ZN(DP_mult_96_n600) );
  INV_X1 DP_mult_96_U692 ( .A(DP_mult_96_n670), .ZN(DP_mult_96_n103) );
  INV_X1 DP_mult_96_U691 ( .A(DP_mult_96_n589), .ZN(DP_mult_96_n87) );
  INV_X1 DP_mult_96_U690 ( .A(DP_mult_96_n594), .ZN(DP_mult_96_n77) );
  AND2_X1 DP_mult_96_U689 ( .A1(DP_mult_96_n403), .A2(DP_mult_96_n481), .ZN(
        DP_mult_96_n687) );
  INV_X1 DP_mult_96_U688 ( .A(DP_mult_96_n111), .ZN(DP_mult_96_n109) );
  INV_X1 DP_mult_96_U687 ( .A(DP_mult_96_n595), .ZN(DP_mult_96_n93) );
  OAI22_X1 DP_mult_96_U686 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n494), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n493), .ZN(DP_mult_96_n415) );
  OAI22_X1 DP_mult_96_U685 ( .A1(DP_mult_96_n586), .A2(DP_mult_96_n506), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n505), .ZN(DP_mult_96_n426) );
  OAI22_X1 DP_mult_96_U684 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n527), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n526), .ZN(DP_mult_96_n445) );
  OAI22_X1 DP_mult_96_U683 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n532), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n531), .ZN(DP_mult_96_n450) );
  OAI22_X1 DP_mult_96_U682 ( .A1(DP_mult_96_n673), .A2(DP_mult_96_n598), .B1(
        DP_mult_96_n509), .B2(DP_mult_96_n592), .ZN(DP_mult_96_n399) );
  OAI22_X1 DP_mult_96_U681 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n490), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n489), .ZN(DP_mult_96_n411) );
  OAI22_X1 DP_mult_96_U680 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n526), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n525), .ZN(DP_mult_96_n444) );
  OAI22_X1 DP_mult_96_U679 ( .A1(DP_mult_96_n673), .A2(DP_mult_96_n507), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n506), .ZN(DP_mult_96_n427) );
  INV_X1 DP_mult_96_U678 ( .A(DP_mult_96_n591), .ZN(DP_mult_96_n14) );
  INV_X1 DP_mult_96_U677 ( .A(DP_mult_96_n524), .ZN(DP_mult_96_n73) );
  OAI21_X1 DP_mult_96_U676 ( .B1(DP_mult_96_n69), .B2(DP_mult_96_n77), .A(
        DP_mult_96_n73), .ZN(DP_mult_96_n443) );
  OAI22_X1 DP_mult_96_U675 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n597), .B1(
        DP_mult_96_n495), .B2(DP_mult_96_n591), .ZN(DP_mult_96_n398) );
  OAI22_X1 DP_mult_96_U674 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n530), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n529), .ZN(DP_mult_96_n448) );
  OAI22_X1 DP_mult_96_U673 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n489), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n488), .ZN(DP_mult_96_n410) );
  OR2_X1 DP_mult_96_U672 ( .A1(DP_mult_96_n413), .A2(DP_mult_96_n424), .ZN(
        DP_mult_96_n336) );
  OAI22_X1 DP_mult_96_U671 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n491), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n490), .ZN(DP_mult_96_n412) );
  OAI22_X1 DP_mult_96_U670 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n531), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n530), .ZN(DP_mult_96_n449) );
  OAI22_X1 DP_mult_96_U669 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n535), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n534), .ZN(DP_mult_96_n453) );
  OAI22_X1 DP_mult_96_U668 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n533), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n532), .ZN(DP_mult_96_n451) );
  OAI21_X1 DP_mult_96_U667 ( .B1(DP_mult_96_n87), .B2(DP_mult_96_n93), .A(
        DP_mult_96_n89), .ZN(DP_mult_96_n456) );
  INV_X1 DP_mult_96_U666 ( .A(DP_mult_96_n592), .ZN(DP_mult_96_n30) );
  INV_X1 DP_mult_96_U665 ( .A(DP_mult_96_n294), .ZN(DP_mult_96_n295) );
  OAI22_X1 DP_mult_96_U664 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n487), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n486), .ZN(DP_mult_96_n408) );
  OAI22_X1 DP_mult_96_U663 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n528), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n527), .ZN(DP_mult_96_n446) );
  OAI22_X1 DP_mult_96_U662 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n529), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n528), .ZN(DP_mult_96_n447) );
  OAI22_X1 DP_mult_96_U661 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n600), .B1(
        DP_mult_96_n537), .B2(DP_mult_96_n594), .ZN(DP_mult_96_n401) );
  XNOR2_X1 DP_mult_96_U660 ( .A(DP_mult_96_n607), .B(DP_mult_96_n576), .ZN(
        DP_mult_96_n548) );
  XNOR2_X1 DP_mult_96_U659 ( .A(DP_mult_96_n607), .B(DP_mult_96_n577), .ZN(
        DP_mult_96_n549) );
  XNOR2_X1 DP_mult_96_U658 ( .A(DP_mult_96_n607), .B(DP_mult_96_n575), .ZN(
        DP_mult_96_n547) );
  XNOR2_X1 DP_mult_96_U657 ( .A(DP_mult_96_n607), .B(DP_mult_96_n567), .ZN(
        DP_mult_96_n539) );
  XNOR2_X1 DP_mult_96_U656 ( .A(DP_mult_96_n607), .B(DP_mult_96_n572), .ZN(
        DP_mult_96_n544) );
  XNOR2_X1 DP_mult_96_U655 ( .A(DP_mult_96_n607), .B(DP_mult_96_n568), .ZN(
        DP_mult_96_n540) );
  XNOR2_X1 DP_mult_96_U654 ( .A(DP_mult_96_n607), .B(DP_mult_96_n571), .ZN(
        DP_mult_96_n543) );
  XNOR2_X1 DP_mult_96_U653 ( .A(DP_mult_96_n607), .B(DP_mult_96_n569), .ZN(
        DP_mult_96_n541) );
  XNOR2_X1 DP_mult_96_U652 ( .A(DP_mult_96_n607), .B(DP_mult_96_n570), .ZN(
        DP_mult_96_n542) );
  BUF_X2 DP_mult_96_U651 ( .A(DP_mult_96_n620), .Z(DP_mult_96_n596) );
  CLKBUF_X3 DP_mult_96_U650 ( .A(DP_mult_96_n619), .Z(DP_mult_96_n595) );
  OAI22_X1 DP_mult_96_U649 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n493), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n492), .ZN(DP_mult_96_n414) );
  OAI22_X1 DP_mult_96_U648 ( .A1(DP_mult_96_n586), .A2(DP_mult_96_n505), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n504), .ZN(DP_mult_96_n425) );
  OAI22_X1 DP_mult_96_U647 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n536), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n535), .ZN(DP_mult_96_n454) );
  XNOR2_X1 DP_mult_96_U646 ( .A(DP_mult_96_n607), .B(DP_mult_96_n566), .ZN(
        DP_mult_96_n538) );
  OAI22_X1 DP_mult_96_U645 ( .A1(DP_mult_96_n588), .A2(DP_mult_96_n534), .B1(
        DP_mult_96_n594), .B2(DP_mult_96_n533), .ZN(DP_mult_96_n452) );
  CLKBUF_X3 DP_mult_96_U644 ( .A(DP_mult_96_n616), .Z(DP_mult_96_n592) );
  OAI22_X1 DP_mult_96_U643 ( .A1(DP_mult_96_n586), .A2(DP_mult_96_n508), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n507), .ZN(DP_mult_96_n428) );
  INV_X1 DP_mult_96_U642 ( .A(DP_mult_96_n593), .ZN(DP_mult_96_n57) );
  INV_X1 DP_mult_96_U641 ( .A(DP_mult_96_n510), .ZN(DP_mult_96_n48) );
  OAI21_X1 DP_mult_96_U640 ( .B1(DP_mult_96_n40), .B2(DP_mult_96_n57), .A(
        DP_mult_96_n48), .ZN(DP_mult_96_n430) );
  BUF_X2 DP_mult_96_U639 ( .A(DP_mult_96_n618), .Z(DP_mult_96_n594) );
  CLKBUF_X3 DP_mult_96_U638 ( .A(DP_mult_96_n615), .Z(DP_mult_96_n591) );
  OAI22_X1 DP_mult_96_U637 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n492), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n491), .ZN(DP_mult_96_n413) );
  OAI22_X1 DP_mult_96_U636 ( .A1(DP_mult_96_n673), .A2(DP_mult_96_n504), .B1(
        DP_mult_96_n592), .B2(DP_mult_96_n503), .ZN(DP_mult_96_n424) );
  OR2_X1 DP_mult_96_U635 ( .A1(DP_mult_96_n111), .A2(DP_mult_96_n601), .ZN(
        DP_mult_96_n551) );
  INV_X1 DP_mult_96_U634 ( .A(DP_mult_96_n496), .ZN(DP_mult_96_n26) );
  NAND2_X1 DP_mult_96_U633 ( .A1(DP_mult_96_n280), .A2(DP_mult_96_n279), .ZN(
        DP_mult_96_n135) );
  NAND2_X1 DP_mult_96_U632 ( .A1(DP_mult_96_n281), .A2(DP_mult_96_n282), .ZN(
        DP_mult_96_n145) );
  NAND2_X1 DP_mult_96_U631 ( .A1(DP_mult_96_n287), .A2(DP_mult_96_n290), .ZN(
        DP_mult_96_n165) );
  NAND2_X1 DP_mult_96_U630 ( .A1(DP_mult_96_n283), .A2(DP_mult_96_n286), .ZN(
        DP_mult_96_n154) );
  OAI21_X1 DP_mult_96_U629 ( .B1(DP_mult_96_n137), .B2(DP_mult_96_n134), .A(
        DP_mult_96_n135), .ZN(DP_mult_96_n133) );
  AOI21_X1 DP_mult_96_U628 ( .B1(DP_mult_96_n168), .B2(DP_mult_96_n132), .A(
        DP_mult_96_n133), .ZN(DP_mult_96_n131) );
  NAND2_X1 DP_mult_96_U627 ( .A1(DP_mult_96_n404), .A2(DP_mult_96_n278), .ZN(
        DP_mult_96_n129) );
  OAI21_X1 DP_mult_96_U626 ( .B1(DP_mult_96_n131), .B2(DP_mult_96_n128), .A(
        DP_mult_96_n129), .ZN(DP_mult_96_n127) );
  INV_X1 DP_mult_96_U625 ( .A(DP_mult_96_n278), .ZN(DP_mult_96_n279) );
  NOR2_X1 DP_mult_96_U624 ( .A1(DP_mult_96_n280), .A2(DP_mult_96_n279), .ZN(
        DP_mult_96_n134) );
  NOR2_X1 DP_mult_96_U623 ( .A1(DP_mult_96_n404), .A2(DP_mult_96_n278), .ZN(
        DP_mult_96_n128) );
  OR2_X1 DP_mult_96_U622 ( .A1(DP_mult_96_n381), .A2(DP_mult_96_n386), .ZN(
        DP_mult_96_n686) );
  AND2_X1 DP_mult_96_U621 ( .A1(DP_mult_96_n381), .A2(DP_mult_96_n386), .ZN(
        DP_mult_96_n685) );
  AND2_X1 DP_mult_96_U620 ( .A1(DP_mult_96_n367), .A2(DP_mult_96_n374), .ZN(
        DP_mult_96_n684) );
  AND2_X1 DP_mult_96_U619 ( .A1(DP_mult_96_n375), .A2(DP_mult_96_n377), .ZN(
        DP_mult_96_n683) );
  INV_X1 DP_mult_96_U618 ( .A(DP_mult_96_n538), .ZN(DP_mult_96_n89) );
  OR2_X1 DP_mult_96_U617 ( .A1(DP_mult_96_n375), .A2(DP_mult_96_n377), .ZN(
        DP_mult_96_n682) );
  OR2_X1 DP_mult_96_U616 ( .A1(DP_mult_96_n367), .A2(DP_mult_96_n374), .ZN(
        DP_mult_96_n681) );
  AND2_X1 DP_mult_96_U615 ( .A1(DP_mult_96_n669), .A2(DP_mult_96_n480), .ZN(
        DP_mult_96_n680) );
  OR2_X1 DP_mult_96_U614 ( .A1(DP_mult_96_n669), .A2(DP_mult_96_n480), .ZN(
        DP_mult_96_n679) );
  INV_X1 DP_mult_96_U613 ( .A(DP_mult_96_n552), .ZN(DP_mult_96_n105) );
  AOI21_X1 DP_mult_96_U612 ( .B1(DP_mult_96_n679), .B2(DP_mult_96_n687), .A(
        DP_mult_96_n680), .ZN(DP_mult_96_n260) );
  NOR2_X1 DP_mult_96_U611 ( .A1(DP_mult_96_n397), .A2(DP_mult_96_n402), .ZN(
        DP_mult_96_n258) );
  NAND2_X1 DP_mult_96_U610 ( .A1(DP_mult_96_n397), .A2(DP_mult_96_n402), .ZN(
        DP_mult_96_n259) );
  OAI21_X1 DP_mult_96_U609 ( .B1(DP_mult_96_n260), .B2(DP_mult_96_n258), .A(
        DP_mult_96_n259), .ZN(DP_mult_96_n257) );
  INV_X1 DP_mult_96_U608 ( .A(DP_mult_96_n596), .ZN(DP_mult_96_n104) );
  XNOR2_X1 DP_mult_96_U607 ( .A(DP_mult_96_n413), .B(DP_mult_96_n424), .ZN(
        DP_mult_96_n337) );
  OAI21_X1 DP_mult_96_U606 ( .B1(DP_mult_96_n103), .B2(DP_mult_96_n104), .A(
        DP_mult_96_n105), .ZN(DP_mult_96_n469) );
  XOR2_X1 DP_mult_96_U605 ( .A(DP_mult_96_n207), .B(DP_mult_96_n121), .Z(
        DP_sw0_a1_3_) );
  XOR2_X1 DP_mult_96_U604 ( .A(DP_mult_96_n200), .B(DP_mult_96_n120), .Z(
        DP_sw0_a1_4_) );
  XOR2_X1 DP_mult_96_U603 ( .A(DP_mult_96_n184), .B(DP_mult_96_n118), .Z(
        DP_sw0_a1_6_) );
  XOR2_X1 DP_mult_96_U602 ( .A(DP_mult_96_n166), .B(DP_mult_96_n116), .Z(
        DP_sw0_a1_8_) );
  XOR2_X1 DP_mult_96_U601 ( .A(DP_mult_96_n175), .B(DP_mult_96_n117), .Z(
        DP_sw0_a1_7_) );
  XOR2_X1 DP_mult_96_U600 ( .A(DP_mult_96_n155), .B(DP_mult_96_n115), .Z(
        DP_sw0_a1_9_) );
  XOR2_X1 DP_mult_96_U599 ( .A(DP_mult_96_n146), .B(DP_mult_96_n114), .Z(
        DP_sw0_a1_10_) );
  OAI21_X1 DP_mult_96_U598 ( .B1(DP_mult_96_n250), .B2(DP_mult_96_n248), .A(
        DP_mult_96_n249), .ZN(DP_mult_96_n247) );
  NOR2_X1 DP_mult_96_U597 ( .A1(DP_mult_96_n391), .A2(DP_mult_96_n394), .ZN(
        DP_mult_96_n253) );
  NOR2_X1 DP_mult_96_U596 ( .A1(DP_mult_96_n130), .A2(DP_mult_96_n128), .ZN(
        DP_mult_96_n126) );
  AOI21_X1 DP_mult_96_U595 ( .B1(DP_mult_96_n113), .B2(DP_mult_96_n126), .A(
        DP_mult_96_n127), .ZN(DP_sw0_a1_11_) );
  NAND2_X1 DP_mult_96_U594 ( .A1(DP_mult_96_n664), .A2(DP_mult_96_n154), .ZN(
        DP_mult_96_n115) );
  NAND2_X1 DP_mult_96_U593 ( .A1(DP_mult_96_n662), .A2(DP_mult_96_n145), .ZN(
        DP_mult_96_n114) );
  INV_X1 DP_mult_96_U592 ( .A(DP_mult_96_n165), .ZN(DP_mult_96_n163) );
  INV_X1 DP_mult_96_U591 ( .A(DP_mult_96_n154), .ZN(DP_mult_96_n152) );
  NAND2_X1 DP_mult_96_U590 ( .A1(DP_mult_96_n297), .A2(DP_mult_96_n302), .ZN(
        DP_mult_96_n183) );
  INV_X1 DP_mult_96_U589 ( .A(DP_mult_96_n145), .ZN(DP_mult_96_n143) );
  AOI21_X1 DP_mult_96_U588 ( .B1(DP_mult_96_n662), .B2(DP_mult_96_n152), .A(
        DP_mult_96_n143), .ZN(DP_mult_96_n141) );
  INV_X1 DP_mult_96_U587 ( .A(DP_mult_96_n141), .ZN(DP_mult_96_n139) );
  AOI21_X1 DP_mult_96_U586 ( .B1(DP_mult_96_n678), .B2(DP_mult_96_n163), .A(
        DP_mult_96_n139), .ZN(DP_mult_96_n137) );
  NAND2_X1 DP_mult_96_U585 ( .A1(DP_mult_96_n269), .A2(DP_mult_96_n678), .ZN(
        DP_mult_96_n136) );
  NOR2_X1 DP_mult_96_U584 ( .A1(DP_mult_96_n136), .A2(DP_mult_96_n134), .ZN(
        DP_mult_96_n132) );
  INV_X1 DP_mult_96_U583 ( .A(DP_mult_96_n164), .ZN(DP_mult_96_n269) );
  NAND2_X1 DP_mult_96_U582 ( .A1(DP_mult_96_n269), .A2(DP_mult_96_n165), .ZN(
        DP_mult_96_n116) );
  NAND2_X1 DP_mult_96_U581 ( .A1(DP_mult_96_n359), .A2(DP_mult_96_n366), .ZN(
        DP_mult_96_n229) );
  NAND2_X1 DP_mult_96_U580 ( .A1(DP_mult_96_n329), .A2(DP_mult_96_n338), .ZN(
        DP_mult_96_n215) );
  NOR2_X1 DP_mult_96_U579 ( .A1(DP_mult_96_n359), .A2(DP_mult_96_n366), .ZN(
        DP_mult_96_n228) );
  NAND2_X1 DP_mult_96_U578 ( .A1(DP_mult_96_n296), .A2(DP_mult_96_n291), .ZN(
        DP_mult_96_n174) );
  NAND2_X1 DP_mult_96_U577 ( .A1(DP_mult_96_n311), .A2(DP_mult_96_n318), .ZN(
        DP_mult_96_n199) );
  NAND2_X1 DP_mult_96_U576 ( .A1(DP_mult_96_n319), .A2(DP_mult_96_n328), .ZN(
        DP_mult_96_n206) );
  NOR2_X1 DP_mult_96_U575 ( .A1(DP_mult_96_n339), .A2(DP_mult_96_n348), .ZN(
        DP_mult_96_n219) );
  NOR2_X1 DP_mult_96_U574 ( .A1(DP_mult_96_n319), .A2(DP_mult_96_n328), .ZN(
        DP_mult_96_n205) );
  INV_X1 DP_mult_96_U573 ( .A(DP_mult_96_n152), .ZN(DP_mult_96_n150) );
  NAND2_X1 DP_mult_96_U572 ( .A1(DP_mult_96_n189), .A2(DP_mult_96_n192), .ZN(
        DP_mult_96_n119) );
  AND2_X1 DP_mult_96_U571 ( .A1(DP_mult_96_n664), .A2(DP_mult_96_n662), .ZN(
        DP_mult_96_n678) );
  INV_X1 DP_mult_96_U570 ( .A(DP_mult_96_n183), .ZN(DP_mult_96_n181) );
  NAND2_X1 DP_mult_96_U569 ( .A1(DP_mult_96_n167), .A2(DP_mult_96_n132), .ZN(
        DP_mult_96_n130) );
  INV_X1 DP_mult_96_U568 ( .A(DP_mult_96_n214), .ZN(DP_mult_96_n275) );
  NAND2_X1 DP_mult_96_U567 ( .A1(DP_mult_96_n275), .A2(DP_mult_96_n215), .ZN(
        DP_mult_96_n122) );
  NAND2_X1 DP_mult_96_U566 ( .A1(DP_mult_96_n661), .A2(DP_mult_96_n174), .ZN(
        DP_mult_96_n117) );
  INV_X1 DP_mult_96_U565 ( .A(DP_mult_96_n198), .ZN(DP_mult_96_n273) );
  NAND2_X1 DP_mult_96_U564 ( .A1(DP_mult_96_n273), .A2(DP_mult_96_n199), .ZN(
        DP_mult_96_n120) );
  NAND2_X1 DP_mult_96_U563 ( .A1(DP_mult_96_n663), .A2(DP_mult_96_n183), .ZN(
        DP_mult_96_n118) );
  NAND2_X1 DP_mult_96_U562 ( .A1(DP_mult_96_n204), .A2(DP_mult_96_n206), .ZN(
        DP_mult_96_n121) );
  INV_X1 DP_mult_96_U561 ( .A(DP_mult_96_n225), .ZN(DP_mult_96_n277) );
  INV_X1 DP_mult_96_U560 ( .A(DP_mult_96_n269), .ZN(DP_mult_96_n161) );
  INV_X1 DP_mult_96_U559 ( .A(DP_mult_96_n161), .ZN(DP_mult_96_n160) );
  NAND2_X1 DP_mult_96_U558 ( .A1(DP_mult_96_n277), .A2(DP_mult_96_n226), .ZN(
        DP_mult_96_n124) );
  INV_X1 DP_mult_96_U557 ( .A(DP_mult_96_n204), .ZN(DP_mult_96_n203) );
  OAI21_X1 DP_mult_96_U556 ( .B1(DP_mult_96_n211), .B2(DP_mult_96_n203), .A(
        DP_mult_96_n206), .ZN(DP_mult_96_n202) );
  NOR2_X1 DP_mult_96_U555 ( .A1(DP_mult_96_n210), .A2(DP_mult_96_n203), .ZN(
        DP_mult_96_n201) );
  OAI21_X1 DP_mult_96_U554 ( .B1(DP_mult_96_n198), .B2(DP_mult_96_n206), .A(
        DP_mult_96_n199), .ZN(DP_mult_96_n197) );
  INV_X1 DP_mult_96_U553 ( .A(DP_mult_96_n664), .ZN(DP_mult_96_n149) );
  OAI21_X1 DP_mult_96_U552 ( .B1(DP_mult_96_n159), .B2(DP_mult_96_n149), .A(
        DP_mult_96_n150), .ZN(DP_mult_96_n148) );
  NOR2_X1 DP_mult_96_U551 ( .A1(DP_mult_96_n158), .A2(DP_mult_96_n149), .ZN(
        DP_mult_96_n147) );
  AOI21_X1 DP_mult_96_U550 ( .B1(DP_mult_96_n113), .B2(DP_mult_96_n147), .A(
        DP_mult_96_n148), .ZN(DP_mult_96_n146) );
  AND2_X1 DP_mult_96_U549 ( .A1(DP_mult_96_n217), .A2(DP_mult_96_n220), .ZN(
        DP_mult_96_n677) );
  XOR2_X1 DP_mult_96_U548 ( .A(DP_mult_96_n221), .B(DP_mult_96_n677), .Z(
        DP_sw0_a1_1_) );
  INV_X1 DP_mult_96_U547 ( .A(DP_mult_96_n174), .ZN(DP_mult_96_n172) );
  AOI21_X1 DP_mult_96_U546 ( .B1(DP_mult_96_n181), .B2(DP_mult_96_n661), .A(
        DP_mult_96_n172), .ZN(DP_mult_96_n170) );
  OAI21_X1 DP_mult_96_U545 ( .B1(DP_mult_96_n169), .B2(DP_mult_96_n192), .A(
        DP_mult_96_n170), .ZN(DP_mult_96_n168) );
  INV_X1 DP_mult_96_U544 ( .A(DP_mult_96_n220), .ZN(DP_mult_96_n218) );
  AOI21_X1 DP_mult_96_U543 ( .B1(DP_mult_96_n168), .B2(DP_mult_96_n160), .A(
        DP_mult_96_n163), .ZN(DP_mult_96_n159) );
  NOR2_X1 DP_mult_96_U542 ( .A1(DP_mult_96_n191), .A2(DP_mult_96_n169), .ZN(
        DP_mult_96_n167) );
  NOR2_X1 DP_mult_96_U541 ( .A1(DP_mult_96_n205), .A2(DP_mult_96_n198), .ZN(
        DP_mult_96_n196) );
  OAI21_X1 DP_mult_96_U540 ( .B1(DP_mult_96_n214), .B2(DP_mult_96_n220), .A(
        DP_mult_96_n215), .ZN(DP_mult_96_n213) );
  INV_X1 DP_mult_96_U539 ( .A(DP_mult_96_n181), .ZN(DP_mult_96_n179) );
  INV_X1 DP_mult_96_U538 ( .A(DP_mult_96_n213), .ZN(DP_mult_96_n211) );
  NAND2_X1 DP_mult_96_U537 ( .A1(DP_mult_96_n663), .A2(DP_mult_96_n661), .ZN(
        DP_mult_96_n169) );
  NAND2_X1 DP_mult_96_U536 ( .A1(DP_mult_96_n167), .A2(DP_mult_96_n160), .ZN(
        DP_mult_96_n158) );
  INV_X1 DP_mult_96_U535 ( .A(DP_mult_96_n212), .ZN(DP_mult_96_n210) );
  INV_X1 DP_mult_96_U534 ( .A(DP_mult_96_n192), .ZN(DP_mult_96_n186) );
  INV_X1 DP_mult_96_U533 ( .A(DP_mult_96_n191), .ZN(DP_mult_96_n185) );
  AOI21_X1 DP_mult_96_U532 ( .B1(DP_mult_96_n113), .B2(DP_mult_96_n185), .A(
        DP_mult_96_n186), .ZN(DP_mult_96_n184) );
  INV_X1 DP_mult_96_U531 ( .A(DP_mult_96_n159), .ZN(DP_mult_96_n157) );
  INV_X1 DP_mult_96_U530 ( .A(DP_mult_96_n158), .ZN(DP_mult_96_n156) );
  AOI21_X1 DP_mult_96_U529 ( .B1(DP_mult_96_n113), .B2(DP_mult_96_n156), .A(
        DP_mult_96_n157), .ZN(DP_mult_96_n155) );
  INV_X1 DP_mult_96_U528 ( .A(DP_mult_96_n663), .ZN(DP_mult_96_n178) );
  OAI21_X1 DP_mult_96_U527 ( .B1(DP_mult_96_n192), .B2(DP_mult_96_n178), .A(
        DP_mult_96_n179), .ZN(DP_mult_96_n177) );
  NOR2_X1 DP_mult_96_U526 ( .A1(DP_mult_96_n191), .A2(DP_mult_96_n178), .ZN(
        DP_mult_96_n176) );
  AOI21_X1 DP_mult_96_U525 ( .B1(DP_mult_96_n113), .B2(DP_mult_96_n176), .A(
        DP_mult_96_n177), .ZN(DP_mult_96_n175) );
  AOI21_X1 DP_mult_96_U524 ( .B1(DP_mult_96_n113), .B2(DP_mult_96_n167), .A(
        DP_mult_96_n168), .ZN(DP_mult_96_n166) );
  AOI21_X1 DP_mult_96_U523 ( .B1(DP_mult_96_n196), .B2(DP_mult_96_n213), .A(
        DP_mult_96_n197), .ZN(DP_mult_96_n195) );
  NAND2_X1 DP_mult_96_U522 ( .A1(DP_mult_96_n196), .A2(DP_mult_96_n212), .ZN(
        DP_mult_96_n194) );
  BUF_X2 DP_mult_96_U521 ( .A(DP_mult_96_n193), .Z(DP_mult_96_n113) );
  INV_X1 DP_mult_96_U520 ( .A(DP_mult_96_n211), .ZN(DP_mult_96_n209) );
  INV_X1 DP_mult_96_U519 ( .A(DP_mult_96_n210), .ZN(DP_mult_96_n208) );
  BUF_X2 DP_mult_96_U518 ( .A(DP_mult_96_n612), .Z(DP_mult_96_n588) );
  NOR2_X1 DP_mult_96_U517 ( .A1(DP_mult_96_n287), .A2(DP_mult_96_n290), .ZN(
        DP_mult_96_n164) );
  NAND2_X1 DP_mult_96_U516 ( .A1(DP_mult_96_n303), .A2(DP_mult_96_n310), .ZN(
        DP_mult_96_n192) );
  NAND2_X1 DP_mult_96_U515 ( .A1(DP_mult_96_n339), .A2(DP_mult_96_n348), .ZN(
        DP_mult_96_n220) );
  NOR2_X1 DP_mult_96_U514 ( .A1(DP_mult_96_n329), .A2(DP_mult_96_n338), .ZN(
        DP_mult_96_n214) );
  BUF_X2 DP_mult_96_U513 ( .A(DP_mult_96_n610), .Z(DP_mult_96_n586) );
  XNOR2_X1 DP_mult_96_U512 ( .A(DP_mult_96_n671), .B(DP_sw0_3_), .ZN(
        DP_mult_96_n519) );
  CLKBUF_X1 DP_mult_96_U511 ( .A(DP_mult_96_n222), .Z(DP_mult_96_n676) );
  XNOR2_X1 DP_mult_96_U510 ( .A(DP_mult_96_n605), .B(DP_mult_96_n576), .ZN(
        DP_mult_96_n675) );
  BUF_X2 DP_mult_96_U509 ( .A(DP_mult_96_n611), .Z(DP_mult_96_n674) );
  BUF_X2 DP_mult_96_U508 ( .A(DP_mult_96_n610), .Z(DP_mult_96_n673) );
  XNOR2_X1 DP_mult_96_U507 ( .A(DP_a_int[5]), .B(DP_a_int[6]), .ZN(
        DP_mult_96_n672) );
  CLKBUF_X1 DP_mult_96_U506 ( .A(DP_a_int[4]), .Z(DP_mult_96_n671) );
  BUF_X2 DP_mult_96_U505 ( .A(DP_mult_96_n614), .Z(DP_mult_96_n670) );
  NOR2_X1 DP_mult_96_U504 ( .A1(DP_mult_96_n303), .A2(DP_mult_96_n310), .ZN(
        DP_mult_96_n191) );
  CLKBUF_X3 DP_mult_96_U503 ( .A(DP_mult_96_n672), .Z(DP_mult_96_n593) );
  AND2_X1 DP_mult_96_U502 ( .A1(DP_mult_96_n111), .A2(DP_mult_96_n93), .ZN(
        DP_mult_96_n669) );
  AND2_X1 DP_mult_96_U501 ( .A1(DP_mult_96_n111), .A2(DP_mult_96_n30), .ZN(
        DP_mult_96_n668) );
  AND2_X1 DP_mult_96_U500 ( .A1(DP_mult_96_n111), .A2(DP_mult_96_n77), .ZN(
        DP_mult_96_n667) );
  AND2_X1 DP_mult_96_U499 ( .A1(DP_mult_96_n111), .A2(DP_mult_96_n14), .ZN(
        DP_mult_96_n666) );
  AND2_X1 DP_mult_96_U498 ( .A1(DP_mult_96_n111), .A2(DP_mult_96_n57), .ZN(
        DP_mult_96_n665) );
  BUF_X2 DP_mult_96_U497 ( .A(DP_sw0_0_), .Z(DP_mult_96_n111) );
  OR2_X1 DP_mult_96_U496 ( .A1(DP_mult_96_n283), .A2(DP_mult_96_n286), .ZN(
        DP_mult_96_n664) );
  OR2_X1 DP_mult_96_U495 ( .A1(DP_mult_96_n297), .A2(DP_mult_96_n302), .ZN(
        DP_mult_96_n663) );
  OR2_X1 DP_mult_96_U494 ( .A1(DP_mult_96_n281), .A2(DP_mult_96_n282), .ZN(
        DP_mult_96_n662) );
  OR2_X1 DP_mult_96_U493 ( .A1(DP_mult_96_n296), .A2(DP_mult_96_n291), .ZN(
        DP_mult_96_n661) );
  NOR2_X1 DP_mult_96_U492 ( .A1(DP_mult_96_n311), .A2(DP_mult_96_n318), .ZN(
        DP_mult_96_n198) );
  OAI22_X1 DP_mult_96_U491 ( .A1(DP_mult_96_n585), .A2(DP_mult_96_n483), .B1(
        DP_mult_96_n591), .B2(DP_mult_96_n482), .ZN(DP_mult_96_n278) );
  BUF_X2 DP_mult_96_U490 ( .A(DP_mult_96_n609), .Z(DP_mult_96_n585) );
  NOR2_X2 DP_mult_96_U489 ( .A1(DP_mult_96_n349), .A2(DP_mult_96_n358), .ZN(
        DP_mult_96_n225) );
  CLKBUF_X3 DP_mult_96_U488 ( .A(DP_sw0_6_), .Z(DP_mult_96_n572) );
  CLKBUF_X3 DP_mult_96_U487 ( .A(DP_sw0_2_), .Z(DP_mult_96_n576) );
  HA_X1 DP_mult_96_U274 ( .A(DP_mult_96_n467), .B(DP_mult_96_n479), .CO(
        DP_mult_96_n396), .S(DP_mult_96_n397) );
  FA_X1 DP_mult_96_U273 ( .A(DP_mult_96_n466), .B(DP_mult_96_n478), .CI(
        DP_mult_96_n396), .CO(DP_mult_96_n394), .S(DP_mult_96_n395) );
  HA_X1 DP_mult_96_U272 ( .A(DP_mult_96_n454), .B(DP_mult_96_n477), .CO(
        DP_mult_96_n392), .S(DP_mult_96_n393) );
  FA_X1 DP_mult_96_U271 ( .A(DP_mult_96_n401), .B(DP_mult_96_n465), .CI(
        DP_mult_96_n393), .CO(DP_mult_96_n390), .S(DP_mult_96_n391) );
  FA_X1 DP_mult_96_U270 ( .A(DP_mult_96_n476), .B(DP_mult_96_n464), .CI(
        DP_mult_96_n453), .CO(DP_mult_96_n388), .S(DP_mult_96_n389) );
  FA_X1 DP_mult_96_U269 ( .A(DP_mult_96_n665), .B(DP_mult_96_n392), .CI(
        DP_mult_96_n389), .CO(DP_mult_96_n386), .S(DP_mult_96_n387) );
  HA_X1 DP_mult_96_U268 ( .A(DP_mult_96_n441), .B(DP_mult_96_n452), .CO(
        DP_mult_96_n384), .S(DP_mult_96_n385) );
  FA_X1 DP_mult_96_U267 ( .A(DP_mult_96_n475), .B(DP_mult_96_n400), .CI(
        DP_mult_96_n463), .CO(DP_mult_96_n382), .S(DP_mult_96_n383) );
  FA_X1 DP_mult_96_U266 ( .A(DP_mult_96_n388), .B(DP_mult_96_n385), .CI(
        DP_mult_96_n383), .CO(DP_mult_96_n380), .S(DP_mult_96_n381) );
  FA_X1 DP_mult_96_U265 ( .A(DP_mult_96_n462), .B(DP_mult_96_n474), .CI(
        DP_mult_96_n440), .CO(DP_mult_96_n378), .S(DP_mult_96_n379) );
  FA_X1 DP_mult_96_U264 ( .A(DP_mult_96_n384), .B(DP_mult_96_n451), .CI(
        DP_mult_96_n382), .CO(DP_mult_96_n376), .S(DP_mult_96_n377) );
  FA_X1 DP_mult_96_U263 ( .A(DP_mult_96_n379), .B(DP_mult_96_n668), .CI(
        DP_mult_96_n380), .CO(DP_mult_96_n374), .S(DP_mult_96_n375) );
  HA_X1 DP_mult_96_U262 ( .A(DP_mult_96_n428), .B(DP_mult_96_n439), .CO(
        DP_mult_96_n372), .S(DP_mult_96_n373) );
  FA_X1 DP_mult_96_U261 ( .A(DP_mult_96_n461), .B(DP_mult_96_n450), .CI(
        DP_mult_96_n399), .CO(DP_mult_96_n370), .S(DP_mult_96_n371) );
  FA_X1 DP_mult_96_U260 ( .A(DP_mult_96_n373), .B(DP_mult_96_n473), .CI(
        DP_mult_96_n378), .CO(DP_mult_96_n368), .S(DP_mult_96_n369) );
  FA_X1 DP_mult_96_U259 ( .A(DP_mult_96_n376), .B(DP_mult_96_n371), .CI(
        DP_mult_96_n369), .CO(DP_mult_96_n366), .S(DP_mult_96_n367) );
  FA_X1 DP_mult_96_U258 ( .A(DP_mult_96_n427), .B(DP_mult_96_n472), .CI(
        DP_mult_96_n438), .CO(DP_mult_96_n364), .S(DP_mult_96_n365) );
  FA_X1 DP_mult_96_U257 ( .A(DP_mult_96_n449), .B(DP_mult_96_n460), .CI(
        DP_mult_96_n372), .CO(DP_mult_96_n362), .S(DP_mult_96_n363) );
  FA_X1 DP_mult_96_U256 ( .A(DP_mult_96_n666), .B(DP_mult_96_n370), .CI(
        DP_mult_96_n365), .CO(DP_mult_96_n360), .S(DP_mult_96_n361) );
  FA_X1 DP_mult_96_U255 ( .A(DP_mult_96_n368), .B(DP_mult_96_n363), .CI(
        DP_mult_96_n361), .CO(DP_mult_96_n358), .S(DP_mult_96_n359) );
  HA_X1 DP_mult_96_U254 ( .A(DP_mult_96_n415), .B(DP_mult_96_n426), .CO(
        DP_mult_96_n356), .S(DP_mult_96_n357) );
  FA_X1 DP_mult_96_U253 ( .A(DP_mult_96_n471), .B(DP_mult_96_n448), .CI(
        DP_mult_96_n398), .CO(DP_mult_96_n354), .S(DP_mult_96_n355) );
  FA_X1 DP_mult_96_U252 ( .A(DP_mult_96_n437), .B(DP_mult_96_n459), .CI(
        DP_mult_96_n357), .CO(DP_mult_96_n352), .S(DP_mult_96_n353) );
  FA_X1 DP_mult_96_U251 ( .A(DP_mult_96_n362), .B(DP_mult_96_n364), .CI(
        DP_mult_96_n355), .CO(DP_mult_96_n350), .S(DP_mult_96_n351) );
  FA_X1 DP_mult_96_U250 ( .A(DP_mult_96_n360), .B(DP_mult_96_n353), .CI(
        DP_mult_96_n351), .CO(DP_mult_96_n348), .S(DP_mult_96_n349) );
  HA_X1 DP_mult_96_U249 ( .A(DP_mult_96_n414), .B(DP_mult_96_n425), .CO(
        DP_mult_96_n346), .S(DP_mult_96_n347) );
  FA_X1 DP_mult_96_U248 ( .A(DP_mult_96_n470), .B(DP_mult_96_n447), .CI(
        DP_mult_96_n436), .CO(DP_mult_96_n344), .S(DP_mult_96_n345) );
  FA_X1 DP_mult_96_U247 ( .A(DP_mult_96_n356), .B(DP_mult_96_n458), .CI(
        DP_mult_96_n347), .CO(DP_mult_96_n342), .S(DP_mult_96_n343) );
  FA_X1 DP_mult_96_U246 ( .A(DP_mult_96_n345), .B(DP_mult_96_n354), .CI(
        DP_mult_96_n352), .CO(DP_mult_96_n340), .S(DP_mult_96_n341) );
  FA_X1 DP_mult_96_U245 ( .A(DP_mult_96_n350), .B(DP_mult_96_n343), .CI(
        DP_mult_96_n341), .CO(DP_mult_96_n338), .S(DP_mult_96_n339) );
  FA_X1 DP_mult_96_U242 ( .A(DP_mult_96_n457), .B(DP_mult_96_n446), .CI(
        DP_mult_96_n435), .CO(DP_mult_96_n334), .S(DP_mult_96_n335) );
  FA_X1 DP_mult_96_U241 ( .A(DP_mult_96_n337), .B(DP_mult_96_n346), .CI(
        DP_mult_96_n469), .CO(DP_mult_96_n332), .S(DP_mult_96_n333) );
  FA_X1 DP_mult_96_U240 ( .A(DP_mult_96_n335), .B(DP_mult_96_n344), .CI(
        DP_mult_96_n342), .CO(DP_mult_96_n330), .S(DP_mult_96_n331) );
  FA_X1 DP_mult_96_U239 ( .A(DP_mult_96_n340), .B(DP_mult_96_n333), .CI(
        DP_mult_96_n331), .CO(DP_mult_96_n328), .S(DP_mult_96_n329) );
  FA_X1 DP_mult_96_U237 ( .A(DP_mult_96_n445), .B(DP_mult_96_n423), .CI(
        DP_mult_96_n327), .CO(DP_mult_96_n324), .S(DP_mult_96_n325) );
  FA_X1 DP_mult_96_U236 ( .A(DP_mult_96_n412), .B(DP_mult_96_n434), .CI(
        DP_mult_96_n336), .CO(DP_mult_96_n322), .S(DP_mult_96_n323) );
  FA_X1 DP_mult_96_U235 ( .A(DP_mult_96_n325), .B(DP_mult_96_n334), .CI(
        DP_mult_96_n332), .CO(DP_mult_96_n320), .S(DP_mult_96_n321) );
  FA_X1 DP_mult_96_U234 ( .A(DP_mult_96_n330), .B(DP_mult_96_n323), .CI(
        DP_mult_96_n321), .CO(DP_mult_96_n318), .S(DP_mult_96_n319) );
  FA_X1 DP_mult_96_U233 ( .A(DP_mult_96_n444), .B(DP_mult_96_n411), .CI(
        DP_mult_96_n326), .CO(DP_mult_96_n316), .S(DP_mult_96_n317) );
  FA_X1 DP_mult_96_U232 ( .A(DP_mult_96_n422), .B(DP_mult_96_n433), .CI(
        DP_mult_96_n456), .CO(DP_mult_96_n314), .S(DP_mult_96_n315) );
  FA_X1 DP_mult_96_U231 ( .A(DP_mult_96_n322), .B(DP_mult_96_n324), .CI(
        DP_mult_96_n317), .CO(DP_mult_96_n312), .S(DP_mult_96_n313) );
  FA_X1 DP_mult_96_U230 ( .A(DP_mult_96_n320), .B(DP_mult_96_n315), .CI(
        DP_mult_96_n313), .CO(DP_mult_96_n310), .S(DP_mult_96_n311) );
  FA_X1 DP_mult_96_U228 ( .A(DP_mult_96_n421), .B(DP_mult_96_n410), .CI(
        DP_mult_96_n309), .CO(DP_mult_96_n306), .S(DP_mult_96_n307) );
  FA_X1 DP_mult_96_U227 ( .A(DP_mult_96_n316), .B(DP_mult_96_n432), .CI(
        DP_mult_96_n307), .CO(DP_mult_96_n304), .S(DP_mult_96_n305) );
  FA_X1 DP_mult_96_U226 ( .A(DP_mult_96_n312), .B(DP_mult_96_n314), .CI(
        DP_mult_96_n305), .CO(DP_mult_96_n302), .S(DP_mult_96_n303) );
  FA_X1 DP_mult_96_U225 ( .A(DP_mult_96_n420), .B(DP_mult_96_n409), .CI(
        DP_mult_96_n308), .CO(DP_mult_96_n300), .S(DP_mult_96_n301) );
  FA_X1 DP_mult_96_U224 ( .A(DP_mult_96_n443), .B(DP_mult_96_n431), .CI(
        DP_mult_96_n306), .CO(DP_mult_96_n298), .S(DP_mult_96_n299) );
  FA_X1 DP_mult_96_U223 ( .A(DP_mult_96_n304), .B(DP_mult_96_n301), .CI(
        DP_mult_96_n299), .CO(DP_mult_96_n296), .S(DP_mult_96_n297) );
  FA_X1 DP_mult_96_U221 ( .A(DP_mult_96_n408), .B(DP_mult_96_n419), .CI(
        DP_mult_96_n295), .CO(DP_mult_96_n292), .S(DP_mult_96_n293) );
  FA_X1 DP_mult_96_U220 ( .A(DP_mult_96_n293), .B(DP_mult_96_n300), .CI(
        DP_mult_96_n298), .CO(DP_mult_96_n290), .S(DP_mult_96_n291) );
  FA_X1 DP_mult_96_U219 ( .A(DP_mult_96_n418), .B(DP_mult_96_n294), .CI(
        DP_mult_96_n407), .CO(DP_mult_96_n288), .S(DP_mult_96_n289) );
  FA_X1 DP_mult_96_U218 ( .A(DP_mult_96_n292), .B(DP_mult_96_n430), .CI(
        DP_mult_96_n289), .CO(DP_mult_96_n286), .S(DP_mult_96_n287) );
  FA_X1 DP_mult_96_U216 ( .A(DP_mult_96_n285), .B(DP_mult_96_n406), .CI(
        DP_mult_96_n288), .CO(DP_mult_96_n282), .S(DP_mult_96_n283) );
  FA_X1 DP_mult_96_U215 ( .A(DP_mult_96_n405), .B(DP_mult_96_n284), .CI(
        DP_mult_96_n417), .CO(DP_mult_96_n280), .S(DP_mult_96_n281) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U224 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n145), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n69), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n67) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U223 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n74), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n145), .A(
        DP_sub_1_root_sub_0_root_sub_104_n73), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n71) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U222 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n69), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n73), .A(
        DP_sub_1_root_sub_0_root_sub_104_n70), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n68) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U221 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n93), .A2(DP_x_7_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n42) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U220 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n42), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n83) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U219 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n42), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n50), .A(
        DP_sub_1_root_sub_0_root_sub_104_n43), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n41) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U218 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n49), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n42), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n40) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U217 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n88), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n73), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n11) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U216 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n153), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n74) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U215 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n58), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n64), .A(
        DP_sub_1_root_sub_0_root_sub_104_n59), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n57) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U214 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n148), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n38), .A(
        DP_sub_1_root_sub_0_root_sub_104_n39), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n37) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U213 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n66), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n65) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U212 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n1), .B(
        DP_sub_1_root_sub_0_root_sub_104_n5), .ZN(DP_fb_8_) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U211 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n1), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n33), .A(
        DP_sub_1_root_sub_0_root_sub_104_n34), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n32) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U210 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n1), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n28), .A(
        DP_sub_1_root_sub_0_root_sub_104_n29), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n27) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U209 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n1), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n19), .A(
        DP_sub_1_root_sub_0_root_sub_104_n20), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n18) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U208 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n1), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n14), .A(
        DP_sub_1_root_sub_0_root_sub_104_n15), .ZN(DP_fb_12_) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U207 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n87), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n70), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n10) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U206 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n71), .B(
        DP_sub_1_root_sub_0_root_sub_104_n10), .ZN(DP_fb_3_) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U205 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n65), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n61), .A(
        DP_sub_1_root_sub_0_root_sub_104_n62), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n60) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U204 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n65), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n56), .A(
        DP_sub_1_root_sub_0_root_sub_104_n57), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n51) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U203 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n45), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n65), .A(
        DP_sub_1_root_sub_0_root_sub_104_n46), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n44) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U202 ( .A(DP_sw1_a2_6_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n94) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U201 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n30), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n36), .A(
        DP_sub_1_root_sub_0_root_sub_104_n31), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n29) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U200 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n35), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n30), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n28) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U199 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n157), .B(
        DP_sub_1_root_sub_0_root_sub_104_n78), .ZN(DP_fb_1_) );
  OR2_X1 DP_sub_1_root_sub_0_root_sub_104_U198 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n156), .A2(DP_sw1_a2_1_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n77) );
  XOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U197 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n51), .B(
        DP_sub_1_root_sub_0_root_sub_104_n7), .Z(DP_fb_6_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U196 ( .A(DP_sw1_a2_10_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n90) );
  XOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U195 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n32), .B(
        DP_sub_1_root_sub_0_root_sub_104_n4), .Z(DP_fb_9_) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U194 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n40), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n57), .A(
        DP_sub_1_root_sub_0_root_sub_104_n41), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n39) );
  XOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U193 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n44), .B(
        DP_sub_1_root_sub_0_root_sub_104_n6), .Z(DP_fb_7_) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U192 ( .A(DP_x_1_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n156) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U191 ( .A(DP_x_11_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n101) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U190 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n93), .A2(DP_x_7_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n43) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U189 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n95), .A2(DP_x_5_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n59) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U188 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n91), .A2(DP_x_9_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n31) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U187 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n96), .A2(DP_x_4_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n64) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U186 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n90), .A2(DP_x_10_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n26) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U185 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n92), .A2(DP_x_8_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n36) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U184 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n94), .A2(DP_x_6_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n50) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U183 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n83), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n43), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n6) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U182 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n33), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n36), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n5) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U181 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n58), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n85) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U180 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n30), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n81) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U179 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n81), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n31), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n4) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U178 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n48), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n50), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n7) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U177 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n146), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n26), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n3) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U176 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n54), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n49), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n45) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U175 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n55), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n49), .A(
        DP_sub_1_root_sub_0_root_sub_104_n50), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n46) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U174 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n49), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n48) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U173 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n72), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n88) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U172 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n69), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n87) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U171 ( .A1(DP_sw1_a2_11_), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n101), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n17) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U170 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n64), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n62) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U169 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n63), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n61) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U168 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n36), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n34) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U167 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n35), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n33) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U166 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n26), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n24) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U165 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n22), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n20) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U164 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n56), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n40), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n38) );
  BUF_X2 DP_sub_1_root_sub_0_root_sub_104_U163 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n37), .Z(
        DP_sub_1_root_sub_0_root_sub_104_n1) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U162 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n16), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n79) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U161 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n56), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n54) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U160 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n57), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n55) );
  XOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U159 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n27), .B(
        DP_sub_1_root_sub_0_root_sub_104_n3), .Z(DP_fb_10_) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U158 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n22), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n16), .A(
        DP_sub_1_root_sub_0_root_sub_104_n17), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n15) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U157 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n21), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n16), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n14) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U156 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n21), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n19) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U155 ( .A(DP_sw1_a2_9_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n91) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U154 ( .A(DP_sw1_a2_8_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n92) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U153 ( .A(DP_sw1_a2_7_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n93) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U152 ( .A(DP_sw1_a2_4_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n96) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U151 ( .A(DP_sw1_a2_5_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n95) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U150 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n91), .A2(DP_x_9_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n30) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U149 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n94), .A2(DP_x_6_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n49) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U148 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n95), .A2(DP_x_5_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n58) );
  AOI21_X1 DP_sub_1_root_sub_0_root_sub_104_U147 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n29), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n146), .A(
        DP_sub_1_root_sub_0_root_sub_104_n24), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n22) );
  NAND2_X1 DP_sub_1_root_sub_0_root_sub_104_U146 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n28), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n146), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n21) );
  AND2_X1 DP_sub_1_root_sub_0_root_sub_104_U145 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n79), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n17), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n155) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U144 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n18), .B(
        DP_sub_1_root_sub_0_root_sub_104_n155), .ZN(DP_fb_11_) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U143 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n92), .A2(DP_x_8_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n35) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U142 ( .A1(DP_sw1_a2_11_), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n101), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n16) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U141 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n11), .B(
        DP_sub_1_root_sub_0_root_sub_104_n75), .ZN(DP_fb_2_) );
  BUF_X1 DP_sub_1_root_sub_0_root_sub_104_U140 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n75), .Z(
        DP_sub_1_root_sub_0_root_sub_104_n153) );
  AND2_X1 DP_sub_1_root_sub_0_root_sub_104_U139 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n61), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n64), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n151) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U138 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n66), .B(
        DP_sub_1_root_sub_0_root_sub_104_n151), .ZN(DP_fb_4_) );
  AND2_X1 DP_sub_1_root_sub_0_root_sub_104_U137 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n85), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n59), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n150) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U136 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n60), .B(
        DP_sub_1_root_sub_0_root_sub_104_n150), .ZN(DP_fb_5_) );
  AND2_X1 DP_sub_1_root_sub_0_root_sub_104_U135 ( .A1(DP_sw1_a2_0_), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n149), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n78) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U134 ( .A(DP_sw1_a2_1_), .B(
        DP_x_1_), .ZN(DP_sub_1_root_sub_0_root_sub_104_n157) );
  OAI21_X1 DP_sub_1_root_sub_0_root_sub_104_U133 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n147), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n78), .A(
        DP_sub_1_root_sub_0_root_sub_104_n77), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n75) );
  OR2_X1 DP_sub_1_root_sub_0_root_sub_104_U132 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n152), .A2(DP_sw1_a2_3_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n70) );
  OR2_X1 DP_sub_1_root_sub_0_root_sub_104_U131 ( .A1(DP_sw1_a2_2_), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n154), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n73) );
  XNOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U130 ( .A(DP_sw1_a2_0_), .B(
        DP_sub_1_root_sub_0_root_sub_104_n149), .ZN(DP_fb_0_) );
  AND2_X2 DP_sub_1_root_sub_0_root_sub_104_U129 ( .A1(DP_sw1_a2_3_), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n152), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n69) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U128 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n63), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n58), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n56) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U127 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n65), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n148) );
  NOR2_X1 DP_sub_1_root_sub_0_root_sub_104_U126 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n96), .A2(DP_x_4_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n63) );
  AND2_X1 DP_sub_1_root_sub_0_root_sub_104_U125 ( .A1(DP_sw1_a2_1_), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n156), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n147) );
  OR2_X1 DP_sub_1_root_sub_0_root_sub_104_U124 ( .A1(
        DP_sub_1_root_sub_0_root_sub_104_n90), .A2(DP_x_10_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n146) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U123 ( .A(DP_x_2_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n154) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U122 ( .A(DP_x_3_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n152) );
  INV_X1 DP_sub_1_root_sub_0_root_sub_104_U121 ( .A(DP_x_0_), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n149) );
  AOI21_X2 DP_sub_1_root_sub_0_root_sub_104_U120 ( .B1(
        DP_sub_1_root_sub_0_root_sub_104_n67), .B2(
        DP_sub_1_root_sub_0_root_sub_104_n153), .A(
        DP_sub_1_root_sub_0_root_sub_104_n68), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n66) );
  AND2_X1 DP_sub_1_root_sub_0_root_sub_104_U119 ( .A1(DP_sw1_a2_2_), .A2(
        DP_sub_1_root_sub_0_root_sub_104_n154), .ZN(
        DP_sub_1_root_sub_0_root_sub_104_n72) );
  BUF_X1 DP_sub_1_root_sub_0_root_sub_104_U118 ( .A(
        DP_sub_1_root_sub_0_root_sub_104_n72), .Z(
        DP_sub_1_root_sub_0_root_sub_104_n145) );
  XNOR2_X1 DP_mult_105_U982 ( .A(DP_w_11_), .B(DP_mult_105_n608), .ZN(
        DP_mult_105_n553) );
  XNOR2_X1 DP_mult_105_U981 ( .A(DP_w_11_), .B(DP_mult_105_n607), .ZN(
        DP_mult_105_n539) );
  XNOR2_X1 DP_mult_105_U980 ( .A(DP_mult_105_n712), .B(DP_mult_105_n606), .ZN(
        DP_mult_105_n525) );
  XNOR2_X1 DP_mult_105_U979 ( .A(DP_mult_105_n605), .B(DP_mult_105_n712), .ZN(
        DP_mult_105_n511) );
  NAND2_X1 DP_mult_105_U978 ( .A1(DP_mult_105_n349), .A2(DP_mult_105_n358), 
        .ZN(DP_mult_105_n226) );
  OAI21_X1 DP_mult_105_U977 ( .B1(DP_mult_105_n225), .B2(DP_mult_105_n229), 
        .A(DP_mult_105_n226), .ZN(DP_mult_105_n224) );
  XNOR2_X1 DP_mult_105_U976 ( .A(DP_mult_105_n604), .B(DP_mult_105_n712), .ZN(
        DP_mult_105_n497) );
  NOR2_X1 DP_mult_105_U975 ( .A1(DP_mult_105_n228), .A2(DP_mult_105_n225), 
        .ZN(DP_mult_105_n223) );
  XNOR2_X1 DP_mult_105_U974 ( .A(DP_mult_105_n603), .B(DP_mult_105_n712), .ZN(
        DP_mult_105_n483) );
  NOR2_X1 DP_mult_105_U973 ( .A1(DP_mult_105_n203), .A2(DP_mult_105_n198), 
        .ZN(DP_mult_105_n196) );
  OAI21_X1 DP_mult_105_U972 ( .B1(DP_mult_105_n198), .B2(DP_mult_105_n206), 
        .A(DP_mult_105_n199), .ZN(DP_mult_105_n197) );
  AOI21_X1 DP_mult_105_U971 ( .B1(DP_mult_105_n196), .B2(DP_mult_105_n209), 
        .A(DP_mult_105_n197), .ZN(DP_mult_105_n195) );
  NAND2_X1 DP_mult_105_U970 ( .A1(DP_mult_105_n185), .A2(DP_mult_105_n192), 
        .ZN(DP_mult_105_n119) );
  XNOR2_X1 DP_mult_105_U969 ( .A(DP_mult_105_n193), .B(DP_mult_105_n119), .ZN(
        DP_w_b0_5_) );
  XNOR2_X1 DP_mult_105_U968 ( .A(DP_w_12_), .B(DP_mult_105_n606), .ZN(
        DP_mult_105_n524) );
  INV_X1 DP_mult_105_U967 ( .A(DP_mult_105_n308), .ZN(DP_mult_105_n309) );
  XNOR2_X1 DP_mult_105_U966 ( .A(DP_w_12_), .B(DP_mult_105_n608), .ZN(
        DP_mult_105_n552) );
  AOI21_X1 DP_mult_105_U965 ( .B1(DP_mult_105_n223), .B2(DP_mult_105_n231), 
        .A(DP_mult_105_n224), .ZN(DP_mult_105_n222) );
  OAI21_X1 DP_mult_105_U964 ( .B1(DP_mult_105_n194), .B2(DP_mult_105_n763), 
        .A(DP_mult_105_n195), .ZN(DP_mult_105_n193) );
  INV_X1 DP_mult_105_U963 ( .A(DP_mult_105_n552), .ZN(DP_mult_105_n105) );
  NOR2_X1 DP_mult_105_U962 ( .A1(DP_mult_105_n339), .A2(DP_mult_105_n348), 
        .ZN(DP_mult_105_n219) );
  OAI22_X1 DP_mult_105_U961 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n731), 
        .B1(DP_mult_105_n553), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n471) );
  XNOR2_X1 DP_mult_105_U960 ( .A(DP_mult_105_n221), .B(DP_mult_105_n123), .ZN(
        DP_w_b0_1_) );
  NAND2_X1 DP_mult_105_U959 ( .A1(DP_mult_105_n319), .A2(DP_mult_105_n328), 
        .ZN(DP_mult_105_n206) );
  INV_X1 DP_mult_105_U958 ( .A(DP_mult_105_n211), .ZN(DP_mult_105_n209) );
  AOI21_X1 DP_mult_105_U957 ( .B1(DP_mult_105_n747), .B2(DP_mult_105_n208), 
        .A(DP_mult_105_n213), .ZN(DP_mult_105_n207) );
  NAND2_X1 DP_mult_105_U956 ( .A1(DP_mult_105_n732), .A2(DP_mult_105_n220), 
        .ZN(DP_mult_105_n123) );
  INV_X1 DP_mult_105_U955 ( .A(DP_mult_105_n222), .ZN(DP_mult_105_n221) );
  INV_X1 DP_mult_105_U954 ( .A(DP_mult_105_n220), .ZN(DP_mult_105_n218) );
  AOI21_X1 DP_mult_105_U953 ( .B1(DP_mult_105_n689), .B2(DP_mult_105_n727), 
        .A(DP_mult_105_n218), .ZN(DP_mult_105_n216) );
  OAI22_X1 DP_mult_105_U952 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n557), 
        .B1(DP_mult_105_n556), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n474) );
  OAI22_X1 DP_mult_105_U951 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n556), 
        .B1(DP_mult_105_n555), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n473) );
  OAI21_X1 DP_mult_105_U950 ( .B1(DP_mult_105_n214), .B2(DP_mult_105_n220), 
        .A(DP_mult_105_n215), .ZN(DP_mult_105_n213) );
  AOI21_X1 DP_mult_105_U949 ( .B1(DP_mult_105_n201), .B2(DP_mult_105_n747), 
        .A(DP_mult_105_n202), .ZN(DP_mult_105_n200) );
  NOR2_X1 DP_mult_105_U948 ( .A1(DP_mult_105_n329), .A2(DP_mult_105_n338), 
        .ZN(DP_mult_105_n214) );
  NAND2_X1 DP_mult_105_U947 ( .A1(DP_mult_105_n339), .A2(DP_mult_105_n348), 
        .ZN(DP_mult_105_n220) );
  XNOR2_X1 DP_mult_105_U946 ( .A(DP_mult_105_n566), .B(DP_mult_105_n607), .ZN(
        DP_mult_105_n538) );
  XNOR2_X1 DP_mult_105_U945 ( .A(DP_mult_105_n605), .B(DP_mult_105_n566), .ZN(
        DP_mult_105_n510) );
  XNOR2_X1 DP_mult_105_U944 ( .A(DP_mult_105_n604), .B(DP_mult_105_n566), .ZN(
        DP_mult_105_n496) );
  XNOR2_X1 DP_mult_105_U943 ( .A(DP_mult_105_n603), .B(DP_mult_105_n566), .ZN(
        DP_mult_105_n482) );
  INV_X1 DP_mult_105_U942 ( .A(DP_mult_105_n689), .ZN(DP_mult_105_n763) );
  CLKBUF_X1 DP_mult_105_U941 ( .A(DP_mult_105_n717), .Z(DP_mult_105_n762) );
  OAI21_X1 DP_mult_105_U940 ( .B1(DP_mult_105_n230), .B2(DP_mult_105_n228), 
        .A(DP_mult_105_n229), .ZN(DP_mult_105_n227) );
  XNOR2_X1 DP_mult_105_U939 ( .A(DP_w_10_), .B(DP_mult_105_n608), .ZN(
        DP_mult_105_n554) );
  NAND2_X1 DP_mult_105_U938 ( .A1(DP_mult_105_n329), .A2(DP_mult_105_n338), 
        .ZN(DP_mult_105_n215) );
  NAND3_X1 DP_mult_105_U937 ( .A1(DP_mult_105_n759), .A2(DP_mult_105_n760), 
        .A3(DP_mult_105_n761), .ZN(DP_mult_105_n338) );
  NAND2_X1 DP_mult_105_U936 ( .A1(DP_mult_105_n350), .A2(DP_mult_105_n343), 
        .ZN(DP_mult_105_n761) );
  NAND2_X1 DP_mult_105_U935 ( .A1(DP_mult_105_n739), .A2(DP_mult_105_n343), 
        .ZN(DP_mult_105_n760) );
  NAND2_X1 DP_mult_105_U934 ( .A1(DP_mult_105_n739), .A2(DP_mult_105_n350), 
        .ZN(DP_mult_105_n759) );
  NAND3_X1 DP_mult_105_U933 ( .A1(DP_mult_105_n756), .A2(DP_mult_105_n757), 
        .A3(DP_mult_105_n758), .ZN(DP_mult_105_n350) );
  NAND2_X1 DP_mult_105_U932 ( .A1(DP_mult_105_n688), .A2(DP_mult_105_n729), 
        .ZN(DP_mult_105_n758) );
  NAND2_X1 DP_mult_105_U931 ( .A1(DP_mult_105_n362), .A2(DP_mult_105_n729), 
        .ZN(DP_mult_105_n757) );
  NAND2_X1 DP_mult_105_U930 ( .A1(DP_mult_105_n688), .A2(DP_mult_105_n362), 
        .ZN(DP_mult_105_n756) );
  NAND3_X1 DP_mult_105_U929 ( .A1(DP_mult_105_n753), .A2(DP_mult_105_n754), 
        .A3(DP_mult_105_n755), .ZN(DP_mult_105_n354) );
  NAND2_X1 DP_mult_105_U928 ( .A1(DP_mult_105_n448), .A2(DP_mult_105_n728), 
        .ZN(DP_mult_105_n755) );
  NAND2_X1 DP_mult_105_U927 ( .A1(DP_mult_105_n398), .A2(DP_mult_105_n728), 
        .ZN(DP_mult_105_n754) );
  NAND2_X1 DP_mult_105_U926 ( .A1(DP_mult_105_n398), .A2(DP_mult_105_n448), 
        .ZN(DP_mult_105_n753) );
  OAI22_X1 DP_mult_105_U925 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n539), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n538), .ZN(DP_mult_105_n326) );
  INV_X1 DP_mult_105_U924 ( .A(DP_mult_105_n326), .ZN(DP_mult_105_n327) );
  NAND3_X1 DP_mult_105_U923 ( .A1(DP_mult_105_n750), .A2(DP_mult_105_n751), 
        .A3(DP_mult_105_n752), .ZN(DP_mult_105_n340) );
  NAND2_X1 DP_mult_105_U922 ( .A1(DP_mult_105_n354), .A2(DP_mult_105_n352), 
        .ZN(DP_mult_105_n752) );
  NAND2_X1 DP_mult_105_U921 ( .A1(DP_mult_105_n345), .A2(DP_mult_105_n352), 
        .ZN(DP_mult_105_n751) );
  NAND2_X1 DP_mult_105_U920 ( .A1(DP_mult_105_n345), .A2(DP_mult_105_n354), 
        .ZN(DP_mult_105_n750) );
  NOR2_X1 DP_mult_105_U919 ( .A1(DP_mult_105_n359), .A2(DP_mult_105_n366), 
        .ZN(DP_mult_105_n228) );
  INV_X1 DP_mult_105_U918 ( .A(DP_mult_105_n231), .ZN(DP_mult_105_n230) );
  XNOR2_X1 DP_mult_105_U917 ( .A(DP_mult_105_n364), .B(DP_mult_105_n362), .ZN(
        DP_mult_105_n749) );
  XNOR2_X1 DP_mult_105_U916 ( .A(DP_mult_105_n355), .B(DP_mult_105_n749), .ZN(
        DP_mult_105_n351) );
  OAI22_X1 DP_mult_105_U915 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n539), 
        .B1(DP_mult_105_n538), .B2(DP_mult_105_n595), .ZN(DP_mult_105_n748) );
  OAI22_X1 DP_mult_105_U914 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n540), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n539), .ZN(DP_mult_105_n457) );
  INV_X1 DP_mult_105_U913 ( .A(DP_mult_105_n763), .ZN(DP_mult_105_n747) );
  XOR2_X1 DP_mult_105_U912 ( .A(DP_mult_105_n607), .B(DP_mult_105_n566), .Z(
        DP_mult_105_n746) );
  OAI21_X1 DP_mult_105_U911 ( .B1(DP_mult_105_n211), .B2(DP_mult_105_n203), 
        .A(DP_mult_105_n206), .ZN(DP_mult_105_n202) );
  NOR2_X1 DP_mult_105_U910 ( .A1(DP_mult_105_n721), .A2(DP_mult_105_n203), 
        .ZN(DP_mult_105_n201) );
  NAND2_X1 DP_mult_105_U909 ( .A1(DP_mult_105_n196), .A2(DP_mult_105_n212), 
        .ZN(DP_mult_105_n194) );
  XNOR2_X1 DP_mult_105_U908 ( .A(DP_mult_105_n398), .B(DP_mult_105_n448), .ZN(
        DP_mult_105_n745) );
  XNOR2_X1 DP_mult_105_U907 ( .A(DP_mult_105_n471), .B(DP_mult_105_n745), .ZN(
        DP_mult_105_n355) );
  NAND2_X1 DP_mult_105_U906 ( .A1(DP_mult_105_n359), .A2(DP_mult_105_n366), 
        .ZN(DP_mult_105_n229) );
  AOI21_X1 DP_mult_105_U905 ( .B1(DP_mult_105_n704), .B2(DP_mult_105_n673), 
        .A(DP_mult_105_n705), .ZN(DP_mult_105_n233) );
  NAND2_X1 DP_mult_105_U904 ( .A1(DP_mult_105_n704), .A2(DP_mult_105_n709), 
        .ZN(DP_mult_105_n232) );
  XNOR2_X1 DP_mult_105_U903 ( .A(DP_mult_105_n608), .B(DP_mult_105_n570), .ZN(
        DP_mult_105_n556) );
  XNOR2_X1 DP_mult_105_U902 ( .A(DP_mult_105_n354), .B(DP_mult_105_n352), .ZN(
        DP_mult_105_n744) );
  XNOR2_X1 DP_mult_105_U901 ( .A(DP_mult_105_n345), .B(DP_mult_105_n744), .ZN(
        DP_mult_105_n341) );
  NOR2_X1 DP_mult_105_U900 ( .A1(DP_mult_105_n349), .A2(DP_mult_105_n358), 
        .ZN(DP_mult_105_n225) );
  NAND3_X1 DP_mult_105_U899 ( .A1(DP_mult_105_n741), .A2(DP_mult_105_n742), 
        .A3(DP_mult_105_n743), .ZN(DP_mult_105_n358) );
  NAND2_X1 DP_mult_105_U898 ( .A1(DP_mult_105_n368), .A2(DP_mult_105_n363), 
        .ZN(DP_mult_105_n743) );
  NAND2_X1 DP_mult_105_U897 ( .A1(DP_mult_105_n361), .A2(DP_mult_105_n363), 
        .ZN(DP_mult_105_n742) );
  NAND2_X1 DP_mult_105_U896 ( .A1(DP_mult_105_n361), .A2(DP_mult_105_n368), 
        .ZN(DP_mult_105_n741) );
  OAI22_X1 DP_mult_105_U895 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n525), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n524), .ZN(DP_mult_105_n308) );
  INV_X1 DP_mult_105_U894 ( .A(DP_mult_105_n213), .ZN(DP_mult_105_n211) );
  XNOR2_X1 DP_mult_105_U893 ( .A(DP_mult_105_n607), .B(DP_mult_105_n711), .ZN(
        DP_mult_105_n540) );
  XNOR2_X1 DP_mult_105_U892 ( .A(DP_mult_105_n606), .B(DP_mult_105_n711), .ZN(
        DP_mult_105_n526) );
  XNOR2_X1 DP_mult_105_U891 ( .A(DP_mult_105_n605), .B(DP_mult_105_n711), .ZN(
        DP_mult_105_n512) );
  XNOR2_X1 DP_mult_105_U890 ( .A(DP_mult_105_n604), .B(DP_mult_105_n722), .ZN(
        DP_mult_105_n498) );
  XNOR2_X1 DP_mult_105_U889 ( .A(DP_mult_105_n603), .B(DP_mult_105_n722), .ZN(
        DP_mult_105_n484) );
  XOR2_X1 DP_mult_105_U888 ( .A(DP_mult_105_n155), .B(DP_mult_105_n115), .Z(
        DP_w_b0_9_) );
  OR2_X1 DP_mult_105_U887 ( .A1(DP_mult_105_n358), .A2(DP_mult_105_n349), .ZN(
        DP_mult_105_n740) );
  XNOR2_X1 DP_mult_105_U886 ( .A(DP_mult_105_n608), .B(DP_w_9_), .ZN(
        DP_mult_105_n555) );
  OAI22_X1 DP_mult_105_U885 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n511), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n510), .ZN(DP_mult_105_n294) );
  INV_X1 DP_mult_105_U884 ( .A(DP_mult_105_n294), .ZN(DP_mult_105_n295) );
  XNOR2_X1 DP_mult_105_U883 ( .A(DP_mult_105_n345), .B(DP_mult_105_n744), .ZN(
        DP_mult_105_n739) );
  NAND3_X1 DP_mult_105_U882 ( .A1(DP_mult_105_n736), .A2(DP_mult_105_n737), 
        .A3(DP_mult_105_n738), .ZN(DP_mult_105_n320) );
  NAND2_X1 DP_mult_105_U881 ( .A1(DP_mult_105_n332), .A2(DP_mult_105_n325), 
        .ZN(DP_mult_105_n738) );
  NAND2_X1 DP_mult_105_U880 ( .A1(DP_mult_105_n334), .A2(DP_mult_105_n325), 
        .ZN(DP_mult_105_n737) );
  NAND2_X1 DP_mult_105_U879 ( .A1(DP_mult_105_n334), .A2(DP_mult_105_n332), 
        .ZN(DP_mult_105_n736) );
  NAND3_X1 DP_mult_105_U878 ( .A1(DP_mult_105_n733), .A2(DP_mult_105_n734), 
        .A3(DP_mult_105_n735), .ZN(DP_mult_105_n324) );
  NAND2_X1 DP_mult_105_U877 ( .A1(DP_mult_105_n423), .A2(DP_mult_105_n327), 
        .ZN(DP_mult_105_n735) );
  NAND2_X1 DP_mult_105_U876 ( .A1(DP_mult_105_n445), .A2(DP_mult_105_n327), 
        .ZN(DP_mult_105_n734) );
  NAND2_X1 DP_mult_105_U875 ( .A1(DP_mult_105_n445), .A2(DP_mult_105_n423), 
        .ZN(DP_mult_105_n733) );
  OR2_X1 DP_mult_105_U874 ( .A1(DP_mult_105_n339), .A2(DP_mult_105_n348), .ZN(
        DP_mult_105_n732) );
  CLKBUF_X1 DP_mult_105_U873 ( .A(DP_mult_105_n554), .Z(DP_mult_105_n731) );
  NAND2_X1 DP_mult_105_U872 ( .A1(DP_mult_105_n311), .A2(DP_mult_105_n318), 
        .ZN(DP_mult_105_n199) );
  AOI21_X1 DP_mult_105_U871 ( .B1(DP_mult_105_n698), .B2(DP_mult_105_n185), 
        .A(DP_mult_105_n190), .ZN(DP_mult_105_n184) );
  AOI21_X1 DP_mult_105_U870 ( .B1(DP_mult_105_n697), .B2(DP_mult_105_n176), 
        .A(DP_mult_105_n177), .ZN(DP_mult_105_n175) );
  AOI21_X1 DP_mult_105_U869 ( .B1(DP_mult_105_n698), .B2(DP_mult_105_n167), 
        .A(DP_mult_105_n168), .ZN(DP_mult_105_n166) );
  AOI21_X1 DP_mult_105_U868 ( .B1(DP_mult_105_n697), .B2(DP_mult_105_n156), 
        .A(DP_mult_105_n157), .ZN(DP_mult_105_n155) );
  AOI21_X1 DP_mult_105_U867 ( .B1(DP_mult_105_n698), .B2(DP_mult_105_n147), 
        .A(DP_mult_105_n148), .ZN(DP_mult_105_n146) );
  AOI21_X1 DP_mult_105_U866 ( .B1(DP_mult_105_n697), .B2(DP_mult_105_n126), 
        .A(DP_mult_105_n127), .ZN(DP_w_b0_11_) );
  AOI21_X1 DP_mult_105_U865 ( .B1(DP_mult_105_n247), .B2(DP_mult_105_n674), 
        .A(DP_mult_105_n669), .ZN(DP_mult_105_n242) );
  NAND2_X1 DP_mult_105_U864 ( .A1(DP_mult_105_n730), .A2(DP_mult_105_n233), 
        .ZN(DP_mult_105_n231) );
  OR2_X1 DP_mult_105_U863 ( .A1(DP_mult_105_n232), .A2(DP_mult_105_n242), .ZN(
        DP_mult_105_n730) );
  OAI22_X1 DP_mult_105_U862 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n731), 
        .B1(DP_mult_105_n717), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n728) );
  INV_X1 DP_mult_105_U861 ( .A(DP_mult_105_n219), .ZN(DP_mult_105_n727) );
  OAI22_X1 DP_mult_105_U860 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n529), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n528), .ZN(DP_mult_105_n447) );
  OAI22_X1 DP_mult_105_U859 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n517), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n516), .ZN(DP_mult_105_n436) );
  OR2_X1 DP_mult_105_U858 ( .A1(DP_mult_105_n338), .A2(DP_mult_105_n329), .ZN(
        DP_mult_105_n726) );
  NAND3_X1 DP_mult_105_U857 ( .A1(DP_mult_105_n724), .A2(DP_mult_105_n723), 
        .A3(DP_mult_105_n725), .ZN(DP_mult_105_n344) );
  NAND2_X1 DP_mult_105_U856 ( .A1(DP_mult_105_n447), .A2(DP_mult_105_n436), 
        .ZN(DP_mult_105_n725) );
  NAND2_X1 DP_mult_105_U855 ( .A1(DP_mult_105_n718), .A2(DP_mult_105_n436), 
        .ZN(DP_mult_105_n724) );
  NAND2_X1 DP_mult_105_U854 ( .A1(DP_mult_105_n718), .A2(DP_mult_105_n447), 
        .ZN(DP_mult_105_n723) );
  CLKBUF_X1 DP_mult_105_U853 ( .A(DP_mult_105_n711), .Z(DP_mult_105_n722) );
  XNOR2_X1 DP_mult_105_U852 ( .A(DP_mult_105_n607), .B(DP_w_9_), .ZN(
        DP_mult_105_n541) );
  XNOR2_X1 DP_mult_105_U851 ( .A(DP_mult_105_n606), .B(DP_w_9_), .ZN(
        DP_mult_105_n527) );
  XNOR2_X1 DP_mult_105_U850 ( .A(DP_mult_105_n604), .B(DP_mult_105_n569), .ZN(
        DP_mult_105_n499) );
  XNOR2_X1 DP_mult_105_U849 ( .A(DP_mult_105_n605), .B(DP_w_9_), .ZN(
        DP_mult_105_n513) );
  XNOR2_X1 DP_mult_105_U848 ( .A(DP_mult_105_n603), .B(DP_mult_105_n569), .ZN(
        DP_mult_105_n485) );
  XNOR2_X1 DP_mult_105_U847 ( .A(DP_mult_105_n607), .B(DP_mult_105_n570), .ZN(
        DP_mult_105_n542) );
  XNOR2_X1 DP_mult_105_U846 ( .A(DP_mult_105_n606), .B(DP_mult_105_n570), .ZN(
        DP_mult_105_n528) );
  XNOR2_X1 DP_mult_105_U845 ( .A(DP_mult_105_n604), .B(DP_mult_105_n570), .ZN(
        DP_mult_105_n500) );
  XNOR2_X1 DP_mult_105_U844 ( .A(DP_mult_105_n605), .B(DP_mult_105_n570), .ZN(
        DP_mult_105_n514) );
  XNOR2_X1 DP_mult_105_U843 ( .A(DP_mult_105_n603), .B(DP_mult_105_n570), .ZN(
        DP_mult_105_n486) );
  XNOR2_X1 DP_mult_105_U842 ( .A(DP_mult_105_n447), .B(DP_mult_105_n436), .ZN(
        DP_mult_105_n720) );
  XNOR2_X1 DP_mult_105_U841 ( .A(DP_mult_105_n719), .B(DP_mult_105_n720), .ZN(
        DP_mult_105_n345) );
  OAI22_X1 DP_mult_105_U840 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n762), 
        .B1(DP_mult_105_n552), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n718) );
  OAI22_X1 DP_mult_105_U839 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n762), 
        .B1(DP_mult_105_n552), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n719) );
  XNOR2_X1 DP_mult_105_U838 ( .A(DP_w_11_), .B(DP_mult_105_n608), .ZN(
        DP_mult_105_n717) );
  NAND3_X1 DP_mult_105_U837 ( .A1(DP_mult_105_n714), .A2(DP_mult_105_n715), 
        .A3(DP_mult_105_n716), .ZN(DP_mult_105_n366) );
  NAND2_X1 DP_mult_105_U836 ( .A1(DP_mult_105_n376), .A2(DP_mult_105_n371), 
        .ZN(DP_mult_105_n716) );
  NAND2_X1 DP_mult_105_U835 ( .A1(DP_mult_105_n369), .A2(DP_mult_105_n371), 
        .ZN(DP_mult_105_n715) );
  NAND2_X1 DP_mult_105_U834 ( .A1(DP_mult_105_n369), .A2(DP_mult_105_n376), 
        .ZN(DP_mult_105_n714) );
  XNOR2_X1 DP_mult_105_U833 ( .A(DP_mult_105_n334), .B(DP_mult_105_n332), .ZN(
        DP_mult_105_n713) );
  XNOR2_X1 DP_mult_105_U832 ( .A(DP_mult_105_n713), .B(DP_mult_105_n325), .ZN(
        DP_mult_105_n321) );
  CLKBUF_X1 DP_mult_105_U831 ( .A(DP_w_11_), .Z(DP_mult_105_n712) );
  CLKBUF_X1 DP_mult_105_U830 ( .A(DP_w_10_), .Z(DP_mult_105_n711) );
  XNOR2_X1 DP_mult_105_U829 ( .A(DP_mult_105_n445), .B(DP_mult_105_n423), .ZN(
        DP_mult_105_n710) );
  XOR2_X1 DP_mult_105_U828 ( .A(DP_mult_105_n184), .B(DP_mult_105_n118), .Z(
        DP_w_b0_6_) );
  INV_X1 DP_mult_105_U827 ( .A(DP_b_int[11]), .ZN(DP_mult_105_n620) );
  XOR2_X1 DP_mult_105_U826 ( .A(DP_b_int[7]), .B(DP_b_int[6]), .Z(
        DP_mult_105_n582) );
  NAND2_X1 DP_mult_105_U825 ( .A1(DP_mult_105_n582), .A2(DP_mult_105_n618), 
        .ZN(DP_mult_105_n612) );
  BUF_X1 DP_mult_105_U824 ( .A(DP_mult_105_n612), .Z(DP_mult_105_n588) );
  XOR2_X1 DP_mult_105_U823 ( .A(DP_b_int[5]), .B(DP_b_int[4]), .Z(
        DP_mult_105_n581) );
  NAND2_X1 DP_mult_105_U822 ( .A1(DP_mult_105_n581), .A2(DP_mult_105_n617), 
        .ZN(DP_mult_105_n611) );
  BUF_X1 DP_mult_105_U821 ( .A(DP_mult_105_n611), .Z(DP_mult_105_n587) );
  XOR2_X1 DP_mult_105_U820 ( .A(DP_b_int[9]), .B(DP_b_int[8]), .Z(
        DP_mult_105_n583) );
  NAND2_X1 DP_mult_105_U819 ( .A1(DP_mult_105_n583), .A2(DP_mult_105_n619), 
        .ZN(DP_mult_105_n613) );
  BUF_X1 DP_mult_105_U818 ( .A(DP_mult_105_n613), .Z(DP_mult_105_n589) );
  XOR2_X1 DP_mult_105_U817 ( .A(DP_b_int[3]), .B(DP_b_int[2]), .Z(
        DP_mult_105_n580) );
  NAND2_X1 DP_mult_105_U816 ( .A1(DP_mult_105_n580), .A2(DP_mult_105_n616), 
        .ZN(DP_mult_105_n610) );
  BUF_X1 DP_mult_105_U815 ( .A(DP_mult_105_n610), .Z(DP_mult_105_n586) );
  XOR2_X1 DP_mult_105_U814 ( .A(DP_b_int[1]), .B(DP_b_int[0]), .Z(
        DP_mult_105_n579) );
  NAND2_X1 DP_mult_105_U813 ( .A1(DP_mult_105_n579), .A2(DP_mult_105_n615), 
        .ZN(DP_mult_105_n609) );
  BUF_X1 DP_mult_105_U812 ( .A(DP_mult_105_n609), .Z(DP_mult_105_n585) );
  XOR2_X1 DP_mult_105_U811 ( .A(DP_b_int[11]), .B(DP_b_int[10]), .Z(
        DP_mult_105_n584) );
  NAND2_X1 DP_mult_105_U810 ( .A1(DP_mult_105_n584), .A2(DP_mult_105_n620), 
        .ZN(DP_mult_105_n614) );
  XNOR2_X1 DP_mult_105_U809 ( .A(DP_b_int[3]), .B(DP_b_int[4]), .ZN(
        DP_mult_105_n616) );
  XNOR2_X1 DP_mult_105_U808 ( .A(DP_b_int[7]), .B(DP_b_int[8]), .ZN(
        DP_mult_105_n618) );
  XNOR2_X1 DP_mult_105_U807 ( .A(DP_b_int[9]), .B(DP_b_int[10]), .ZN(
        DP_mult_105_n619) );
  XNOR2_X1 DP_mult_105_U806 ( .A(DP_b_int[1]), .B(DP_b_int[2]), .ZN(
        DP_mult_105_n615) );
  XNOR2_X1 DP_mult_105_U805 ( .A(DP_b_int[5]), .B(DP_b_int[6]), .ZN(
        DP_mult_105_n617) );
  INV_X1 DP_mult_105_U804 ( .A(DP_mult_105_n586), .ZN(DP_mult_105_n24) );
  INV_X1 DP_mult_105_U803 ( .A(DP_mult_105_n588), .ZN(DP_mult_105_n69) );
  INV_X1 DP_mult_105_U802 ( .A(DP_mult_105_n589), .ZN(DP_mult_105_n87) );
  INV_X1 DP_mult_105_U801 ( .A(DP_mult_105_n590), .ZN(DP_mult_105_n103) );
  INV_X1 DP_mult_105_U800 ( .A(DP_mult_105_n604), .ZN(DP_mult_105_n598) );
  INV_X1 DP_mult_105_U799 ( .A(DP_mult_105_n605), .ZN(DP_mult_105_n599) );
  INV_X1 DP_mult_105_U798 ( .A(DP_mult_105_n608), .ZN(DP_mult_105_n602) );
  XNOR2_X1 DP_mult_105_U797 ( .A(DP_mult_105_n607), .B(DP_mult_105_n111), .ZN(
        DP_mult_105_n550) );
  OAI22_X1 DP_mult_105_U796 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n562), 
        .B1(DP_mult_105_n561), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n479) );
  OAI22_X1 DP_mult_105_U795 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n550), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n549), .ZN(DP_mult_105_n467) );
  XNOR2_X1 DP_mult_105_U794 ( .A(DP_mult_105_n604), .B(DP_mult_105_n111), .ZN(
        DP_mult_105_n508) );
  OAI22_X1 DP_mult_105_U793 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n520), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n519), .ZN(DP_mult_105_n439) );
  OAI22_X1 DP_mult_105_U792 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n508), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n507), .ZN(DP_mult_105_n428) );
  NAND2_X1 DP_mult_105_U791 ( .A1(DP_mult_105_n35), .A2(DP_mult_105_n605), 
        .ZN(DP_mult_105_n523) );
  INV_X1 DP_mult_105_U790 ( .A(DP_mult_105_n111), .ZN(DP_mult_105_n35) );
  NAND2_X1 DP_mult_105_U789 ( .A1(DP_mult_105_n35), .A2(DP_mult_105_n604), 
        .ZN(DP_mult_105_n509) );
  NAND2_X1 DP_mult_105_U788 ( .A1(DP_mult_105_n109), .A2(DP_mult_105_n606), 
        .ZN(DP_mult_105_n537) );
  INV_X1 DP_mult_105_U787 ( .A(DP_mult_105_n111), .ZN(DP_mult_105_n109) );
  NAND2_X1 DP_mult_105_U786 ( .A1(DP_mult_105_n109), .A2(DP_mult_105_n608), 
        .ZN(DP_mult_105_n565) );
  XNOR2_X1 DP_mult_105_U785 ( .A(DP_mult_105_n605), .B(DP_mult_105_n573), .ZN(
        DP_mult_105_n517) );
  OAI22_X1 DP_mult_105_U784 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n505), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n504), .ZN(DP_mult_105_n425) );
  OAI22_X1 DP_mult_105_U783 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n493), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n492), .ZN(DP_mult_105_n414) );
  XNOR2_X1 DP_mult_105_U782 ( .A(DP_mult_105_n603), .B(DP_mult_105_n111), .ZN(
        DP_mult_105_n494) );
  OAI22_X1 DP_mult_105_U781 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n506), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n505), .ZN(DP_mult_105_n426) );
  OAI22_X1 DP_mult_105_U780 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n494), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n493), .ZN(DP_mult_105_n415) );
  XNOR2_X1 DP_mult_105_U779 ( .A(DP_mult_105_n608), .B(DP_mult_105_n577), .ZN(
        DP_mult_105_n563) );
  XNOR2_X1 DP_mult_105_U778 ( .A(DP_mult_105_n608), .B(DP_mult_105_n576), .ZN(
        DP_mult_105_n562) );
  XNOR2_X1 DP_mult_105_U777 ( .A(DP_mult_105_n608), .B(DP_mult_105_n575), .ZN(
        DP_mult_105_n561) );
  XNOR2_X1 DP_mult_105_U776 ( .A(DP_mult_105_n603), .B(DP_mult_105_n574), .ZN(
        DP_mult_105_n490) );
  XNOR2_X1 DP_mult_105_U775 ( .A(DP_mult_105_n603), .B(DP_mult_105_n573), .ZN(
        DP_mult_105_n489) );
  XNOR2_X1 DP_mult_105_U774 ( .A(DP_mult_105_n603), .B(DP_mult_105_n576), .ZN(
        DP_mult_105_n492) );
  XNOR2_X1 DP_mult_105_U773 ( .A(DP_mult_105_n603), .B(DP_mult_105_n575), .ZN(
        DP_mult_105_n491) );
  XNOR2_X1 DP_mult_105_U772 ( .A(DP_mult_105_n603), .B(DP_mult_105_n572), .ZN(
        DP_mult_105_n488) );
  XNOR2_X1 DP_mult_105_U771 ( .A(DP_mult_105_n603), .B(DP_w_7_), .ZN(
        DP_mult_105_n487) );
  XNOR2_X1 DP_mult_105_U770 ( .A(DP_mult_105_n603), .B(DP_mult_105_n577), .ZN(
        DP_mult_105_n493) );
  XNOR2_X1 DP_mult_105_U769 ( .A(DP_mult_105_n604), .B(DP_w_7_), .ZN(
        DP_mult_105_n501) );
  XNOR2_X1 DP_mult_105_U768 ( .A(DP_mult_105_n604), .B(DP_mult_105_n574), .ZN(
        DP_mult_105_n504) );
  XNOR2_X1 DP_mult_105_U767 ( .A(DP_mult_105_n604), .B(DP_mult_105_n572), .ZN(
        DP_mult_105_n502) );
  XNOR2_X1 DP_mult_105_U766 ( .A(DP_mult_105_n604), .B(DP_mult_105_n573), .ZN(
        DP_mult_105_n503) );
  XNOR2_X1 DP_mult_105_U765 ( .A(DP_mult_105_n605), .B(DP_mult_105_n577), .ZN(
        DP_mult_105_n521) );
  XNOR2_X1 DP_mult_105_U764 ( .A(DP_mult_105_n604), .B(DP_mult_105_n575), .ZN(
        DP_mult_105_n505) );
  XNOR2_X1 DP_mult_105_U763 ( .A(DP_mult_105_n605), .B(DP_mult_105_n576), .ZN(
        DP_mult_105_n520) );
  XNOR2_X1 DP_mult_105_U762 ( .A(DP_mult_105_n604), .B(DP_mult_105_n577), .ZN(
        DP_mult_105_n507) );
  XNOR2_X1 DP_mult_105_U761 ( .A(DP_mult_105_n604), .B(DP_mult_105_n576), .ZN(
        DP_mult_105_n506) );
  XNOR2_X1 DP_mult_105_U760 ( .A(DP_mult_105_n605), .B(DP_mult_105_n575), .ZN(
        DP_mult_105_n519) );
  XNOR2_X1 DP_mult_105_U759 ( .A(DP_mult_105_n605), .B(DP_mult_105_n574), .ZN(
        DP_mult_105_n518) );
  XNOR2_X1 DP_mult_105_U758 ( .A(DP_mult_105_n606), .B(DP_mult_105_n577), .ZN(
        DP_mult_105_n535) );
  XNOR2_X1 DP_mult_105_U757 ( .A(DP_mult_105_n606), .B(DP_mult_105_n576), .ZN(
        DP_mult_105_n534) );
  XNOR2_X1 DP_mult_105_U756 ( .A(DP_mult_105_n606), .B(DP_mult_105_n575), .ZN(
        DP_mult_105_n533) );
  XNOR2_X1 DP_mult_105_U755 ( .A(DP_mult_105_n606), .B(DP_mult_105_n574), .ZN(
        DP_mult_105_n532) );
  XNOR2_X1 DP_mult_105_U754 ( .A(DP_mult_105_n607), .B(DP_mult_105_n577), .ZN(
        DP_mult_105_n549) );
  XNOR2_X1 DP_mult_105_U753 ( .A(DP_mult_105_n607), .B(DP_mult_105_n576), .ZN(
        DP_mult_105_n548) );
  XNOR2_X1 DP_mult_105_U752 ( .A(DP_mult_105_n607), .B(DP_mult_105_n575), .ZN(
        DP_mult_105_n547) );
  XNOR2_X1 DP_mult_105_U751 ( .A(DP_mult_105_n605), .B(DP_mult_105_n111), .ZN(
        DP_mult_105_n522) );
  OAI22_X1 DP_mult_105_U750 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n534), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n533), .ZN(DP_mult_105_n452) );
  OAI22_X1 DP_mult_105_U749 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n522), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n521), .ZN(DP_mult_105_n441) );
  BUF_X1 DP_mult_105_U748 ( .A(DP_mult_105_n618), .Z(DP_mult_105_n594) );
  BUF_X1 DP_mult_105_U747 ( .A(DP_mult_105_n617), .Z(DP_mult_105_n593) );
  XNOR2_X1 DP_mult_105_U746 ( .A(DP_mult_105_n608), .B(DP_mult_105_n111), .ZN(
        DP_mult_105_n564) );
  OAI22_X1 DP_mult_105_U745 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n602), 
        .B1(DP_mult_105_n565), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n403) );
  OAI22_X1 DP_mult_105_U744 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n564), 
        .B1(DP_mult_105_n563), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n481) );
  INV_X1 DP_mult_105_U743 ( .A(DP_mult_105_n603), .ZN(DP_mult_105_n597) );
  OAI22_X1 DP_mult_105_U742 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n597), 
        .B1(DP_mult_105_n495), .B2(DP_mult_105_n591), .ZN(DP_mult_105_n398) );
  BUF_X1 DP_mult_105_U741 ( .A(DP_mult_105_n619), .Z(DP_mult_105_n595) );
  BUF_X1 DP_mult_105_U740 ( .A(DP_mult_105_n616), .Z(DP_mult_105_n592) );
  BUF_X1 DP_mult_105_U739 ( .A(DP_mult_105_n615), .Z(DP_mult_105_n591) );
  OAI22_X1 DP_mult_105_U738 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n503), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n502), .ZN(DP_mult_105_n423) );
  OAI22_X1 DP_mult_105_U737 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n492), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n491), .ZN(DP_mult_105_n413) );
  INV_X1 DP_mult_105_U736 ( .A(DP_mult_105_n482), .ZN(DP_mult_105_n10) );
  INV_X1 DP_mult_105_U735 ( .A(DP_mult_105_n585), .ZN(DP_mult_105_n8) );
  OAI21_X1 DP_mult_105_U734 ( .B1(DP_mult_105_n8), .B2(DP_mult_105_n14), .A(
        DP_mult_105_n10), .ZN(DP_mult_105_n404) );
  OAI22_X1 DP_mult_105_U733 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n504), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n503), .ZN(DP_mult_105_n424) );
  NAND2_X1 DP_mult_105_U732 ( .A1(DP_mult_105_n109), .A2(DP_mult_105_n607), 
        .ZN(DP_mult_105_n551) );
  INV_X1 DP_mult_105_U731 ( .A(DP_mult_105_n607), .ZN(DP_mult_105_n601) );
  OAI22_X1 DP_mult_105_U730 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n601), 
        .B1(DP_mult_105_n551), .B2(DP_mult_105_n595), .ZN(DP_mult_105_n402) );
  OAI22_X1 DP_mult_105_U729 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n563), 
        .B1(DP_mult_105_n562), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n480) );
  OAI22_X1 DP_mult_105_U728 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n499), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n498), .ZN(DP_mult_105_n419) );
  OAI22_X1 DP_mult_105_U727 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n487), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n486), .ZN(DP_mult_105_n408) );
  OAI22_X1 DP_mult_105_U726 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n545), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n544), .ZN(DP_mult_105_n462) );
  OAI22_X1 DP_mult_105_U725 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n521), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n520), .ZN(DP_mult_105_n440) );
  OAI22_X1 DP_mult_105_U724 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n526), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n525), .ZN(DP_mult_105_n444) );
  OAI22_X1 DP_mult_105_U723 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n490), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n489), .ZN(DP_mult_105_n411) );
  OAI22_X1 DP_mult_105_U722 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n498), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n497), .ZN(DP_mult_105_n418) );
  OAI22_X1 DP_mult_105_U721 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n486), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n485), .ZN(DP_mult_105_n407) );
  OAI22_X1 DP_mult_105_U720 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n519), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n518), .ZN(DP_mult_105_n438) );
  OAI22_X1 DP_mult_105_U719 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n507), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n506), .ZN(DP_mult_105_n427) );
  OAI21_X1 DP_mult_105_U718 ( .B1(DP_mult_105_n69), .B2(DP_mult_105_n77), .A(
        DP_mult_105_n73), .ZN(DP_mult_105_n443) );
  OAI22_X1 DP_mult_105_U717 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n512), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n511), .ZN(DP_mult_105_n431) );
  OAI22_X1 DP_mult_105_U716 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n501), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n500), .ZN(DP_mult_105_n421) );
  OAI22_X1 DP_mult_105_U715 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n489), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n488), .ZN(DP_mult_105_n410) );
  OAI22_X1 DP_mult_105_U714 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n558), 
        .B1(DP_mult_105_n557), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n475) );
  OAI22_X1 DP_mult_105_U713 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n546), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n545), .ZN(DP_mult_105_n463) );
  OAI22_X1 DP_mult_105_U712 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n599), 
        .B1(DP_mult_105_n523), .B2(DP_mult_105_n593), .ZN(DP_mult_105_n400) );
  OAI22_X1 DP_mult_105_U711 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n513), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n512), .ZN(DP_mult_105_n432) );
  OAI22_X1 DP_mult_105_U710 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n500), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n499), .ZN(DP_mult_105_n420) );
  OAI22_X1 DP_mult_105_U709 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n488), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n487), .ZN(DP_mult_105_n409) );
  OAI22_X1 DP_mult_105_U708 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n542), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n541), .ZN(DP_mult_105_n459) );
  OAI22_X1 DP_mult_105_U707 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n518), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n517), .ZN(DP_mult_105_n437) );
  OAI22_X1 DP_mult_105_U706 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n528), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n527), .ZN(DP_mult_105_n446) );
  OAI22_X1 DP_mult_105_U705 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n516), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n515), .ZN(DP_mult_105_n435) );
  OAI21_X1 DP_mult_105_U704 ( .B1(DP_mult_105_n87), .B2(DP_mult_105_n93), .A(
        DP_mult_105_n746), .ZN(DP_mult_105_n456) );
  OAI22_X1 DP_mult_105_U703 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n514), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n513), .ZN(DP_mult_105_n433) );
  OAI22_X1 DP_mult_105_U702 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n502), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n501), .ZN(DP_mult_105_n422) );
  OAI22_X1 DP_mult_105_U701 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n543), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n542), .ZN(DP_mult_105_n460) );
  OAI22_X1 DP_mult_105_U700 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n531), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n530), .ZN(DP_mult_105_n449) );
  OAI22_X1 DP_mult_105_U699 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n533), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n532), .ZN(DP_mult_105_n451) );
  OAI22_X1 DP_mult_105_U698 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n544), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n543), .ZN(DP_mult_105_n461) );
  OAI22_X1 DP_mult_105_U697 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n532), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n531), .ZN(DP_mult_105_n450) );
  OAI22_X1 DP_mult_105_U696 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n598), 
        .B1(DP_mult_105_n509), .B2(DP_mult_105_n592), .ZN(DP_mult_105_n399) );
  XNOR2_X1 DP_mult_105_U695 ( .A(DP_mult_105_n608), .B(DP_w_7_), .ZN(
        DP_mult_105_n557) );
  XNOR2_X1 DP_mult_105_U694 ( .A(DP_mult_105_n606), .B(DP_w_7_), .ZN(
        DP_mult_105_n529) );
  XNOR2_X1 DP_mult_105_U693 ( .A(DP_mult_105_n605), .B(DP_mult_105_n572), .ZN(
        DP_mult_105_n516) );
  XNOR2_X1 DP_mult_105_U692 ( .A(DP_mult_105_n606), .B(DP_mult_105_n111), .ZN(
        DP_mult_105_n536) );
  OAI22_X1 DP_mult_105_U691 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n560), 
        .B1(DP_mult_105_n559), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n477) );
  OAI22_X1 DP_mult_105_U690 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n536), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n535), .ZN(DP_mult_105_n454) );
  XNOR2_X1 DP_mult_105_U689 ( .A(DP_mult_105_n608), .B(DP_mult_105_n574), .ZN(
        DP_mult_105_n560) );
  XNOR2_X1 DP_mult_105_U688 ( .A(DP_mult_105_n608), .B(DP_mult_105_n573), .ZN(
        DP_mult_105_n559) );
  XNOR2_X1 DP_mult_105_U687 ( .A(DP_mult_105_n608), .B(DP_mult_105_n572), .ZN(
        DP_mult_105_n558) );
  XNOR2_X1 DP_mult_105_U686 ( .A(DP_mult_105_n605), .B(DP_w_7_), .ZN(
        DP_mult_105_n515) );
  XNOR2_X1 DP_mult_105_U685 ( .A(DP_mult_105_n606), .B(DP_mult_105_n573), .ZN(
        DP_mult_105_n531) );
  XNOR2_X1 DP_mult_105_U684 ( .A(DP_mult_105_n606), .B(DP_mult_105_n572), .ZN(
        DP_mult_105_n530) );
  XNOR2_X1 DP_mult_105_U683 ( .A(DP_mult_105_n607), .B(DP_mult_105_n574), .ZN(
        DP_mult_105_n546) );
  XNOR2_X1 DP_mult_105_U682 ( .A(DP_mult_105_n607), .B(DP_mult_105_n573), .ZN(
        DP_mult_105_n545) );
  XNOR2_X1 DP_mult_105_U681 ( .A(DP_mult_105_n607), .B(DP_mult_105_n572), .ZN(
        DP_mult_105_n544) );
  XNOR2_X1 DP_mult_105_U680 ( .A(DP_mult_105_n607), .B(DP_w_7_), .ZN(
        DP_mult_105_n543) );
  OAI22_X1 DP_mult_105_U679 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n541), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n540), .ZN(DP_mult_105_n458) );
  OAI22_X1 DP_mult_105_U678 ( .A1(DP_mult_105_n587), .A2(DP_mult_105_n515), 
        .B1(DP_mult_105_n593), .B2(DP_mult_105_n514), .ZN(DP_mult_105_n434) );
  OR2_X1 DP_mult_105_U677 ( .A1(DP_mult_105_n413), .A2(DP_mult_105_n424), .ZN(
        DP_mult_105_n336) );
  OAI22_X1 DP_mult_105_U676 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n491), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n490), .ZN(DP_mult_105_n412) );
  OAI22_X1 DP_mult_105_U675 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n559), 
        .B1(DP_mult_105_n558), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n476) );
  OAI22_X1 DP_mult_105_U674 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n547), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n546), .ZN(DP_mult_105_n464) );
  OAI22_X1 DP_mult_105_U673 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n535), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n534), .ZN(DP_mult_105_n453) );
  INV_X1 DP_mult_105_U672 ( .A(DP_mult_105_n587), .ZN(DP_mult_105_n40) );
  OAI21_X1 DP_mult_105_U671 ( .B1(DP_mult_105_n40), .B2(DP_mult_105_n57), .A(
        DP_mult_105_n48), .ZN(DP_mult_105_n430) );
  OAI22_X1 DP_mult_105_U670 ( .A1(DP_mult_105_n590), .A2(DP_mult_105_n561), 
        .B1(DP_mult_105_n560), .B2(DP_mult_105_n596), .ZN(DP_mult_105_n478) );
  OAI22_X1 DP_mult_105_U669 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n549), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n548), .ZN(DP_mult_105_n466) );
  INV_X1 DP_mult_105_U668 ( .A(DP_mult_105_n606), .ZN(DP_mult_105_n600) );
  OAI22_X1 DP_mult_105_U667 ( .A1(DP_mult_105_n589), .A2(DP_mult_105_n548), 
        .B1(DP_mult_105_n595), .B2(DP_mult_105_n547), .ZN(DP_mult_105_n465) );
  OAI22_X1 DP_mult_105_U666 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n600), 
        .B1(DP_mult_105_n537), .B2(DP_mult_105_n594), .ZN(DP_mult_105_n401) );
  INV_X1 DP_mult_105_U665 ( .A(DP_mult_105_n284), .ZN(DP_mult_105_n285) );
  OAI22_X1 DP_mult_105_U664 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n485), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n484), .ZN(DP_mult_105_n406) );
  OAI21_X1 DP_mult_105_U663 ( .B1(DP_mult_105_n24), .B2(DP_mult_105_n30), .A(
        DP_mult_105_n26), .ZN(DP_mult_105_n417) );
  OAI22_X1 DP_mult_105_U662 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n484), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n483), .ZN(DP_mult_105_n405) );
  OAI22_X1 DP_mult_105_U661 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n527), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n526), .ZN(DP_mult_105_n445) );
  OAI22_X1 DP_mult_105_U660 ( .A1(DP_mult_105_n588), .A2(DP_mult_105_n530), 
        .B1(DP_mult_105_n594), .B2(DP_mult_105_n529), .ZN(DP_mult_105_n448) );
  OAI22_X1 DP_mult_105_U659 ( .A1(DP_mult_105_n586), .A2(DP_mult_105_n497), 
        .B1(DP_mult_105_n592), .B2(DP_mult_105_n496), .ZN(DP_mult_105_n284) );
  INV_X1 DP_mult_105_U658 ( .A(DP_mult_105_n595), .ZN(DP_mult_105_n93) );
  INV_X1 DP_mult_105_U657 ( .A(DP_mult_105_n594), .ZN(DP_mult_105_n77) );
  INV_X1 DP_mult_105_U656 ( .A(DP_mult_105_n496), .ZN(DP_mult_105_n26) );
  BUF_X4 DP_mult_105_U655 ( .A(DP_w_0_), .Z(DP_mult_105_n111) );
  NOR2_X1 DP_mult_105_U654 ( .A1(DP_mult_105_n397), .A2(DP_mult_105_n402), 
        .ZN(DP_mult_105_n258) );
  NAND2_X1 DP_mult_105_U653 ( .A1(DP_mult_105_n397), .A2(DP_mult_105_n402), 
        .ZN(DP_mult_105_n259) );
  NAND2_X1 DP_mult_105_U652 ( .A1(DP_mult_105_n404), .A2(DP_mult_105_n278), 
        .ZN(DP_mult_105_n129) );
  INV_X1 DP_mult_105_U651 ( .A(DP_mult_105_n278), .ZN(DP_mult_105_n279) );
  BUF_X1 DP_mult_105_U650 ( .A(DP_w_1_), .Z(DP_mult_105_n577) );
  AOI21_X1 DP_mult_105_U649 ( .B1(DP_mult_105_n668), .B2(DP_mult_105_n665), 
        .A(DP_mult_105_n672), .ZN(DP_mult_105_n260) );
  NOR2_X1 DP_mult_105_U648 ( .A1(DP_mult_105_n280), .A2(DP_mult_105_n279), 
        .ZN(DP_mult_105_n134) );
  NOR2_X1 DP_mult_105_U647 ( .A1(DP_mult_105_n404), .A2(DP_mult_105_n278), 
        .ZN(DP_mult_105_n128) );
  OR2_X1 DP_mult_105_U646 ( .A1(DP_mult_105_n375), .A2(DP_mult_105_n377), .ZN(
        DP_mult_105_n709) );
  INV_X1 DP_mult_105_U645 ( .A(DP_mult_105_n524), .ZN(DP_mult_105_n73) );
  INV_X1 DP_mult_105_U644 ( .A(DP_mult_105_n510), .ZN(DP_mult_105_n48) );
  NAND2_X1 DP_mult_105_U643 ( .A1(DP_mult_105_n395), .A2(DP_mult_105_n670), 
        .ZN(DP_mult_105_n256) );
  NAND2_X1 DP_mult_105_U642 ( .A1(DP_mult_105_n391), .A2(DP_mult_105_n394), 
        .ZN(DP_mult_105_n254) );
  NAND2_X1 DP_mult_105_U641 ( .A1(DP_mult_105_n387), .A2(DP_mult_105_n390), 
        .ZN(DP_mult_105_n249) );
  NAND2_X1 DP_mult_105_U640 ( .A1(DP_mult_105_n281), .A2(DP_mult_105_n282), 
        .ZN(DP_mult_105_n145) );
  NAND2_X1 DP_mult_105_U639 ( .A1(DP_mult_105_n287), .A2(DP_mult_105_n290), 
        .ZN(DP_mult_105_n165) );
  NAND2_X1 DP_mult_105_U638 ( .A1(DP_mult_105_n283), .A2(DP_mult_105_n286), 
        .ZN(DP_mult_105_n154) );
  INV_X1 DP_mult_105_U637 ( .A(DP_mult_105_n591), .ZN(DP_mult_105_n14) );
  INV_X1 DP_mult_105_U636 ( .A(DP_mult_105_n592), .ZN(DP_mult_105_n30) );
  NOR2_X1 DP_mult_105_U635 ( .A1(DP_mult_105_n387), .A2(DP_mult_105_n390), 
        .ZN(DP_mult_105_n248) );
  NOR2_X1 DP_mult_105_U634 ( .A1(DP_mult_105_n395), .A2(DP_mult_105_n670), 
        .ZN(DP_mult_105_n255) );
  AOI21_X1 DP_mult_105_U633 ( .B1(DP_mult_105_n703), .B2(DP_mult_105_n163), 
        .A(DP_mult_105_n139), .ZN(DP_mult_105_n137) );
  NAND2_X1 DP_mult_105_U632 ( .A1(DP_mult_105_n280), .A2(DP_mult_105_n279), 
        .ZN(DP_mult_105_n135) );
  OAI21_X1 DP_mult_105_U631 ( .B1(DP_mult_105_n137), .B2(DP_mult_105_n134), 
        .A(DP_mult_105_n135), .ZN(DP_mult_105_n133) );
  AOI21_X1 DP_mult_105_U630 ( .B1(DP_mult_105_n168), .B2(DP_mult_105_n132), 
        .A(DP_mult_105_n133), .ZN(DP_mult_105_n131) );
  OAI21_X1 DP_mult_105_U629 ( .B1(DP_mult_105_n103), .B2(DP_b_int[11]), .A(
        DP_mult_105_n105), .ZN(DP_mult_105_n469) );
  XNOR2_X1 DP_mult_105_U628 ( .A(DP_mult_105_n413), .B(DP_mult_105_n424), .ZN(
        DP_mult_105_n337) );
  NOR2_X1 DP_mult_105_U627 ( .A1(DP_mult_105_n391), .A2(DP_mult_105_n394), 
        .ZN(DP_mult_105_n253) );
  XNOR2_X1 DP_mult_105_U626 ( .A(DP_mult_105_n376), .B(DP_mult_105_n371), .ZN(
        DP_mult_105_n708) );
  XNOR2_X1 DP_mult_105_U625 ( .A(DP_mult_105_n369), .B(DP_mult_105_n708), .ZN(
        DP_mult_105_n367) );
  XNOR2_X1 DP_mult_105_U624 ( .A(DP_mult_105_n368), .B(DP_mult_105_n363), .ZN(
        DP_mult_105_n707) );
  XNOR2_X1 DP_mult_105_U623 ( .A(DP_mult_105_n361), .B(DP_mult_105_n707), .ZN(
        DP_mult_105_n359) );
  INV_X1 DP_mult_105_U622 ( .A(DP_mult_105_n593), .ZN(DP_mult_105_n57) );
  XNOR2_X1 DP_mult_105_U621 ( .A(DP_mult_105_n350), .B(DP_mult_105_n343), .ZN(
        DP_mult_105_n706) );
  XNOR2_X1 DP_mult_105_U620 ( .A(DP_mult_105_n706), .B(DP_mult_105_n341), .ZN(
        DP_mult_105_n339) );
  BUF_X1 DP_mult_105_U619 ( .A(DP_w_3_), .Z(DP_mult_105_n575) );
  BUF_X1 DP_mult_105_U618 ( .A(DP_w_2_), .Z(DP_mult_105_n576) );
  OAI21_X1 DP_mult_105_U617 ( .B1(DP_mult_105_n250), .B2(DP_mult_105_n248), 
        .A(DP_mult_105_n249), .ZN(DP_mult_105_n247) );
  INV_X1 DP_mult_105_U616 ( .A(DP_mult_105_n145), .ZN(DP_mult_105_n143) );
  AOI21_X1 DP_mult_105_U615 ( .B1(DP_mult_105_n664), .B2(DP_mult_105_n152), 
        .A(DP_mult_105_n143), .ZN(DP_mult_105_n141) );
  INV_X1 DP_mult_105_U614 ( .A(DP_mult_105_n141), .ZN(DP_mult_105_n139) );
  OAI21_X1 DP_mult_105_U613 ( .B1(DP_mult_105_n131), .B2(DP_mult_105_n128), 
        .A(DP_mult_105_n129), .ZN(DP_mult_105_n127) );
  NOR2_X1 DP_mult_105_U612 ( .A1(DP_mult_105_n130), .A2(DP_mult_105_n128), 
        .ZN(DP_mult_105_n126) );
  AND2_X1 DP_mult_105_U611 ( .A1(DP_mult_105_n367), .A2(DP_mult_105_n374), 
        .ZN(DP_mult_105_n705) );
  INV_X1 DP_mult_105_U610 ( .A(DP_mult_105_n165), .ZN(DP_mult_105_n163) );
  INV_X1 DP_mult_105_U609 ( .A(DP_mult_105_n154), .ZN(DP_mult_105_n152) );
  OR2_X1 DP_mult_105_U608 ( .A1(DP_mult_105_n367), .A2(DP_mult_105_n374), .ZN(
        DP_mult_105_n704) );
  NAND2_X1 DP_mult_105_U607 ( .A1(DP_mult_105_n661), .A2(DP_mult_105_n165), 
        .ZN(DP_mult_105_n116) );
  XOR2_X1 DP_mult_105_U606 ( .A(DP_mult_105_n166), .B(DP_mult_105_n116), .Z(
        DP_w_b0_8_) );
  NAND2_X1 DP_mult_105_U605 ( .A1(DP_mult_105_n667), .A2(DP_mult_105_n154), 
        .ZN(DP_mult_105_n115) );
  NAND2_X1 DP_mult_105_U604 ( .A1(DP_mult_105_n664), .A2(DP_mult_105_n145), 
        .ZN(DP_mult_105_n114) );
  XOR2_X1 DP_mult_105_U603 ( .A(DP_mult_105_n146), .B(DP_mult_105_n114), .Z(
        DP_w_b0_10_) );
  NAND2_X1 DP_mult_105_U602 ( .A1(DP_mult_105_n296), .A2(DP_mult_105_n291), 
        .ZN(DP_mult_105_n174) );
  NAND2_X1 DP_mult_105_U601 ( .A1(DP_mult_105_n297), .A2(DP_mult_105_n302), 
        .ZN(DP_mult_105_n183) );
  BUF_X2 DP_mult_105_U600 ( .A(DP_w_8_), .Z(DP_mult_105_n570) );
  BUF_X1 DP_mult_105_U599 ( .A(DP_w_4_), .Z(DP_mult_105_n574) );
  BUF_X1 DP_mult_105_U598 ( .A(DP_w_5_), .Z(DP_mult_105_n573) );
  BUF_X1 DP_mult_105_U597 ( .A(DP_w_6_), .Z(DP_mult_105_n572) );
  OAI21_X1 DP_mult_105_U596 ( .B1(DP_mult_105_n253), .B2(DP_mult_105_n256), 
        .A(DP_mult_105_n254), .ZN(DP_mult_105_n252) );
  NOR2_X1 DP_mult_105_U595 ( .A1(DP_mult_105_n253), .A2(DP_mult_105_n255), 
        .ZN(DP_mult_105_n251) );
  OAI21_X1 DP_mult_105_U594 ( .B1(DP_mult_105_n260), .B2(DP_mult_105_n258), 
        .A(DP_mult_105_n259), .ZN(DP_mult_105_n257) );
  AOI21_X1 DP_mult_105_U593 ( .B1(DP_mult_105_n251), .B2(DP_mult_105_n257), 
        .A(DP_mult_105_n252), .ZN(DP_mult_105_n250) );
  NAND2_X1 DP_mult_105_U592 ( .A1(DP_mult_105_n661), .A2(DP_mult_105_n703), 
        .ZN(DP_mult_105_n136) );
  NOR2_X1 DP_mult_105_U591 ( .A1(DP_mult_105_n136), .A2(DP_mult_105_n134), 
        .ZN(DP_mult_105_n132) );
  NAND2_X1 DP_mult_105_U590 ( .A1(DP_mult_105_n303), .A2(DP_mult_105_n310), 
        .ZN(DP_mult_105_n192) );
  NOR2_X1 DP_mult_105_U589 ( .A1(DP_mult_105_n303), .A2(DP_mult_105_n310), 
        .ZN(DP_mult_105_n191) );
  INV_X1 DP_mult_105_U588 ( .A(DP_mult_105_n675), .ZN(DP_mult_105_n203) );
  INV_X1 DP_mult_105_U587 ( .A(DP_mult_105_n198), .ZN(DP_mult_105_n273) );
  INV_X1 DP_mult_105_U586 ( .A(DP_mult_105_n192), .ZN(DP_mult_105_n190) );
  AND2_X1 DP_mult_105_U585 ( .A1(DP_mult_105_n667), .A2(DP_mult_105_n664), 
        .ZN(DP_mult_105_n703) );
  INV_X1 DP_mult_105_U584 ( .A(DP_mult_105_n661), .ZN(DP_mult_105_n161) );
  INV_X1 DP_mult_105_U583 ( .A(DP_mult_105_n161), .ZN(DP_mult_105_n160) );
  INV_X1 DP_mult_105_U582 ( .A(DP_mult_105_n183), .ZN(DP_mult_105_n181) );
  INV_X1 DP_mult_105_U581 ( .A(DP_mult_105_n667), .ZN(DP_mult_105_n149) );
  AND2_X1 DP_mult_105_U580 ( .A1(DP_mult_105_n740), .A2(DP_mult_105_n226), 
        .ZN(DP_mult_105_n702) );
  XOR2_X1 DP_mult_105_U579 ( .A(DP_mult_105_n227), .B(DP_mult_105_n702), .Z(
        DP_w_b0_0_) );
  INV_X1 DP_mult_105_U578 ( .A(DP_mult_105_n152), .ZN(DP_mult_105_n150) );
  OAI21_X1 DP_mult_105_U577 ( .B1(DP_mult_105_n159), .B2(DP_mult_105_n149), 
        .A(DP_mult_105_n150), .ZN(DP_mult_105_n148) );
  NAND2_X1 DP_mult_105_U576 ( .A1(DP_mult_105_n167), .A2(DP_mult_105_n132), 
        .ZN(DP_mult_105_n130) );
  NAND2_X1 DP_mult_105_U575 ( .A1(DP_mult_105_n666), .A2(DP_mult_105_n183), 
        .ZN(DP_mult_105_n118) );
  NAND2_X1 DP_mult_105_U574 ( .A1(DP_mult_105_n663), .A2(DP_mult_105_n174), 
        .ZN(DP_mult_105_n117) );
  XOR2_X1 DP_mult_105_U573 ( .A(DP_mult_105_n175), .B(DP_mult_105_n117), .Z(
        DP_w_b0_7_) );
  OR2_X1 DP_mult_105_U572 ( .A1(DP_mult_105_n214), .A2(DP_mult_105_n219), .ZN(
        DP_mult_105_n721) );
  INV_X1 DP_mult_105_U571 ( .A(DP_mult_105_n174), .ZN(DP_mult_105_n172) );
  AOI21_X1 DP_mult_105_U570 ( .B1(DP_mult_105_n181), .B2(DP_mult_105_n663), 
        .A(DP_mult_105_n172), .ZN(DP_mult_105_n170) );
  OAI21_X1 DP_mult_105_U569 ( .B1(DP_mult_105_n169), .B2(DP_mult_105_n192), 
        .A(DP_mult_105_n170), .ZN(DP_mult_105_n168) );
  AOI21_X1 DP_mult_105_U568 ( .B1(DP_mult_105_n168), .B2(DP_mult_105_n160), 
        .A(DP_mult_105_n163), .ZN(DP_mult_105_n159) );
  NOR2_X1 DP_mult_105_U567 ( .A1(DP_mult_105_n191), .A2(DP_mult_105_n169), 
        .ZN(DP_mult_105_n167) );
  INV_X1 DP_mult_105_U566 ( .A(DP_mult_105_n191), .ZN(DP_mult_105_n185) );
  INV_X1 DP_mult_105_U565 ( .A(DP_mult_105_n721), .ZN(DP_mult_105_n212) );
  INV_X1 DP_mult_105_U564 ( .A(DP_mult_105_n159), .ZN(DP_mult_105_n157) );
  INV_X1 DP_mult_105_U563 ( .A(DP_mult_105_n721), .ZN(DP_mult_105_n208) );
  NOR2_X1 DP_mult_105_U562 ( .A1(DP_mult_105_n191), .A2(DP_mult_105_n178), 
        .ZN(DP_mult_105_n176) );
  NOR2_X1 DP_mult_105_U561 ( .A1(DP_mult_105_n158), .A2(DP_mult_105_n149), 
        .ZN(DP_mult_105_n147) );
  INV_X1 DP_mult_105_U560 ( .A(DP_mult_105_n666), .ZN(DP_mult_105_n178) );
  NAND2_X1 DP_mult_105_U559 ( .A1(DP_mult_105_n666), .A2(DP_mult_105_n663), 
        .ZN(DP_mult_105_n169) );
  INV_X1 DP_mult_105_U558 ( .A(DP_mult_105_n181), .ZN(DP_mult_105_n179) );
  OAI21_X1 DP_mult_105_U557 ( .B1(DP_mult_105_n192), .B2(DP_mult_105_n178), 
        .A(DP_mult_105_n179), .ZN(DP_mult_105_n177) );
  NAND2_X1 DP_mult_105_U556 ( .A1(DP_mult_105_n167), .A2(DP_mult_105_n160), 
        .ZN(DP_mult_105_n158) );
  INV_X1 DP_mult_105_U555 ( .A(DP_mult_105_n158), .ZN(DP_mult_105_n156) );
  BUF_X1 DP_mult_105_U554 ( .A(DP_b_int[0]), .Z(DP_mult_105_n603) );
  BUF_X1 DP_mult_105_U553 ( .A(DP_b_int[2]), .Z(DP_mult_105_n604) );
  BUF_X1 DP_mult_105_U552 ( .A(DP_b_int[8]), .Z(DP_mult_105_n607) );
  BUF_X1 DP_mult_105_U551 ( .A(DP_mult_105_n620), .Z(DP_mult_105_n596) );
  OR2_X1 DP_mult_105_U550 ( .A1(DP_mult_105_n111), .A2(DP_mult_105_n597), .ZN(
        DP_mult_105_n495) );
  AND2_X1 DP_mult_105_U549 ( .A1(DP_mult_105_n111), .A2(DP_mult_105_n14), .ZN(
        DP_mult_105_n701) );
  AND2_X1 DP_mult_105_U548 ( .A1(DP_mult_105_n111), .A2(DP_mult_105_n30), .ZN(
        DP_mult_105_n700) );
  AND2_X1 DP_mult_105_U547 ( .A1(DP_mult_105_n111), .A2(DP_mult_105_n57), .ZN(
        DP_mult_105_n699) );
  CLKBUF_X1 DP_mult_105_U546 ( .A(DP_mult_105_n698), .Z(DP_mult_105_n697) );
  CLKBUF_X1 DP_mult_105_U545 ( .A(DP_w_9_), .Z(DP_mult_105_n569) );
  NAND3_X1 DP_mult_105_U544 ( .A1(DP_mult_105_n694), .A2(DP_mult_105_n695), 
        .A3(DP_mult_105_n696), .ZN(DP_mult_105_n360) );
  NAND2_X1 DP_mult_105_U543 ( .A1(DP_mult_105_n370), .A2(DP_mult_105_n701), 
        .ZN(DP_mult_105_n696) );
  NAND2_X1 DP_mult_105_U542 ( .A1(DP_mult_105_n365), .A2(DP_mult_105_n701), 
        .ZN(DP_mult_105_n695) );
  NAND2_X1 DP_mult_105_U541 ( .A1(DP_mult_105_n365), .A2(DP_mult_105_n370), 
        .ZN(DP_mult_105_n694) );
  NAND3_X1 DP_mult_105_U540 ( .A1(DP_mult_105_n691), .A2(DP_mult_105_n692), 
        .A3(DP_mult_105_n693), .ZN(DP_mult_105_n328) );
  NAND2_X1 DP_mult_105_U539 ( .A1(DP_mult_105_n340), .A2(DP_mult_105_n333), 
        .ZN(DP_mult_105_n693) );
  NAND2_X1 DP_mult_105_U538 ( .A1(DP_mult_105_n331), .A2(DP_mult_105_n333), 
        .ZN(DP_mult_105_n692) );
  NAND2_X1 DP_mult_105_U537 ( .A1(DP_mult_105_n331), .A2(DP_mult_105_n340), 
        .ZN(DP_mult_105_n691) );
  XNOR2_X1 DP_mult_105_U536 ( .A(DP_mult_105_n340), .B(DP_mult_105_n333), .ZN(
        DP_mult_105_n690) );
  XNOR2_X1 DP_mult_105_U535 ( .A(DP_mult_105_n331), .B(DP_mult_105_n690), .ZN(
        DP_mult_105_n329) );
  BUF_X2 DP_mult_105_U534 ( .A(DP_w_12_), .Z(DP_mult_105_n566) );
  BUF_X1 DP_mult_105_U533 ( .A(DP_mult_105_n364), .Z(DP_mult_105_n688) );
  BUF_X1 DP_mult_105_U532 ( .A(DP_mult_105_n193), .Z(DP_mult_105_n698) );
  NAND3_X1 DP_mult_105_U531 ( .A1(DP_mult_105_n685), .A2(DP_mult_105_n686), 
        .A3(DP_mult_105_n687), .ZN(DP_mult_105_n310) );
  NAND2_X1 DP_mult_105_U530 ( .A1(DP_mult_105_n315), .A2(DP_mult_105_n313), 
        .ZN(DP_mult_105_n687) );
  NAND2_X1 DP_mult_105_U529 ( .A1(DP_mult_105_n320), .A2(DP_mult_105_n313), 
        .ZN(DP_mult_105_n686) );
  NAND2_X1 DP_mult_105_U528 ( .A1(DP_mult_105_n320), .A2(DP_mult_105_n315), 
        .ZN(DP_mult_105_n685) );
  NAND3_X1 DP_mult_105_U527 ( .A1(DP_mult_105_n682), .A2(DP_mult_105_n683), 
        .A3(DP_mult_105_n684), .ZN(DP_mult_105_n312) );
  NAND2_X1 DP_mult_105_U526 ( .A1(DP_mult_105_n324), .A2(DP_mult_105_n317), 
        .ZN(DP_mult_105_n684) );
  NAND2_X1 DP_mult_105_U525 ( .A1(DP_mult_105_n322), .A2(DP_mult_105_n317), 
        .ZN(DP_mult_105_n683) );
  NAND2_X1 DP_mult_105_U524 ( .A1(DP_mult_105_n322), .A2(DP_mult_105_n324), 
        .ZN(DP_mult_105_n682) );
  CLKBUF_X1 DP_mult_105_U523 ( .A(DP_mult_105_n365), .Z(DP_mult_105_n681) );
  BUF_X1 DP_mult_105_U522 ( .A(DP_mult_105_n221), .Z(DP_mult_105_n689) );
  AND2_X1 DP_mult_105_U521 ( .A1(DP_mult_105_n273), .A2(DP_mult_105_n199), 
        .ZN(DP_mult_105_n680) );
  XNOR2_X1 DP_mult_105_U520 ( .A(DP_mult_105_n200), .B(DP_mult_105_n680), .ZN(
        DP_w_b0_4_) );
  XNOR2_X1 DP_mult_105_U519 ( .A(DP_mult_105_n320), .B(DP_mult_105_n315), .ZN(
        DP_mult_105_n679) );
  XNOR2_X1 DP_mult_105_U518 ( .A(DP_mult_105_n679), .B(DP_mult_105_n313), .ZN(
        DP_mult_105_n311) );
  XNOR2_X1 DP_mult_105_U517 ( .A(DP_mult_105_n322), .B(DP_mult_105_n324), .ZN(
        DP_mult_105_n678) );
  XNOR2_X1 DP_mult_105_U516 ( .A(DP_mult_105_n678), .B(DP_mult_105_n317), .ZN(
        DP_mult_105_n313) );
  CLKBUF_X1 DP_mult_105_U515 ( .A(DP_mult_105_n355), .Z(DP_mult_105_n729) );
  XNOR2_X1 DP_mult_105_U514 ( .A(DP_mult_105_n370), .B(DP_mult_105_n701), .ZN(
        DP_mult_105_n677) );
  XNOR2_X1 DP_mult_105_U513 ( .A(DP_mult_105_n681), .B(DP_mult_105_n677), .ZN(
        DP_mult_105_n361) );
  XOR2_X1 DP_mult_105_U512 ( .A(DP_mult_105_n710), .B(DP_mult_105_n326), .Z(
        DP_mult_105_n325) );
  OAI22_X1 DP_mult_105_U511 ( .A1(DP_mult_105_n596), .A2(DP_mult_105_n554), 
        .B1(DP_mult_105_n555), .B2(DP_mult_105_n614), .ZN(DP_mult_105_n472) );
  AND2_X1 DP_mult_105_U510 ( .A1(DP_mult_105_n675), .A2(DP_mult_105_n206), 
        .ZN(DP_mult_105_n676) );
  XNOR2_X1 DP_mult_105_U509 ( .A(DP_mult_105_n207), .B(DP_mult_105_n676), .ZN(
        DP_w_b0_3_) );
  OR2_X1 DP_mult_105_U508 ( .A1(DP_mult_105_n319), .A2(DP_mult_105_n328), .ZN(
        DP_mult_105_n675) );
  OR2_X1 DP_mult_105_U507 ( .A1(DP_mult_105_n381), .A2(DP_mult_105_n386), .ZN(
        DP_mult_105_n674) );
  AND2_X1 DP_mult_105_U506 ( .A1(DP_mult_105_n375), .A2(DP_mult_105_n377), 
        .ZN(DP_mult_105_n673) );
  AND2_X1 DP_mult_105_U505 ( .A1(DP_mult_105_n671), .A2(DP_mult_105_n480), 
        .ZN(DP_mult_105_n672) );
  AND2_X1 DP_mult_105_U504 ( .A1(DP_mult_105_n111), .A2(DP_mult_105_n93), .ZN(
        DP_mult_105_n671) );
  AND2_X1 DP_mult_105_U503 ( .A1(DP_mult_105_n111), .A2(DP_mult_105_n77), .ZN(
        DP_mult_105_n670) );
  AND2_X1 DP_mult_105_U502 ( .A1(DP_mult_105_n381), .A2(DP_mult_105_n386), 
        .ZN(DP_mult_105_n669) );
  OR2_X1 DP_mult_105_U501 ( .A1(DP_mult_105_n671), .A2(DP_mult_105_n480), .ZN(
        DP_mult_105_n668) );
  OR2_X1 DP_mult_105_U500 ( .A1(DP_mult_105_n283), .A2(DP_mult_105_n286), .ZN(
        DP_mult_105_n667) );
  OR2_X1 DP_mult_105_U499 ( .A1(DP_mult_105_n297), .A2(DP_mult_105_n302), .ZN(
        DP_mult_105_n666) );
  AND2_X1 DP_mult_105_U498 ( .A1(DP_mult_105_n403), .A2(DP_mult_105_n481), 
        .ZN(DP_mult_105_n665) );
  OR2_X1 DP_mult_105_U497 ( .A1(DP_mult_105_n281), .A2(DP_mult_105_n282), .ZN(
        DP_mult_105_n664) );
  OR2_X1 DP_mult_105_U496 ( .A1(DP_mult_105_n296), .A2(DP_mult_105_n291), .ZN(
        DP_mult_105_n663) );
  NOR2_X1 DP_mult_105_U495 ( .A1(DP_mult_105_n311), .A2(DP_mult_105_n318), 
        .ZN(DP_mult_105_n198) );
  OAI22_X1 DP_mult_105_U494 ( .A1(DP_mult_105_n585), .A2(DP_mult_105_n483), 
        .B1(DP_mult_105_n591), .B2(DP_mult_105_n482), .ZN(DP_mult_105_n278) );
  BUF_X1 DP_mult_105_U493 ( .A(DP_mult_105_n614), .Z(DP_mult_105_n590) );
  BUF_X1 DP_mult_105_U492 ( .A(DP_b_int[10]), .Z(DP_mult_105_n608) );
  BUF_X1 DP_mult_105_U491 ( .A(DP_b_int[4]), .Z(DP_mult_105_n605) );
  BUF_X1 DP_mult_105_U490 ( .A(DP_b_int[6]), .Z(DP_mult_105_n606) );
  AND2_X1 DP_mult_105_U489 ( .A1(DP_mult_105_n215), .A2(DP_mult_105_n726), 
        .ZN(DP_mult_105_n662) );
  XNOR2_X1 DP_mult_105_U488 ( .A(DP_mult_105_n662), .B(DP_mult_105_n216), .ZN(
        DP_w_b0_2_) );
  OR2_X2 DP_mult_105_U487 ( .A1(DP_mult_105_n287), .A2(DP_mult_105_n290), .ZN(
        DP_mult_105_n661) );
  HA_X1 DP_mult_105_U274 ( .A(DP_mult_105_n467), .B(DP_mult_105_n479), .CO(
        DP_mult_105_n396), .S(DP_mult_105_n397) );
  FA_X1 DP_mult_105_U273 ( .A(DP_mult_105_n466), .B(DP_mult_105_n478), .CI(
        DP_mult_105_n396), .CO(DP_mult_105_n394), .S(DP_mult_105_n395) );
  HA_X1 DP_mult_105_U272 ( .A(DP_mult_105_n454), .B(DP_mult_105_n477), .CO(
        DP_mult_105_n392), .S(DP_mult_105_n393) );
  FA_X1 DP_mult_105_U271 ( .A(DP_mult_105_n401), .B(DP_mult_105_n465), .CI(
        DP_mult_105_n393), .CO(DP_mult_105_n390), .S(DP_mult_105_n391) );
  FA_X1 DP_mult_105_U270 ( .A(DP_mult_105_n476), .B(DP_mult_105_n464), .CI(
        DP_mult_105_n453), .CO(DP_mult_105_n388), .S(DP_mult_105_n389) );
  FA_X1 DP_mult_105_U269 ( .A(DP_mult_105_n699), .B(DP_mult_105_n392), .CI(
        DP_mult_105_n389), .CO(DP_mult_105_n386), .S(DP_mult_105_n387) );
  HA_X1 DP_mult_105_U268 ( .A(DP_mult_105_n441), .B(DP_mult_105_n452), .CO(
        DP_mult_105_n384), .S(DP_mult_105_n385) );
  FA_X1 DP_mult_105_U267 ( .A(DP_mult_105_n463), .B(DP_mult_105_n475), .CI(
        DP_mult_105_n400), .CO(DP_mult_105_n382), .S(DP_mult_105_n383) );
  FA_X1 DP_mult_105_U266 ( .A(DP_mult_105_n388), .B(DP_mult_105_n385), .CI(
        DP_mult_105_n383), .CO(DP_mult_105_n380), .S(DP_mult_105_n381) );
  FA_X1 DP_mult_105_U265 ( .A(DP_mult_105_n462), .B(DP_mult_105_n440), .CI(
        DP_mult_105_n474), .CO(DP_mult_105_n378), .S(DP_mult_105_n379) );
  FA_X1 DP_mult_105_U264 ( .A(DP_mult_105_n384), .B(DP_mult_105_n451), .CI(
        DP_mult_105_n382), .CO(DP_mult_105_n376), .S(DP_mult_105_n377) );
  FA_X1 DP_mult_105_U263 ( .A(DP_mult_105_n379), .B(DP_mult_105_n700), .CI(
        DP_mult_105_n380), .CO(DP_mult_105_n374), .S(DP_mult_105_n375) );
  HA_X1 DP_mult_105_U262 ( .A(DP_mult_105_n428), .B(DP_mult_105_n439), .CO(
        DP_mult_105_n372), .S(DP_mult_105_n373) );
  FA_X1 DP_mult_105_U261 ( .A(DP_mult_105_n461), .B(DP_mult_105_n450), .CI(
        DP_mult_105_n399), .CO(DP_mult_105_n370), .S(DP_mult_105_n371) );
  FA_X1 DP_mult_105_U260 ( .A(DP_mult_105_n473), .B(DP_mult_105_n373), .CI(
        DP_mult_105_n378), .CO(DP_mult_105_n368), .S(DP_mult_105_n369) );
  FA_X1 DP_mult_105_U258 ( .A(DP_mult_105_n427), .B(DP_mult_105_n438), .CI(
        DP_mult_105_n472), .CO(DP_mult_105_n364), .S(DP_mult_105_n365) );
  FA_X1 DP_mult_105_U257 ( .A(DP_mult_105_n449), .B(DP_mult_105_n460), .CI(
        DP_mult_105_n372), .CO(DP_mult_105_n362), .S(DP_mult_105_n363) );
  HA_X1 DP_mult_105_U254 ( .A(DP_mult_105_n415), .B(DP_mult_105_n426), .CO(
        DP_mult_105_n356), .S(DP_mult_105_n357) );
  FA_X1 DP_mult_105_U252 ( .A(DP_mult_105_n437), .B(DP_mult_105_n459), .CI(
        DP_mult_105_n357), .CO(DP_mult_105_n352), .S(DP_mult_105_n353) );
  FA_X1 DP_mult_105_U250 ( .A(DP_mult_105_n353), .B(DP_mult_105_n360), .CI(
        DP_mult_105_n351), .CO(DP_mult_105_n348), .S(DP_mult_105_n349) );
  HA_X1 DP_mult_105_U249 ( .A(DP_mult_105_n414), .B(DP_mult_105_n425), .CO(
        DP_mult_105_n346), .S(DP_mult_105_n347) );
  FA_X1 DP_mult_105_U247 ( .A(DP_mult_105_n356), .B(DP_mult_105_n458), .CI(
        DP_mult_105_n347), .CO(DP_mult_105_n342), .S(DP_mult_105_n343) );
  FA_X1 DP_mult_105_U242 ( .A(DP_mult_105_n457), .B(DP_mult_105_n446), .CI(
        DP_mult_105_n435), .CO(DP_mult_105_n334), .S(DP_mult_105_n335) );
  FA_X1 DP_mult_105_U241 ( .A(DP_mult_105_n337), .B(DP_mult_105_n346), .CI(
        DP_mult_105_n469), .CO(DP_mult_105_n332), .S(DP_mult_105_n333) );
  FA_X1 DP_mult_105_U240 ( .A(DP_mult_105_n335), .B(DP_mult_105_n342), .CI(
        DP_mult_105_n344), .CO(DP_mult_105_n330), .S(DP_mult_105_n331) );
  FA_X1 DP_mult_105_U236 ( .A(DP_mult_105_n412), .B(DP_mult_105_n434), .CI(
        DP_mult_105_n336), .CO(DP_mult_105_n322), .S(DP_mult_105_n323) );
  FA_X1 DP_mult_105_U234 ( .A(DP_mult_105_n330), .B(DP_mult_105_n323), .CI(
        DP_mult_105_n321), .CO(DP_mult_105_n318), .S(DP_mult_105_n319) );
  FA_X1 DP_mult_105_U233 ( .A(DP_mult_105_n444), .B(DP_mult_105_n411), .CI(
        DP_mult_105_n748), .CO(DP_mult_105_n316), .S(DP_mult_105_n317) );
  FA_X1 DP_mult_105_U232 ( .A(DP_mult_105_n422), .B(DP_mult_105_n433), .CI(
        DP_mult_105_n456), .CO(DP_mult_105_n314), .S(DP_mult_105_n315) );
  FA_X1 DP_mult_105_U228 ( .A(DP_mult_105_n421), .B(DP_mult_105_n410), .CI(
        DP_mult_105_n309), .CO(DP_mult_105_n306), .S(DP_mult_105_n307) );
  FA_X1 DP_mult_105_U227 ( .A(DP_mult_105_n316), .B(DP_mult_105_n432), .CI(
        DP_mult_105_n307), .CO(DP_mult_105_n304), .S(DP_mult_105_n305) );
  FA_X1 DP_mult_105_U226 ( .A(DP_mult_105_n312), .B(DP_mult_105_n314), .CI(
        DP_mult_105_n305), .CO(DP_mult_105_n302), .S(DP_mult_105_n303) );
  FA_X1 DP_mult_105_U225 ( .A(DP_mult_105_n420), .B(DP_mult_105_n409), .CI(
        DP_mult_105_n308), .CO(DP_mult_105_n300), .S(DP_mult_105_n301) );
  FA_X1 DP_mult_105_U224 ( .A(DP_mult_105_n443), .B(DP_mult_105_n431), .CI(
        DP_mult_105_n306), .CO(DP_mult_105_n298), .S(DP_mult_105_n299) );
  FA_X1 DP_mult_105_U223 ( .A(DP_mult_105_n304), .B(DP_mult_105_n301), .CI(
        DP_mult_105_n299), .CO(DP_mult_105_n296), .S(DP_mult_105_n297) );
  FA_X1 DP_mult_105_U221 ( .A(DP_mult_105_n408), .B(DP_mult_105_n419), .CI(
        DP_mult_105_n295), .CO(DP_mult_105_n292), .S(DP_mult_105_n293) );
  FA_X1 DP_mult_105_U220 ( .A(DP_mult_105_n293), .B(DP_mult_105_n300), .CI(
        DP_mult_105_n298), .CO(DP_mult_105_n290), .S(DP_mult_105_n291) );
  FA_X1 DP_mult_105_U219 ( .A(DP_mult_105_n418), .B(DP_mult_105_n294), .CI(
        DP_mult_105_n407), .CO(DP_mult_105_n288), .S(DP_mult_105_n289) );
  FA_X1 DP_mult_105_U218 ( .A(DP_mult_105_n292), .B(DP_mult_105_n430), .CI(
        DP_mult_105_n289), .CO(DP_mult_105_n286), .S(DP_mult_105_n287) );
  FA_X1 DP_mult_105_U216 ( .A(DP_mult_105_n285), .B(DP_mult_105_n406), .CI(
        DP_mult_105_n288), .CO(DP_mult_105_n282), .S(DP_mult_105_n283) );
  FA_X1 DP_mult_105_U215 ( .A(DP_mult_105_n405), .B(DP_mult_105_n284), .CI(
        DP_mult_105_n417), .CO(DP_mult_105_n280), .S(DP_mult_105_n281) );
  INV_X1 CU_U14 ( .A(vOut), .ZN(CU_n5) );
  NAND2_X1 CU_U13 ( .A1(CU_n3), .A2(CU_n8), .ZN(CU_n6) );
  AOI21_X1 CU_U12 ( .B1(CU_n5), .B2(CU_n6), .A(CU_n1), .ZN(CU_nextState[1]) );
  NAND2_X1 CU_U11 ( .A1(CU_presentState_1_), .A2(CU_n8), .ZN(CU_n4) );
  INV_X1 CU_U10 ( .A(vIn), .ZN(CU_n1) );
  AOI21_X1 CU_U9 ( .B1(CU_presentState_2_), .B2(CU_presentState_0_), .A(vIn), 
        .ZN(CU_n12) );
  AOI21_X1 CU_U8 ( .B1(CU_n11), .B2(CU_n8), .A(CU_n12), .ZN(CU_n10) );
  OAI22_X1 CU_U7 ( .A1(CU_n1), .A2(CU_n4), .B1(CU_presentState_1_), .B2(CU_n10), .ZN(CU_nextState[0]) );
  NOR2_X1 CU_U6 ( .A1(CU_n3), .A2(CU_n9), .ZN(vOut) );
  NOR2_X1 CU_U5 ( .A1(vIn), .A2(CU_n4), .ZN(CU_N20) );
  INV_X1 CU_U4 ( .A(CU_n4), .ZN(reg_sw0_en_int) );
  XOR2_X1 CU_U16 ( .A(CU_presentState_1_), .B(CU_presentState_0_), .Z(CU_n3)
         );
  XOR2_X1 CU_U15 ( .A(CU_n8), .B(CU_presentState_0_), .Z(CU_n9) );
  NOR3_X2 CU_U3 ( .A1(CU_n3), .A2(CU_presentState_2_), .A3(CU_presentState_0_), 
        .ZN(regs_clr_int) );
  DFFR_X1 CU_presentState_reg_2_ ( .D(CU_N20), .CK(clk), .RN(rst_n), .Q(
        CU_presentState_2_), .QN(CU_n8) );
  DFFR_X1 CU_presentState_reg_1_ ( .D(CU_nextState[1]), .CK(clk), .RN(rst_n), 
        .Q(CU_presentState_1_) );
  DFFR_X1 CU_presentState_reg_0_ ( .D(CU_nextState[0]), .CK(clk), .RN(rst_n), 
        .Q(CU_presentState_0_), .QN(CU_n11) );
endmodule

