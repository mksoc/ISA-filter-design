
module iir_filter ( clk, rst_n, vIn, dIn, a, b, dOut, vOut );
  input [11:0] dIn;
  input [23:0] a;
  input [35:0] b;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   sw_regs_en_int, delayed_controls_0__1_, delayed_controls_1__0_,
         delayed_controls_1__1_, delayed_controls_2__0_, DP_n13, DP_n12,
         DP_n11, DP_n10, DP_n9, DP_n8, DP_n7, DP_n6, DP_n5, DP_n4, DP_n3,
         DP_n2, DP_n1, DP_fb_10_, DP_fb_11_, DP_fb_12_, DP_fb_13_, DP_fb_14_,
         DP_fb_15_, DP_fb_16_, DP_fb_17_, DP_fb_18_, DP_fb_19_, DP_fb_1_,
         DP_fb_20_, DP_fb_21_, DP_fb_22_, DP_fb_23_, DP_fb_2_, DP_fb_3_,
         DP_fb_4_, DP_fb_5_, DP_fb_6_, DP_fb_7_, DP_fb_8_, DP_fb_9_, DP_N123,
         DP_N124, DP_N125, DP_N126, DP_N127, DP_N128, DP_N129, DP_N130,
         DP_N131, DP_N132, DP_N133, DP_N134, DP_N135, DP_N136, DP_N137,
         DP_N138, DP_N139, DP_N140, DP_N141, DP_N142, DP_N143, DP_N144,
         DP_N145, DP_N100, DP_N101, DP_N102, DP_N103, DP_N104, DP_N105,
         DP_N106, DP_N107, DP_N108, DP_N109, DP_N110, DP_N111, DP_N112,
         DP_N113, DP_N114, DP_N115, DP_N116, DP_N117, DP_N118, DP_N119,
         DP_N120, DP_N121, DP_N99, DP_N75, DP_N76, DP_N77, DP_N78, DP_N79,
         DP_N80, DP_N81, DP_N82, DP_N83, DP_N84, DP_N85, DP_N86, DP_N87,
         DP_N88, DP_N89, DP_N90, DP_N91, DP_N92, DP_N93, DP_N94, DP_N95,
         DP_N96, DP_N97, DP_N51, DP_N52, DP_N53, DP_N54, DP_N55, DP_N56,
         DP_N57, DP_N58, DP_N59, DP_N60, DP_N61, DP_N62, DP_N63, DP_N64,
         DP_N65, DP_N66, DP_N67, DP_N68, DP_N69, DP_N70, DP_N71, DP_N72,
         DP_N73, DP_N10, DP_N11, DP_N12, DP_N13, DP_N14, DP_N15, DP_N16,
         DP_N17, DP_N18, DP_N19, DP_N20, DP_N21, DP_N22, DP_N23, DP_N24,
         DP_N25, DP_N37, DP_N38, DP_N39, DP_N4, DP_N40, DP_N41, DP_N42, DP_N43,
         DP_N44, DP_N45, DP_N46, DP_N47, DP_N49, DP_N5, DP_N6, DP_N7, DP_N8,
         DP_N9, DP_ff_0_, DP_ff_10_, DP_ff_11_, DP_ff_12_, DP_ff_13_,
         DP_ff_14_, DP_ff_15_, DP_ff_16_, DP_ff_17_, DP_ff_18_, DP_ff_19_,
         DP_ff_1_, DP_ff_20_, DP_ff_21_, DP_ff_22_, DP_ff_23_, DP_ff_2_,
         DP_ff_3_, DP_ff_4_, DP_ff_5_, DP_ff_6_, DP_ff_7_, DP_ff_8_, DP_ff_9_,
         DP_ff_part_0_, DP_ff_part_10_, DP_ff_part_11_, DP_ff_part_12_,
         DP_ff_part_13_, DP_ff_part_14_, DP_ff_part_15_, DP_ff_part_16_,
         DP_ff_part_17_, DP_ff_part_18_, DP_ff_part_19_, DP_ff_part_1_,
         DP_ff_part_20_, DP_ff_part_21_, DP_ff_part_22_, DP_ff_part_23_,
         DP_ff_part_2_, DP_ff_part_3_, DP_ff_part_4_, DP_ff_part_5_,
         DP_ff_part_6_, DP_ff_part_7_, DP_ff_part_8_, DP_ff_part_9_, DP_n66,
         DP_n65, DP_n64, DP_n63, DP_n62, DP_n61, DP_n60, DP_n59, DP_n58,
         DP_n57, DP_n56, DP_n55, DP_n54, DP_N148, DP_N146, DP_y_0_, DP_y_1_,
         DP_y_2_, DP_y_3_, DP_y_4_, DP_y_5_, DP_y_6_, DP_y_7_, DP_y_8_,
         DP_y_9_, DP_y_10_, DP_y_11_, DP_y_23, DP_sw1_0_, DP_sw1_1_, DP_sw1_2_,
         DP_sw1_3_, DP_sw1_4_, DP_sw1_5_, DP_sw1_6_, DP_sw1_7_, DP_sw1_8_,
         DP_sw1_9_, DP_sw1_10_, DP_sw1_11_, DP_sw1_12_, DP_sw1_13_, DP_sw1_14_,
         DP_sw1_15_, DP_sw1_16_, DP_sw1_17_, DP_sw1_18_, DP_sw1_19_,
         DP_sw1_20_, DP_sw1_21_, DP_sw1_22_, DP_sw1_23_, DP_sw0_0_, DP_sw0_1_,
         DP_sw0_2_, DP_sw0_3_, DP_sw0_4_, DP_sw0_5_, DP_sw0_6_, DP_sw0_7_,
         DP_sw0_8_, DP_sw0_9_, DP_sw0_10_, DP_sw0_11_, DP_sw0_12_, DP_sw0_13_,
         DP_sw0_14_, DP_sw0_15_, DP_sw0_16_, DP_sw0_17_, DP_sw0_18_,
         DP_sw0_19_, DP_sw0_20_, DP_sw0_21_, DP_sw0_22_, DP_sw0_23_, DP_w_0_,
         DP_w_1_, DP_w_2_, DP_w_3_, DP_w_4_, DP_w_5_, DP_w_6_, DP_w_7_,
         DP_w_8_, DP_w_9_, DP_w_10_, DP_w_11_, DP_w_12_, DP_w_13_, DP_w_14_,
         DP_w_15_, DP_w_16_, DP_w_17_, DP_w_18_, DP_w_19_, DP_w_20_, DP_w_21_,
         DP_w_22_, DP_w_23_, DP_b_int_2__0_, DP_b_int_2__1_, DP_b_int_2__2_,
         DP_b_int_2__3_, DP_b_int_2__4_, DP_b_int_2__5_, DP_b_int_2__6_,
         DP_b_int_2__7_, DP_b_int_2__8_, DP_b_int_2__9_, DP_b_int_2__10_,
         DP_b_int_2__11_, DP_b_int_1__0_, DP_b_int_1__1_, DP_b_int_1__2_,
         DP_b_int_1__3_, DP_b_int_1__4_, DP_b_int_1__5_, DP_b_int_1__6_,
         DP_b_int_1__7_, DP_b_int_1__8_, DP_b_int_1__9_, DP_b_int_1__10_,
         DP_b_int_1__11_, DP_b_int_0__0_, DP_b_int_0__1_, DP_b_int_0__2_,
         DP_b_int_0__3_, DP_b_int_0__4_, DP_b_int_0__5_, DP_b_int_0__6_,
         DP_b_int_0__7_, DP_b_int_0__8_, DP_b_int_0__9_, DP_b_int_0__10_,
         DP_b_int_0__11_, DP_a_int_1__1_, DP_a_int_1__2_, DP_a_int_1__3_,
         DP_a_int_1__4_, DP_a_int_1__5_, DP_a_int_1__6_, DP_a_int_1__7_,
         DP_a_int_1__8_, DP_a_int_1__9_, DP_a_int_1__10_, DP_a_int_1__11_,
         DP_x_0_, DP_x_1_, DP_x_2_, DP_x_3_, DP_x_4_, DP_x_5_, DP_x_6_,
         DP_x_7_, DP_x_8_, DP_x_9_, DP_x_10_, DP_x_11_, DP_reg_in_n39,
         DP_reg_in_n38, DP_reg_in_n37, DP_reg_in_n36, DP_reg_in_n35,
         DP_reg_in_n34, DP_reg_in_n33, DP_reg_in_n32, DP_reg_in_n31,
         DP_reg_in_n30, DP_reg_in_n29, DP_reg_in_n28, DP_reg_in_n27,
         DP_reg_in_n26, DP_reg_in_n25, DP_reg_in_n24, DP_reg_in_n23,
         DP_reg_in_n22, DP_reg_in_n21, DP_reg_in_n20, DP_reg_in_n19,
         DP_reg_in_n18, DP_reg_in_n17, DP_reg_in_n16, DP_reg_in_n15,
         DP_reg_in_n14, DP_reg_in_n13, DP_reg_in_n12, DP_reg_in_n11,
         DP_reg_in_n10, DP_reg_in_n9, DP_reg_in_n8, DP_reg_in_n7, DP_reg_in_n6,
         DP_reg_in_n5, DP_reg_in_n4, DP_reg_in_n3, DP_reg_in_n2, DP_reg_in_n1,
         DP_reg_a_i_1_n75, DP_reg_a_i_1_n74, DP_reg_a_i_1_n73,
         DP_reg_a_i_1_n72, DP_reg_a_i_1_n71, DP_reg_a_i_1_n70,
         DP_reg_a_i_1_n69, DP_reg_a_i_1_n68, DP_reg_a_i_1_n67,
         DP_reg_a_i_1_n66, DP_reg_a_i_1_n65, DP_reg_a_i_1_n64,
         DP_reg_a_i_1_n63, DP_reg_a_i_1_n62, DP_reg_a_i_1_n61,
         DP_reg_a_i_1_n60, DP_reg_a_i_1_n59, DP_reg_a_i_1_n58,
         DP_reg_a_i_1_n57, DP_reg_a_i_1_n56, DP_reg_a_i_1_n55,
         DP_reg_a_i_1_n54, DP_reg_a_i_1_n53, DP_reg_a_i_1_n52,
         DP_reg_a_i_1_n51, DP_reg_a_i_1_n50, DP_reg_a_i_1_n49,
         DP_reg_a_i_1_n48, DP_reg_a_i_1_n47, DP_reg_a_i_1_n46,
         DP_reg_a_i_1_n45, DP_reg_a_i_1_n44, DP_reg_a_i_1_n43,
         DP_reg_a_i_1_n42, DP_reg_a_i_1_n41, DP_reg_a_i_1_n40,
         DP_reg_a_i_1_n39, DP_reg_a_i_1_n38, DP_reg_a_i_1_n37,
         DP_reg_a_i_2_n75, DP_reg_a_i_2_n74, DP_reg_a_i_2_n73,
         DP_reg_a_i_2_n72, DP_reg_a_i_2_n71, DP_reg_a_i_2_n70,
         DP_reg_a_i_2_n69, DP_reg_a_i_2_n68, DP_reg_a_i_2_n67,
         DP_reg_a_i_2_n66, DP_reg_a_i_2_n65, DP_reg_a_i_2_n64,
         DP_reg_a_i_2_n63, DP_reg_a_i_2_n62, DP_reg_a_i_2_n61,
         DP_reg_a_i_2_n60, DP_reg_a_i_2_n59, DP_reg_a_i_2_n58,
         DP_reg_a_i_2_n57, DP_reg_a_i_2_n56, DP_reg_a_i_2_n55,
         DP_reg_a_i_2_n54, DP_reg_a_i_2_n53, DP_reg_a_i_2_n52,
         DP_reg_a_i_2_n51, DP_reg_a_i_2_n50, DP_reg_a_i_2_n49,
         DP_reg_a_i_2_n48, DP_reg_a_i_2_n47, DP_reg_a_i_2_n46,
         DP_reg_a_i_2_n45, DP_reg_a_i_2_n44, DP_reg_a_i_2_n43,
         DP_reg_a_i_2_n42, DP_reg_a_i_2_n41, DP_reg_a_i_2_n40,
         DP_reg_a_i_2_n39, DP_reg_a_i_2_n38, DP_reg_a_i_2_n37,
         DP_reg_b_i_0_n75, DP_reg_b_i_0_n74, DP_reg_b_i_0_n73,
         DP_reg_b_i_0_n72, DP_reg_b_i_0_n71, DP_reg_b_i_0_n70,
         DP_reg_b_i_0_n69, DP_reg_b_i_0_n68, DP_reg_b_i_0_n67,
         DP_reg_b_i_0_n66, DP_reg_b_i_0_n65, DP_reg_b_i_0_n64,
         DP_reg_b_i_0_n63, DP_reg_b_i_0_n62, DP_reg_b_i_0_n61,
         DP_reg_b_i_0_n60, DP_reg_b_i_0_n59, DP_reg_b_i_0_n58,
         DP_reg_b_i_0_n57, DP_reg_b_i_0_n56, DP_reg_b_i_0_n55,
         DP_reg_b_i_0_n54, DP_reg_b_i_0_n53, DP_reg_b_i_0_n52,
         DP_reg_b_i_0_n51, DP_reg_b_i_0_n50, DP_reg_b_i_0_n49,
         DP_reg_b_i_0_n48, DP_reg_b_i_0_n47, DP_reg_b_i_0_n46,
         DP_reg_b_i_0_n45, DP_reg_b_i_0_n44, DP_reg_b_i_0_n43,
         DP_reg_b_i_0_n42, DP_reg_b_i_0_n41, DP_reg_b_i_0_n40,
         DP_reg_b_i_0_n39, DP_reg_b_i_0_n38, DP_reg_b_i_0_n37,
         DP_reg_b_i_1_n75, DP_reg_b_i_1_n74, DP_reg_b_i_1_n73,
         DP_reg_b_i_1_n72, DP_reg_b_i_1_n71, DP_reg_b_i_1_n70,
         DP_reg_b_i_1_n69, DP_reg_b_i_1_n68, DP_reg_b_i_1_n67,
         DP_reg_b_i_1_n66, DP_reg_b_i_1_n65, DP_reg_b_i_1_n64,
         DP_reg_b_i_1_n63, DP_reg_b_i_1_n62, DP_reg_b_i_1_n61,
         DP_reg_b_i_1_n60, DP_reg_b_i_1_n59, DP_reg_b_i_1_n58,
         DP_reg_b_i_1_n57, DP_reg_b_i_1_n56, DP_reg_b_i_1_n55,
         DP_reg_b_i_1_n54, DP_reg_b_i_1_n53, DP_reg_b_i_1_n52,
         DP_reg_b_i_1_n51, DP_reg_b_i_1_n50, DP_reg_b_i_1_n49,
         DP_reg_b_i_1_n48, DP_reg_b_i_1_n47, DP_reg_b_i_1_n46,
         DP_reg_b_i_1_n45, DP_reg_b_i_1_n44, DP_reg_b_i_1_n43,
         DP_reg_b_i_1_n42, DP_reg_b_i_1_n41, DP_reg_b_i_1_n40,
         DP_reg_b_i_1_n39, DP_reg_b_i_1_n38, DP_reg_b_i_1_n37,
         DP_reg_b_i_2_n75, DP_reg_b_i_2_n74, DP_reg_b_i_2_n73,
         DP_reg_b_i_2_n72, DP_reg_b_i_2_n71, DP_reg_b_i_2_n70,
         DP_reg_b_i_2_n69, DP_reg_b_i_2_n68, DP_reg_b_i_2_n67,
         DP_reg_b_i_2_n66, DP_reg_b_i_2_n65, DP_reg_b_i_2_n64,
         DP_reg_b_i_2_n63, DP_reg_b_i_2_n62, DP_reg_b_i_2_n61,
         DP_reg_b_i_2_n60, DP_reg_b_i_2_n59, DP_reg_b_i_2_n58,
         DP_reg_b_i_2_n57, DP_reg_b_i_2_n56, DP_reg_b_i_2_n55,
         DP_reg_b_i_2_n54, DP_reg_b_i_2_n53, DP_reg_b_i_2_n52,
         DP_reg_b_i_2_n51, DP_reg_b_i_2_n50, DP_reg_b_i_2_n49,
         DP_reg_b_i_2_n48, DP_reg_b_i_2_n47, DP_reg_b_i_2_n46,
         DP_reg_b_i_2_n45, DP_reg_b_i_2_n44, DP_reg_b_i_2_n43,
         DP_reg_b_i_2_n42, DP_reg_b_i_2_n41, DP_reg_b_i_2_n40,
         DP_reg_b_i_2_n39, DP_reg_b_i_2_n38, DP_reg_b_i_2_n37, DP_reg_sw0_n80,
         DP_reg_sw0_n79, DP_reg_sw0_n78, DP_reg_sw0_n77, DP_reg_sw0_n76,
         DP_reg_sw0_n75, DP_reg_sw0_n74, DP_reg_sw0_n73, DP_reg_sw0_n72,
         DP_reg_sw0_n71, DP_reg_sw0_n70, DP_reg_sw0_n69, DP_reg_sw0_n68,
         DP_reg_sw0_n67, DP_reg_sw0_n66, DP_reg_sw0_n65, DP_reg_sw0_n64,
         DP_reg_sw0_n63, DP_reg_sw0_n62, DP_reg_sw0_n61, DP_reg_sw0_n60,
         DP_reg_sw0_n59, DP_reg_sw0_n58, DP_reg_sw0_n57, DP_reg_sw0_n56,
         DP_reg_sw0_n55, DP_reg_sw0_n54, DP_reg_sw0_n53, DP_reg_sw0_n52,
         DP_reg_sw0_n51, DP_reg_sw0_n50, DP_reg_sw0_n49, DP_reg_sw0_n48,
         DP_reg_sw0_n47, DP_reg_sw0_n46, DP_reg_sw0_n45, DP_reg_sw0_n44,
         DP_reg_sw0_n43, DP_reg_sw0_n42, DP_reg_sw0_n41, DP_reg_sw0_n40,
         DP_reg_sw0_n39, DP_reg_sw0_n38, DP_reg_sw0_n37, DP_reg_sw0_n36,
         DP_reg_sw0_n35, DP_reg_sw0_n34, DP_reg_sw0_n33, DP_reg_sw0_n32,
         DP_reg_sw0_n31, DP_reg_sw0_n30, DP_reg_sw0_n29, DP_reg_sw0_n28,
         DP_reg_sw0_n27, DP_reg_sw0_n26, DP_reg_sw0_n25, DP_reg_sw0_n24,
         DP_reg_sw0_n23, DP_reg_sw0_n22, DP_reg_sw0_n21, DP_reg_sw0_n20,
         DP_reg_sw0_n19, DP_reg_sw0_n18, DP_reg_sw0_n17, DP_reg_sw0_n16,
         DP_reg_sw0_n15, DP_reg_sw0_n14, DP_reg_sw0_n13, DP_reg_sw0_n12,
         DP_reg_sw0_n11, DP_reg_sw0_n10, DP_reg_sw0_n9, DP_reg_sw0_n8,
         DP_reg_sw0_n7, DP_reg_sw0_n6, DP_reg_sw0_n5, DP_reg_sw0_n4,
         DP_reg_sw0_n3, DP_reg_sw0_n2, DP_reg_sw0_n1, DP_reg_sw1_n152,
         DP_reg_sw1_n151, DP_reg_sw1_n150, DP_reg_sw1_n149, DP_reg_sw1_n148,
         DP_reg_sw1_n147, DP_reg_sw1_n146, DP_reg_sw1_n145, DP_reg_sw1_n144,
         DP_reg_sw1_n143, DP_reg_sw1_n142, DP_reg_sw1_n141, DP_reg_sw1_n140,
         DP_reg_sw1_n139, DP_reg_sw1_n138, DP_reg_sw1_n137, DP_reg_sw1_n136,
         DP_reg_sw1_n135, DP_reg_sw1_n134, DP_reg_sw1_n133, DP_reg_sw1_n132,
         DP_reg_sw1_n131, DP_reg_sw1_n130, DP_reg_sw1_n129, DP_reg_sw1_n128,
         DP_reg_sw1_n127, DP_reg_sw1_n126, DP_reg_sw1_n125, DP_reg_sw1_n124,
         DP_reg_sw1_n123, DP_reg_sw1_n122, DP_reg_sw1_n121, DP_reg_sw1_n120,
         DP_reg_sw1_n119, DP_reg_sw1_n118, DP_reg_sw1_n117, DP_reg_sw1_n116,
         DP_reg_sw1_n115, DP_reg_sw1_n114, DP_reg_sw1_n113, DP_reg_sw1_n112,
         DP_reg_sw1_n111, DP_reg_sw1_n110, DP_reg_sw1_n109, DP_reg_sw1_n108,
         DP_reg_sw1_n107, DP_reg_sw1_n106, DP_reg_sw1_n105, DP_reg_sw1_n104,
         DP_reg_sw1_n103, DP_reg_sw1_n102, DP_reg_sw1_n101, DP_reg_sw1_n100,
         DP_reg_sw1_n99, DP_reg_sw1_n98, DP_reg_sw1_n97, DP_reg_sw1_n96,
         DP_reg_sw1_n95, DP_reg_sw1_n94, DP_reg_sw1_n93, DP_reg_sw1_n92,
         DP_reg_sw1_n91, DP_reg_sw1_n90, DP_reg_sw1_n89, DP_reg_sw1_n88,
         DP_reg_sw1_n87, DP_reg_sw1_n86, DP_reg_sw1_n85, DP_reg_sw1_n84,
         DP_reg_sw1_n83, DP_reg_sw1_n82, DP_reg_sw1_n81, DP_reg_sw1_n80,
         DP_reg_sw1_n79, DP_reg_sw1_n78, DP_reg_sw1_n77, DP_reg_sw1_n76,
         DP_reg_sw1_n75, DP_reg_sw1_n74, DP_reg_sw1_n73, DP_reg_sw2_n152,
         DP_reg_sw2_n151, DP_reg_sw2_n150, DP_reg_sw2_n149, DP_reg_sw2_n148,
         DP_reg_sw2_n147, DP_reg_sw2_n146, DP_reg_sw2_n145, DP_reg_sw2_n144,
         DP_reg_sw2_n143, DP_reg_sw2_n142, DP_reg_sw2_n141, DP_reg_sw2_n140,
         DP_reg_sw2_n139, DP_reg_sw2_n138, DP_reg_sw2_n137, DP_reg_sw2_n136,
         DP_reg_sw2_n135, DP_reg_sw2_n134, DP_reg_sw2_n133, DP_reg_sw2_n132,
         DP_reg_sw2_n131, DP_reg_sw2_n130, DP_reg_sw2_n129, DP_reg_sw2_n128,
         DP_reg_sw2_n127, DP_reg_sw2_n126, DP_reg_sw2_n125, DP_reg_sw2_n124,
         DP_reg_sw2_n123, DP_reg_sw2_n122, DP_reg_sw2_n121, DP_reg_sw2_n120,
         DP_reg_sw2_n119, DP_reg_sw2_n118, DP_reg_sw2_n117, DP_reg_sw2_n116,
         DP_reg_sw2_n115, DP_reg_sw2_n114, DP_reg_sw2_n113, DP_reg_sw2_n112,
         DP_reg_sw2_n111, DP_reg_sw2_n110, DP_reg_sw2_n109, DP_reg_sw2_n108,
         DP_reg_sw2_n107, DP_reg_sw2_n106, DP_reg_sw2_n105, DP_reg_sw2_n104,
         DP_reg_sw2_n103, DP_reg_sw2_n102, DP_reg_sw2_n101, DP_reg_sw2_n100,
         DP_reg_sw2_n99, DP_reg_sw2_n98, DP_reg_sw2_n97, DP_reg_sw2_n96,
         DP_reg_sw2_n95, DP_reg_sw2_n94, DP_reg_sw2_n93, DP_reg_sw2_n92,
         DP_reg_sw2_n91, DP_reg_sw2_n90, DP_reg_sw2_n89, DP_reg_sw2_n88,
         DP_reg_sw2_n87, DP_reg_sw2_n86, DP_reg_sw2_n85, DP_reg_sw2_n84,
         DP_reg_sw2_n83, DP_reg_sw2_n82, DP_reg_sw2_n81, DP_reg_sw2_n80,
         DP_reg_sw2_n79, DP_reg_sw2_n78, DP_reg_sw2_n77, DP_reg_sw2_n76,
         DP_reg_sw2_n75, DP_reg_sw2_n74, DP_reg_sw2_n73, DP_reg_ret0_n146,
         DP_reg_ret0_n145, DP_reg_ret0_n144, DP_reg_ret0_n143,
         DP_reg_ret0_n142, DP_reg_ret0_n141, DP_reg_ret0_n140,
         DP_reg_ret0_n139, DP_reg_ret0_n138, DP_reg_ret0_n137,
         DP_reg_ret0_n136, DP_reg_ret0_n135, DP_reg_ret0_n134,
         DP_reg_ret0_n133, DP_reg_ret0_n132, DP_reg_ret0_n131,
         DP_reg_ret0_n130, DP_reg_ret0_n129, DP_reg_ret0_n128,
         DP_reg_ret0_n127, DP_reg_ret0_n126, DP_reg_ret0_n125,
         DP_reg_ret0_n124, DP_reg_ret0_n123, DP_reg_ret0_n122,
         DP_reg_ret0_n121, DP_reg_ret0_n120, DP_reg_ret0_n119,
         DP_reg_ret0_n118, DP_reg_ret0_n117, DP_reg_ret0_n116,
         DP_reg_ret0_n115, DP_reg_ret0_n114, DP_reg_ret0_n113,
         DP_reg_ret0_n112, DP_reg_ret0_n111, DP_reg_ret0_n110,
         DP_reg_ret0_n109, DP_reg_ret0_n108, DP_reg_ret0_n107,
         DP_reg_ret0_n106, DP_reg_ret0_n105, DP_reg_ret0_n104,
         DP_reg_ret0_n103, DP_reg_ret0_n102, DP_reg_ret0_n101,
         DP_reg_ret0_n100, DP_reg_ret0_n99, DP_reg_ret0_n98, DP_reg_ret0_n97,
         DP_reg_ret0_n96, DP_reg_ret0_n95, DP_reg_ret0_n94, DP_reg_ret0_n93,
         DP_reg_ret0_n92, DP_reg_ret0_n91, DP_reg_ret0_n90, DP_reg_ret0_n89,
         DP_reg_ret0_n88, DP_reg_ret0_n87, DP_reg_ret0_n86, DP_reg_ret0_n85,
         DP_reg_ret0_n84, DP_reg_ret0_n83, DP_reg_ret0_n82, DP_reg_ret0_n81,
         DP_reg_ret0_n80, DP_reg_ret0_n79, DP_reg_ret0_n78, DP_reg_ret0_n77,
         DP_reg_ret0_n76, DP_reg_ret0_n75, DP_reg_ret0_n74, DP_reg_ret0_n73,
         DP_reg_ret1_n146, DP_reg_ret1_n145, DP_reg_ret1_n144,
         DP_reg_ret1_n143, DP_reg_ret1_n142, DP_reg_ret1_n141,
         DP_reg_ret1_n140, DP_reg_ret1_n139, DP_reg_ret1_n138,
         DP_reg_ret1_n137, DP_reg_ret1_n136, DP_reg_ret1_n135,
         DP_reg_ret1_n134, DP_reg_ret1_n133, DP_reg_ret1_n132,
         DP_reg_ret1_n131, DP_reg_ret1_n130, DP_reg_ret1_n129,
         DP_reg_ret1_n128, DP_reg_ret1_n127, DP_reg_ret1_n126,
         DP_reg_ret1_n125, DP_reg_ret1_n124, DP_reg_ret1_n123,
         DP_reg_ret1_n122, DP_reg_ret1_n121, DP_reg_ret1_n120,
         DP_reg_ret1_n119, DP_reg_ret1_n118, DP_reg_ret1_n117,
         DP_reg_ret1_n116, DP_reg_ret1_n115, DP_reg_ret1_n114,
         DP_reg_ret1_n113, DP_reg_ret1_n112, DP_reg_ret1_n111,
         DP_reg_ret1_n110, DP_reg_ret1_n109, DP_reg_ret1_n108,
         DP_reg_ret1_n107, DP_reg_ret1_n106, DP_reg_ret1_n105,
         DP_reg_ret1_n104, DP_reg_ret1_n103, DP_reg_ret1_n102,
         DP_reg_ret1_n101, DP_reg_ret1_n100, DP_reg_ret1_n99, DP_reg_ret1_n98,
         DP_reg_ret1_n97, DP_reg_ret1_n96, DP_reg_ret1_n95, DP_reg_ret1_n94,
         DP_reg_ret1_n93, DP_reg_ret1_n92, DP_reg_ret1_n91, DP_reg_ret1_n90,
         DP_reg_ret1_n89, DP_reg_ret1_n88, DP_reg_ret1_n87, DP_reg_ret1_n86,
         DP_reg_ret1_n85, DP_reg_ret1_n84, DP_reg_ret1_n83, DP_reg_ret1_n82,
         DP_reg_ret1_n81, DP_reg_ret1_n80, DP_reg_ret1_n79, DP_reg_ret1_n78,
         DP_reg_ret1_n77, DP_reg_ret1_n76, DP_reg_ret1_n75, DP_reg_ret1_n74,
         DP_reg_ret1_n73, DP_reg_pipe00_n146, DP_reg_pipe00_n145,
         DP_reg_pipe00_n144, DP_reg_pipe00_n143, DP_reg_pipe00_n142,
         DP_reg_pipe00_n141, DP_reg_pipe00_n140, DP_reg_pipe00_n139,
         DP_reg_pipe00_n138, DP_reg_pipe00_n137, DP_reg_pipe00_n136,
         DP_reg_pipe00_n135, DP_reg_pipe00_n134, DP_reg_pipe00_n133,
         DP_reg_pipe00_n132, DP_reg_pipe00_n131, DP_reg_pipe00_n130,
         DP_reg_pipe00_n129, DP_reg_pipe00_n128, DP_reg_pipe00_n127,
         DP_reg_pipe00_n126, DP_reg_pipe00_n125, DP_reg_pipe00_n124,
         DP_reg_pipe00_n123, DP_reg_pipe00_n122, DP_reg_pipe00_n121,
         DP_reg_pipe00_n120, DP_reg_pipe00_n119, DP_reg_pipe00_n118,
         DP_reg_pipe00_n117, DP_reg_pipe00_n116, DP_reg_pipe00_n115,
         DP_reg_pipe00_n114, DP_reg_pipe00_n113, DP_reg_pipe00_n112,
         DP_reg_pipe00_n111, DP_reg_pipe00_n110, DP_reg_pipe00_n109,
         DP_reg_pipe00_n108, DP_reg_pipe00_n107, DP_reg_pipe00_n106,
         DP_reg_pipe00_n105, DP_reg_pipe00_n104, DP_reg_pipe00_n103,
         DP_reg_pipe00_n102, DP_reg_pipe00_n101, DP_reg_pipe00_n100,
         DP_reg_pipe00_n99, DP_reg_pipe00_n98, DP_reg_pipe00_n97,
         DP_reg_pipe00_n96, DP_reg_pipe00_n95, DP_reg_pipe00_n94,
         DP_reg_pipe00_n93, DP_reg_pipe00_n92, DP_reg_pipe00_n91,
         DP_reg_pipe00_n90, DP_reg_pipe00_n89, DP_reg_pipe00_n88,
         DP_reg_pipe00_n87, DP_reg_pipe00_n86, DP_reg_pipe00_n85,
         DP_reg_pipe00_n84, DP_reg_pipe00_n83, DP_reg_pipe00_n82,
         DP_reg_pipe00_n81, DP_reg_pipe00_n80, DP_reg_pipe00_n79,
         DP_reg_pipe00_n78, DP_reg_pipe00_n77, DP_reg_pipe00_n76,
         DP_reg_pipe00_n75, DP_reg_pipe00_n74, DP_reg_pipe00_n73,
         DP_reg_pipe01_n146, DP_reg_pipe01_n145, DP_reg_pipe01_n144,
         DP_reg_pipe01_n143, DP_reg_pipe01_n142, DP_reg_pipe01_n141,
         DP_reg_pipe01_n140, DP_reg_pipe01_n139, DP_reg_pipe01_n138,
         DP_reg_pipe01_n137, DP_reg_pipe01_n136, DP_reg_pipe01_n135,
         DP_reg_pipe01_n134, DP_reg_pipe01_n133, DP_reg_pipe01_n132,
         DP_reg_pipe01_n131, DP_reg_pipe01_n130, DP_reg_pipe01_n129,
         DP_reg_pipe01_n128, DP_reg_pipe01_n127, DP_reg_pipe01_n126,
         DP_reg_pipe01_n125, DP_reg_pipe01_n124, DP_reg_pipe01_n123,
         DP_reg_pipe01_n122, DP_reg_pipe01_n121, DP_reg_pipe01_n120,
         DP_reg_pipe01_n119, DP_reg_pipe01_n118, DP_reg_pipe01_n117,
         DP_reg_pipe01_n116, DP_reg_pipe01_n115, DP_reg_pipe01_n114,
         DP_reg_pipe01_n113, DP_reg_pipe01_n112, DP_reg_pipe01_n111,
         DP_reg_pipe01_n110, DP_reg_pipe01_n109, DP_reg_pipe01_n108,
         DP_reg_pipe01_n107, DP_reg_pipe01_n106, DP_reg_pipe01_n105,
         DP_reg_pipe01_n104, DP_reg_pipe01_n103, DP_reg_pipe01_n102,
         DP_reg_pipe01_n101, DP_reg_pipe01_n100, DP_reg_pipe01_n99,
         DP_reg_pipe01_n98, DP_reg_pipe01_n97, DP_reg_pipe01_n96,
         DP_reg_pipe01_n95, DP_reg_pipe01_n94, DP_reg_pipe01_n93,
         DP_reg_pipe01_n92, DP_reg_pipe01_n91, DP_reg_pipe01_n90,
         DP_reg_pipe01_n89, DP_reg_pipe01_n88, DP_reg_pipe01_n87,
         DP_reg_pipe01_n86, DP_reg_pipe01_n85, DP_reg_pipe01_n84,
         DP_reg_pipe01_n83, DP_reg_pipe01_n82, DP_reg_pipe01_n81,
         DP_reg_pipe01_n80, DP_reg_pipe01_n79, DP_reg_pipe01_n78,
         DP_reg_pipe01_n77, DP_reg_pipe01_n76, DP_reg_pipe01_n75,
         DP_reg_pipe01_n74, DP_reg_pipe01_n73, DP_reg_pipe02_n146,
         DP_reg_pipe02_n145, DP_reg_pipe02_n144, DP_reg_pipe02_n143,
         DP_reg_pipe02_n142, DP_reg_pipe02_n141, DP_reg_pipe02_n140,
         DP_reg_pipe02_n139, DP_reg_pipe02_n138, DP_reg_pipe02_n137,
         DP_reg_pipe02_n136, DP_reg_pipe02_n135, DP_reg_pipe02_n134,
         DP_reg_pipe02_n133, DP_reg_pipe02_n132, DP_reg_pipe02_n131,
         DP_reg_pipe02_n130, DP_reg_pipe02_n129, DP_reg_pipe02_n128,
         DP_reg_pipe02_n127, DP_reg_pipe02_n126, DP_reg_pipe02_n125,
         DP_reg_pipe02_n124, DP_reg_pipe02_n123, DP_reg_pipe02_n122,
         DP_reg_pipe02_n121, DP_reg_pipe02_n120, DP_reg_pipe02_n119,
         DP_reg_pipe02_n118, DP_reg_pipe02_n117, DP_reg_pipe02_n116,
         DP_reg_pipe02_n115, DP_reg_pipe02_n114, DP_reg_pipe02_n113,
         DP_reg_pipe02_n112, DP_reg_pipe02_n111, DP_reg_pipe02_n110,
         DP_reg_pipe02_n109, DP_reg_pipe02_n108, DP_reg_pipe02_n107,
         DP_reg_pipe02_n106, DP_reg_pipe02_n105, DP_reg_pipe02_n104,
         DP_reg_pipe02_n103, DP_reg_pipe02_n102, DP_reg_pipe02_n101,
         DP_reg_pipe02_n100, DP_reg_pipe02_n99, DP_reg_pipe02_n98,
         DP_reg_pipe02_n97, DP_reg_pipe02_n96, DP_reg_pipe02_n95,
         DP_reg_pipe02_n94, DP_reg_pipe02_n93, DP_reg_pipe02_n92,
         DP_reg_pipe02_n91, DP_reg_pipe02_n90, DP_reg_pipe02_n89,
         DP_reg_pipe02_n88, DP_reg_pipe02_n87, DP_reg_pipe02_n86,
         DP_reg_pipe02_n85, DP_reg_pipe02_n84, DP_reg_pipe02_n83,
         DP_reg_pipe02_n82, DP_reg_pipe02_n81, DP_reg_pipe02_n80,
         DP_reg_pipe02_n79, DP_reg_pipe02_n78, DP_reg_pipe02_n77,
         DP_reg_pipe02_n76, DP_reg_pipe02_n75, DP_reg_pipe02_n74,
         DP_reg_pipe02_n73, DP_reg_pipe03_n146, DP_reg_pipe03_n145,
         DP_reg_pipe03_n144, DP_reg_pipe03_n143, DP_reg_pipe03_n142,
         DP_reg_pipe03_n141, DP_reg_pipe03_n140, DP_reg_pipe03_n139,
         DP_reg_pipe03_n138, DP_reg_pipe03_n137, DP_reg_pipe03_n136,
         DP_reg_pipe03_n135, DP_reg_pipe03_n134, DP_reg_pipe03_n133,
         DP_reg_pipe03_n132, DP_reg_pipe03_n131, DP_reg_pipe03_n130,
         DP_reg_pipe03_n129, DP_reg_pipe03_n128, DP_reg_pipe03_n127,
         DP_reg_pipe03_n126, DP_reg_pipe03_n125, DP_reg_pipe03_n124,
         DP_reg_pipe03_n123, DP_reg_pipe03_n122, DP_reg_pipe03_n121,
         DP_reg_pipe03_n120, DP_reg_pipe03_n119, DP_reg_pipe03_n118,
         DP_reg_pipe03_n117, DP_reg_pipe03_n116, DP_reg_pipe03_n115,
         DP_reg_pipe03_n114, DP_reg_pipe03_n113, DP_reg_pipe03_n112,
         DP_reg_pipe03_n111, DP_reg_pipe03_n110, DP_reg_pipe03_n109,
         DP_reg_pipe03_n108, DP_reg_pipe03_n107, DP_reg_pipe03_n106,
         DP_reg_pipe03_n105, DP_reg_pipe03_n104, DP_reg_pipe03_n103,
         DP_reg_pipe03_n102, DP_reg_pipe03_n101, DP_reg_pipe03_n100,
         DP_reg_pipe03_n99, DP_reg_pipe03_n98, DP_reg_pipe03_n97,
         DP_reg_pipe03_n96, DP_reg_pipe03_n95, DP_reg_pipe03_n94,
         DP_reg_pipe03_n93, DP_reg_pipe03_n92, DP_reg_pipe03_n91,
         DP_reg_pipe03_n90, DP_reg_pipe03_n89, DP_reg_pipe03_n88,
         DP_reg_pipe03_n87, DP_reg_pipe03_n86, DP_reg_pipe03_n85,
         DP_reg_pipe03_n84, DP_reg_pipe03_n83, DP_reg_pipe03_n82,
         DP_reg_pipe03_n81, DP_reg_pipe03_n80, DP_reg_pipe03_n79,
         DP_reg_pipe03_n78, DP_reg_pipe03_n77, DP_reg_pipe03_n76,
         DP_reg_pipe03_n75, DP_reg_pipe03_n74, DP_reg_pipe03_n73,
         DP_reg_pipe10_n146, DP_reg_pipe10_n145, DP_reg_pipe10_n144,
         DP_reg_pipe10_n143, DP_reg_pipe10_n142, DP_reg_pipe10_n141,
         DP_reg_pipe10_n140, DP_reg_pipe10_n139, DP_reg_pipe10_n138,
         DP_reg_pipe10_n137, DP_reg_pipe10_n136, DP_reg_pipe10_n135,
         DP_reg_pipe10_n134, DP_reg_pipe10_n133, DP_reg_pipe10_n132,
         DP_reg_pipe10_n131, DP_reg_pipe10_n130, DP_reg_pipe10_n129,
         DP_reg_pipe10_n128, DP_reg_pipe10_n127, DP_reg_pipe10_n126,
         DP_reg_pipe10_n125, DP_reg_pipe10_n124, DP_reg_pipe10_n123,
         DP_reg_pipe10_n122, DP_reg_pipe10_n121, DP_reg_pipe10_n120,
         DP_reg_pipe10_n119, DP_reg_pipe10_n118, DP_reg_pipe10_n117,
         DP_reg_pipe10_n116, DP_reg_pipe10_n115, DP_reg_pipe10_n114,
         DP_reg_pipe10_n113, DP_reg_pipe10_n112, DP_reg_pipe10_n111,
         DP_reg_pipe10_n110, DP_reg_pipe10_n109, DP_reg_pipe10_n108,
         DP_reg_pipe10_n107, DP_reg_pipe10_n106, DP_reg_pipe10_n105,
         DP_reg_pipe10_n104, DP_reg_pipe10_n103, DP_reg_pipe10_n102,
         DP_reg_pipe10_n101, DP_reg_pipe10_n100, DP_reg_pipe10_n99,
         DP_reg_pipe10_n98, DP_reg_pipe10_n97, DP_reg_pipe10_n96,
         DP_reg_pipe10_n95, DP_reg_pipe10_n94, DP_reg_pipe10_n93,
         DP_reg_pipe10_n92, DP_reg_pipe10_n91, DP_reg_pipe10_n90,
         DP_reg_pipe10_n89, DP_reg_pipe10_n88, DP_reg_pipe10_n87,
         DP_reg_pipe10_n86, DP_reg_pipe10_n85, DP_reg_pipe10_n84,
         DP_reg_pipe10_n83, DP_reg_pipe10_n82, DP_reg_pipe10_n81,
         DP_reg_pipe10_n80, DP_reg_pipe10_n79, DP_reg_pipe10_n78,
         DP_reg_pipe10_n77, DP_reg_pipe10_n76, DP_reg_pipe10_n75,
         DP_reg_pipe10_n74, DP_reg_pipe10_n73, DP_reg_pipe11_n146,
         DP_reg_pipe11_n145, DP_reg_pipe11_n144, DP_reg_pipe11_n143,
         DP_reg_pipe11_n142, DP_reg_pipe11_n141, DP_reg_pipe11_n140,
         DP_reg_pipe11_n139, DP_reg_pipe11_n138, DP_reg_pipe11_n137,
         DP_reg_pipe11_n136, DP_reg_pipe11_n135, DP_reg_pipe11_n134,
         DP_reg_pipe11_n133, DP_reg_pipe11_n132, DP_reg_pipe11_n131,
         DP_reg_pipe11_n130, DP_reg_pipe11_n129, DP_reg_pipe11_n128,
         DP_reg_pipe11_n127, DP_reg_pipe11_n126, DP_reg_pipe11_n125,
         DP_reg_pipe11_n124, DP_reg_pipe11_n123, DP_reg_pipe11_n122,
         DP_reg_pipe11_n121, DP_reg_pipe11_n120, DP_reg_pipe11_n119,
         DP_reg_pipe11_n118, DP_reg_pipe11_n117, DP_reg_pipe11_n116,
         DP_reg_pipe11_n115, DP_reg_pipe11_n114, DP_reg_pipe11_n113,
         DP_reg_pipe11_n112, DP_reg_pipe11_n111, DP_reg_pipe11_n110,
         DP_reg_pipe11_n109, DP_reg_pipe11_n108, DP_reg_pipe11_n107,
         DP_reg_pipe11_n106, DP_reg_pipe11_n105, DP_reg_pipe11_n104,
         DP_reg_pipe11_n103, DP_reg_pipe11_n102, DP_reg_pipe11_n101,
         DP_reg_pipe11_n100, DP_reg_pipe11_n99, DP_reg_pipe11_n98,
         DP_reg_pipe11_n97, DP_reg_pipe11_n96, DP_reg_pipe11_n95,
         DP_reg_pipe11_n94, DP_reg_pipe11_n93, DP_reg_pipe11_n92,
         DP_reg_pipe11_n91, DP_reg_pipe11_n90, DP_reg_pipe11_n89,
         DP_reg_pipe11_n88, DP_reg_pipe11_n87, DP_reg_pipe11_n86,
         DP_reg_pipe11_n85, DP_reg_pipe11_n84, DP_reg_pipe11_n83,
         DP_reg_pipe11_n82, DP_reg_pipe11_n81, DP_reg_pipe11_n80,
         DP_reg_pipe11_n79, DP_reg_pipe11_n78, DP_reg_pipe11_n77,
         DP_reg_pipe11_n76, DP_reg_pipe11_n75, DP_reg_pipe11_n74,
         DP_reg_pipe11_n73, DP_reg_pipe12_n146, DP_reg_pipe12_n145,
         DP_reg_pipe12_n144, DP_reg_pipe12_n143, DP_reg_pipe12_n142,
         DP_reg_pipe12_n141, DP_reg_pipe12_n140, DP_reg_pipe12_n139,
         DP_reg_pipe12_n138, DP_reg_pipe12_n137, DP_reg_pipe12_n136,
         DP_reg_pipe12_n135, DP_reg_pipe12_n134, DP_reg_pipe12_n133,
         DP_reg_pipe12_n132, DP_reg_pipe12_n131, DP_reg_pipe12_n130,
         DP_reg_pipe12_n129, DP_reg_pipe12_n128, DP_reg_pipe12_n127,
         DP_reg_pipe12_n126, DP_reg_pipe12_n125, DP_reg_pipe12_n124,
         DP_reg_pipe12_n123, DP_reg_pipe12_n122, DP_reg_pipe12_n121,
         DP_reg_pipe12_n120, DP_reg_pipe12_n119, DP_reg_pipe12_n118,
         DP_reg_pipe12_n117, DP_reg_pipe12_n116, DP_reg_pipe12_n115,
         DP_reg_pipe12_n114, DP_reg_pipe12_n113, DP_reg_pipe12_n112,
         DP_reg_pipe12_n111, DP_reg_pipe12_n110, DP_reg_pipe12_n109,
         DP_reg_pipe12_n108, DP_reg_pipe12_n107, DP_reg_pipe12_n106,
         DP_reg_pipe12_n105, DP_reg_pipe12_n104, DP_reg_pipe12_n103,
         DP_reg_pipe12_n102, DP_reg_pipe12_n101, DP_reg_pipe12_n100,
         DP_reg_pipe12_n99, DP_reg_pipe12_n98, DP_reg_pipe12_n97,
         DP_reg_pipe12_n96, DP_reg_pipe12_n95, DP_reg_pipe12_n94,
         DP_reg_pipe12_n93, DP_reg_pipe12_n92, DP_reg_pipe12_n91,
         DP_reg_pipe12_n90, DP_reg_pipe12_n89, DP_reg_pipe12_n88,
         DP_reg_pipe12_n87, DP_reg_pipe12_n86, DP_reg_pipe12_n85,
         DP_reg_pipe12_n84, DP_reg_pipe12_n83, DP_reg_pipe12_n82,
         DP_reg_pipe12_n81, DP_reg_pipe12_n80, DP_reg_pipe12_n79,
         DP_reg_pipe12_n78, DP_reg_pipe12_n77, DP_reg_pipe12_n76,
         DP_reg_pipe12_n75, DP_reg_pipe12_n74, DP_reg_pipe12_n73,
         DP_reg_pipe13_n146, DP_reg_pipe13_n145, DP_reg_pipe13_n144,
         DP_reg_pipe13_n143, DP_reg_pipe13_n142, DP_reg_pipe13_n141,
         DP_reg_pipe13_n140, DP_reg_pipe13_n139, DP_reg_pipe13_n138,
         DP_reg_pipe13_n137, DP_reg_pipe13_n136, DP_reg_pipe13_n135,
         DP_reg_pipe13_n134, DP_reg_pipe13_n133, DP_reg_pipe13_n132,
         DP_reg_pipe13_n131, DP_reg_pipe13_n130, DP_reg_pipe13_n129,
         DP_reg_pipe13_n128, DP_reg_pipe13_n127, DP_reg_pipe13_n126,
         DP_reg_pipe13_n125, DP_reg_pipe13_n124, DP_reg_pipe13_n123,
         DP_reg_pipe13_n122, DP_reg_pipe13_n121, DP_reg_pipe13_n120,
         DP_reg_pipe13_n119, DP_reg_pipe13_n118, DP_reg_pipe13_n117,
         DP_reg_pipe13_n116, DP_reg_pipe13_n115, DP_reg_pipe13_n114,
         DP_reg_pipe13_n113, DP_reg_pipe13_n112, DP_reg_pipe13_n111,
         DP_reg_pipe13_n110, DP_reg_pipe13_n109, DP_reg_pipe13_n108,
         DP_reg_pipe13_n107, DP_reg_pipe13_n106, DP_reg_pipe13_n105,
         DP_reg_pipe13_n104, DP_reg_pipe13_n103, DP_reg_pipe13_n102,
         DP_reg_pipe13_n101, DP_reg_pipe13_n100, DP_reg_pipe13_n99,
         DP_reg_pipe13_n98, DP_reg_pipe13_n97, DP_reg_pipe13_n96,
         DP_reg_pipe13_n95, DP_reg_pipe13_n94, DP_reg_pipe13_n93,
         DP_reg_pipe13_n92, DP_reg_pipe13_n91, DP_reg_pipe13_n90,
         DP_reg_pipe13_n89, DP_reg_pipe13_n88, DP_reg_pipe13_n87,
         DP_reg_pipe13_n86, DP_reg_pipe13_n85, DP_reg_pipe13_n84,
         DP_reg_pipe13_n83, DP_reg_pipe13_n82, DP_reg_pipe13_n81,
         DP_reg_pipe13_n80, DP_reg_pipe13_n79, DP_reg_pipe13_n78,
         DP_reg_pipe13_n77, DP_reg_pipe13_n76, DP_reg_pipe13_n75,
         DP_reg_pipe13_n74, DP_reg_pipe13_n73, DP_reg_out_n75, DP_reg_out_n74,
         DP_reg_out_n73, DP_reg_out_n72, DP_reg_out_n71, DP_reg_out_n70,
         DP_reg_out_n69, DP_reg_out_n68, DP_reg_out_n67, DP_reg_out_n66,
         DP_reg_out_n65, DP_reg_out_n64, DP_reg_out_n63, DP_reg_out_n62,
         DP_reg_out_n61, DP_reg_out_n60, DP_reg_out_n59, DP_reg_out_n58,
         DP_reg_out_n57, DP_reg_out_n56, DP_reg_out_n55, DP_reg_out_n54,
         DP_reg_out_n53, DP_reg_out_n52, DP_reg_out_n51, DP_reg_out_n50,
         DP_reg_out_n49, DP_reg_out_n48, DP_reg_out_n47, DP_reg_out_n46,
         DP_reg_out_n45, DP_reg_out_n44, DP_reg_out_n43, DP_reg_out_n42,
         DP_reg_out_n41, DP_reg_out_n40, DP_reg_out_n39, DP_reg_out_n38,
         DP_reg_out_n37, DP_add_1_root_add_0_root_add_233_carry_1_,
         DP_add_1_root_add_0_root_add_233_carry_2_,
         DP_add_1_root_add_0_root_add_233_carry_3_,
         DP_add_1_root_add_0_root_add_233_carry_4_,
         DP_add_1_root_add_0_root_add_233_carry_5_,
         DP_add_1_root_add_0_root_add_233_carry_6_,
         DP_add_1_root_add_0_root_add_233_carry_7_,
         DP_add_1_root_add_0_root_add_233_carry_8_,
         DP_add_1_root_add_0_root_add_233_carry_9_,
         DP_add_1_root_add_0_root_add_233_carry_10_,
         DP_add_1_root_add_0_root_add_233_carry_11_,
         DP_add_1_root_add_0_root_add_233_carry_12_,
         DP_add_1_root_add_0_root_add_233_carry_13_,
         DP_add_1_root_add_0_root_add_233_carry_14_,
         DP_add_1_root_add_0_root_add_233_carry_15_,
         DP_add_1_root_add_0_root_add_233_carry_16_,
         DP_add_1_root_add_0_root_add_233_carry_17_,
         DP_add_1_root_add_0_root_add_233_carry_18_,
         DP_add_1_root_add_0_root_add_233_carry_19_,
         DP_add_1_root_add_0_root_add_233_carry_20_,
         DP_add_1_root_add_0_root_add_233_carry_21_,
         DP_add_1_root_add_0_root_add_233_carry_22_,
         DP_add_1_root_add_0_root_add_233_carry_23_,
         DP_add_2_root_add_0_root_add_233_carry_1_,
         DP_add_2_root_add_0_root_add_233_carry_2_,
         DP_add_2_root_add_0_root_add_233_carry_3_,
         DP_add_2_root_add_0_root_add_233_carry_4_,
         DP_add_2_root_add_0_root_add_233_carry_5_,
         DP_add_2_root_add_0_root_add_233_carry_6_,
         DP_add_2_root_add_0_root_add_233_carry_7_,
         DP_add_2_root_add_0_root_add_233_carry_8_,
         DP_add_2_root_add_0_root_add_233_carry_9_,
         DP_add_2_root_add_0_root_add_233_carry_10_,
         DP_add_2_root_add_0_root_add_233_carry_11_,
         DP_add_2_root_add_0_root_add_233_carry_12_,
         DP_add_2_root_add_0_root_add_233_carry_13_,
         DP_add_2_root_add_0_root_add_233_carry_14_,
         DP_add_2_root_add_0_root_add_233_carry_15_,
         DP_add_2_root_add_0_root_add_233_carry_16_,
         DP_add_2_root_add_0_root_add_233_carry_17_,
         DP_add_2_root_add_0_root_add_233_carry_18_,
         DP_add_2_root_add_0_root_add_233_carry_19_,
         DP_add_2_root_add_0_root_add_233_carry_20_,
         DP_add_2_root_add_0_root_add_233_carry_21_,
         DP_add_2_root_add_0_root_add_233_carry_22_,
         DP_add_2_root_add_0_root_add_233_carry_23_,
         DP_add_0_root_add_0_root_add_233_n37,
         DP_add_0_root_add_0_root_add_233_n36,
         DP_add_0_root_add_0_root_add_233_n35,
         DP_add_0_root_add_0_root_add_233_n34,
         DP_add_0_root_add_0_root_add_233_n33,
         DP_add_0_root_add_0_root_add_233_n32,
         DP_add_0_root_add_0_root_add_233_n31,
         DP_add_0_root_add_0_root_add_233_n30,
         DP_add_0_root_add_0_root_add_233_n29,
         DP_add_0_root_add_0_root_add_233_n28,
         DP_add_0_root_add_0_root_add_233_n27,
         DP_add_0_root_add_0_root_add_233_n26,
         DP_add_0_root_add_0_root_add_233_n25,
         DP_add_0_root_add_0_root_add_233_n24,
         DP_add_0_root_add_0_root_add_233_n23,
         DP_add_0_root_add_0_root_add_233_n22,
         DP_add_0_root_add_0_root_add_233_n21,
         DP_add_0_root_add_0_root_add_233_n20,
         DP_add_0_root_add_0_root_add_233_n19,
         DP_add_0_root_add_0_root_add_233_n18,
         DP_add_0_root_add_0_root_add_233_n17,
         DP_add_0_root_add_0_root_add_233_n16,
         DP_add_0_root_add_0_root_add_233_n15,
         DP_add_0_root_add_0_root_add_233_n14,
         DP_add_0_root_add_0_root_add_233_n13,
         DP_add_0_root_add_0_root_add_233_n12,
         DP_add_0_root_add_0_root_add_233_n11,
         DP_add_0_root_add_0_root_add_233_n10,
         DP_add_0_root_add_0_root_add_233_n9,
         DP_add_0_root_add_0_root_add_233_n8,
         DP_add_0_root_add_0_root_add_233_n7,
         DP_add_0_root_add_0_root_add_233_n6,
         DP_add_0_root_add_0_root_add_233_n5,
         DP_add_0_root_add_0_root_add_233_n4,
         DP_add_0_root_add_0_root_add_233_n3,
         DP_add_0_root_add_0_root_add_233_n2,
         DP_add_0_root_add_0_root_add_233_n1,
         DP_add_0_root_add_0_root_add_233_carry_11_,
         DP_add_0_root_add_0_root_add_233_carry_12_,
         DP_add_0_root_add_0_root_add_233_carry_13_,
         DP_add_0_root_add_0_root_add_233_carry_14_,
         DP_add_0_root_add_0_root_add_233_carry_15_,
         DP_add_0_root_add_0_root_add_233_carry_16_,
         DP_add_0_root_add_0_root_add_233_carry_17_,
         DP_add_0_root_add_0_root_add_233_carry_18_,
         DP_add_0_root_add_0_root_add_233_carry_19_,
         DP_add_0_root_add_0_root_add_233_carry_20_,
         DP_add_0_root_add_0_root_add_233_carry_21_,
         DP_add_0_root_add_0_root_add_233_carry_22_,
         DP_add_0_root_add_0_root_add_233_carry_23_, DP_mult_219_n2162,
         DP_mult_219_n2161, DP_mult_219_n2160, DP_mult_219_n2159,
         DP_mult_219_n2158, DP_mult_219_n2157, DP_mult_219_n2156,
         DP_mult_219_n2155, DP_mult_219_n2154, DP_mult_219_n2153,
         DP_mult_219_n2152, DP_mult_219_n2151, DP_mult_219_n2150,
         DP_mult_219_n2149, DP_mult_219_n2148, DP_mult_219_n2147,
         DP_mult_219_n2146, DP_mult_219_n2145, DP_mult_219_n2144,
         DP_mult_219_n2143, DP_mult_219_n2142, DP_mult_219_n2141,
         DP_mult_219_n2140, DP_mult_219_n2139, DP_mult_219_n2138,
         DP_mult_219_n2137, DP_mult_219_n2136, DP_mult_219_n2135,
         DP_mult_219_n2134, DP_mult_219_n2133, DP_mult_219_n2132,
         DP_mult_219_n2131, DP_mult_219_n2130, DP_mult_219_n2129,
         DP_mult_219_n2128, DP_mult_219_n2127, DP_mult_219_n2126,
         DP_mult_219_n2125, DP_mult_219_n2124, DP_mult_219_n2123,
         DP_mult_219_n2122, DP_mult_219_n2121, DP_mult_219_n2120,
         DP_mult_219_n2119, DP_mult_219_n2118, DP_mult_219_n2117,
         DP_mult_219_n2116, DP_mult_219_n2115, DP_mult_219_n2114,
         DP_mult_219_n2113, DP_mult_219_n2112, DP_mult_219_n2111,
         DP_mult_219_n2110, DP_mult_219_n2109, DP_mult_219_n2108,
         DP_mult_219_n2107, DP_mult_219_n2106, DP_mult_219_n2105,
         DP_mult_219_n2104, DP_mult_219_n2103, DP_mult_219_n2102,
         DP_mult_219_n2101, DP_mult_219_n2100, DP_mult_219_n2099,
         DP_mult_219_n2098, DP_mult_219_n2097, DP_mult_219_n2096,
         DP_mult_219_n2095, DP_mult_219_n2094, DP_mult_219_n2093,
         DP_mult_219_n2092, DP_mult_219_n2091, DP_mult_219_n2090,
         DP_mult_219_n2089, DP_mult_219_n2088, DP_mult_219_n2087,
         DP_mult_219_n2086, DP_mult_219_n2085, DP_mult_219_n2084,
         DP_mult_219_n2083, DP_mult_219_n2082, DP_mult_219_n2081,
         DP_mult_219_n2080, DP_mult_219_n2079, DP_mult_219_n2078,
         DP_mult_219_n2077, DP_mult_219_n2076, DP_mult_219_n2075,
         DP_mult_219_n2074, DP_mult_219_n2073, DP_mult_219_n2072,
         DP_mult_219_n2071, DP_mult_219_n2070, DP_mult_219_n2069,
         DP_mult_219_n2068, DP_mult_219_n2067, DP_mult_219_n2066,
         DP_mult_219_n2065, DP_mult_219_n2064, DP_mult_219_n2063,
         DP_mult_219_n2062, DP_mult_219_n2061, DP_mult_219_n2060,
         DP_mult_219_n2059, DP_mult_219_n2058, DP_mult_219_n2057,
         DP_mult_219_n2056, DP_mult_219_n2055, DP_mult_219_n2054,
         DP_mult_219_n2053, DP_mult_219_n2052, DP_mult_219_n2051,
         DP_mult_219_n2050, DP_mult_219_n2049, DP_mult_219_n2048,
         DP_mult_219_n2047, DP_mult_219_n2046, DP_mult_219_n2045,
         DP_mult_219_n2044, DP_mult_219_n2043, DP_mult_219_n2042,
         DP_mult_219_n2041, DP_mult_219_n2040, DP_mult_219_n2039,
         DP_mult_219_n2038, DP_mult_219_n2037, DP_mult_219_n2036,
         DP_mult_219_n2035, DP_mult_219_n2034, DP_mult_219_n2033,
         DP_mult_219_n2032, DP_mult_219_n2031, DP_mult_219_n2030,
         DP_mult_219_n2029, DP_mult_219_n2028, DP_mult_219_n2027,
         DP_mult_219_n2026, DP_mult_219_n2025, DP_mult_219_n2024,
         DP_mult_219_n2023, DP_mult_219_n2022, DP_mult_219_n2021,
         DP_mult_219_n2020, DP_mult_219_n2019, DP_mult_219_n2018,
         DP_mult_219_n2017, DP_mult_219_n2016, DP_mult_219_n2015,
         DP_mult_219_n2014, DP_mult_219_n2013, DP_mult_219_n2012,
         DP_mult_219_n2011, DP_mult_219_n2010, DP_mult_219_n2009,
         DP_mult_219_n2008, DP_mult_219_n2007, DP_mult_219_n2006,
         DP_mult_219_n2005, DP_mult_219_n2004, DP_mult_219_n2003,
         DP_mult_219_n2002, DP_mult_219_n2001, DP_mult_219_n2000,
         DP_mult_219_n1999, DP_mult_219_n1998, DP_mult_219_n1997,
         DP_mult_219_n1996, DP_mult_219_n1995, DP_mult_219_n1994,
         DP_mult_219_n1993, DP_mult_219_n1992, DP_mult_219_n1991,
         DP_mult_219_n1990, DP_mult_219_n1989, DP_mult_219_n1988,
         DP_mult_219_n1987, DP_mult_219_n1986, DP_mult_219_n1985,
         DP_mult_219_n1984, DP_mult_219_n1983, DP_mult_219_n1982,
         DP_mult_219_n1981, DP_mult_219_n1980, DP_mult_219_n1979,
         DP_mult_219_n1978, DP_mult_219_n1977, DP_mult_219_n1976,
         DP_mult_219_n1975, DP_mult_219_n1974, DP_mult_219_n1973,
         DP_mult_219_n1972, DP_mult_219_n1971, DP_mult_219_n1970,
         DP_mult_219_n1969, DP_mult_219_n1968, DP_mult_219_n1967,
         DP_mult_219_n1966, DP_mult_219_n1965, DP_mult_219_n1964,
         DP_mult_219_n1963, DP_mult_219_n1962, DP_mult_219_n1961,
         DP_mult_219_n1960, DP_mult_219_n1959, DP_mult_219_n1958,
         DP_mult_219_n1957, DP_mult_219_n1956, DP_mult_219_n1955,
         DP_mult_219_n1954, DP_mult_219_n1953, DP_mult_219_n1952,
         DP_mult_219_n1951, DP_mult_219_n1950, DP_mult_219_n1949,
         DP_mult_219_n1948, DP_mult_219_n1947, DP_mult_219_n1946,
         DP_mult_219_n1945, DP_mult_219_n1944, DP_mult_219_n1943,
         DP_mult_219_n1942, DP_mult_219_n1941, DP_mult_219_n1940,
         DP_mult_219_n1939, DP_mult_219_n1938, DP_mult_219_n1937,
         DP_mult_219_n1936, DP_mult_219_n1935, DP_mult_219_n1934,
         DP_mult_219_n1933, DP_mult_219_n1932, DP_mult_219_n1931,
         DP_mult_219_n1930, DP_mult_219_n1929, DP_mult_219_n1928,
         DP_mult_219_n1927, DP_mult_219_n1926, DP_mult_219_n1925,
         DP_mult_219_n1924, DP_mult_219_n1923, DP_mult_219_n1922,
         DP_mult_219_n1921, DP_mult_219_n1920, DP_mult_219_n1919,
         DP_mult_219_n1918, DP_mult_219_n1917, DP_mult_219_n1916,
         DP_mult_219_n1915, DP_mult_219_n1914, DP_mult_219_n1913,
         DP_mult_219_n1912, DP_mult_219_n1911, DP_mult_219_n1910,
         DP_mult_219_n1909, DP_mult_219_n1908, DP_mult_219_n1907,
         DP_mult_219_n1906, DP_mult_219_n1905, DP_mult_219_n1904,
         DP_mult_219_n1903, DP_mult_219_n1902, DP_mult_219_n1901,
         DP_mult_219_n1900, DP_mult_219_n1899, DP_mult_219_n1898,
         DP_mult_219_n1897, DP_mult_219_n1896, DP_mult_219_n1895,
         DP_mult_219_n1894, DP_mult_219_n1893, DP_mult_219_n1892,
         DP_mult_219_n1891, DP_mult_219_n1890, DP_mult_219_n1889,
         DP_mult_219_n1888, DP_mult_219_n1887, DP_mult_219_n1886,
         DP_mult_219_n1885, DP_mult_219_n1884, DP_mult_219_n1883,
         DP_mult_219_n1882, DP_mult_219_n1881, DP_mult_219_n1880,
         DP_mult_219_n1879, DP_mult_219_n1878, DP_mult_219_n1877,
         DP_mult_219_n1876, DP_mult_219_n1875, DP_mult_219_n1874,
         DP_mult_219_n1873, DP_mult_219_n1872, DP_mult_219_n1871,
         DP_mult_219_n1870, DP_mult_219_n1869, DP_mult_219_n1868,
         DP_mult_219_n1867, DP_mult_219_n1866, DP_mult_219_n1865,
         DP_mult_219_n1864, DP_mult_219_n1863, DP_mult_219_n1862,
         DP_mult_219_n1861, DP_mult_219_n1860, DP_mult_219_n1859,
         DP_mult_219_n1858, DP_mult_219_n1857, DP_mult_219_n1856,
         DP_mult_219_n1855, DP_mult_219_n1854, DP_mult_219_n1853,
         DP_mult_219_n1852, DP_mult_219_n1851, DP_mult_219_n1850,
         DP_mult_219_n1849, DP_mult_219_n1848, DP_mult_219_n1847,
         DP_mult_219_n1846, DP_mult_219_n1845, DP_mult_219_n1844,
         DP_mult_219_n1843, DP_mult_219_n1842, DP_mult_219_n1841,
         DP_mult_219_n1840, DP_mult_219_n1839, DP_mult_219_n1838,
         DP_mult_219_n1837, DP_mult_219_n1836, DP_mult_219_n1835,
         DP_mult_219_n1834, DP_mult_219_n1833, DP_mult_219_n1832,
         DP_mult_219_n1831, DP_mult_219_n1830, DP_mult_219_n1829,
         DP_mult_219_n1828, DP_mult_219_n1827, DP_mult_219_n1826,
         DP_mult_219_n1825, DP_mult_219_n1824, DP_mult_219_n1823,
         DP_mult_219_n1822, DP_mult_219_n1821, DP_mult_219_n1820,
         DP_mult_219_n1819, DP_mult_219_n1818, DP_mult_219_n1817,
         DP_mult_219_n1816, DP_mult_219_n1815, DP_mult_219_n1814,
         DP_mult_219_n1813, DP_mult_219_n1812, DP_mult_219_n1811,
         DP_mult_219_n1810, DP_mult_219_n1809, DP_mult_219_n1808,
         DP_mult_219_n1807, DP_mult_219_n1806, DP_mult_219_n1805,
         DP_mult_219_n1804, DP_mult_219_n1803, DP_mult_219_n1802,
         DP_mult_219_n1801, DP_mult_219_n1800, DP_mult_219_n1799,
         DP_mult_219_n1798, DP_mult_219_n1797, DP_mult_219_n1796,
         DP_mult_219_n1795, DP_mult_219_n1794, DP_mult_219_n1793,
         DP_mult_219_n1792, DP_mult_219_n1791, DP_mult_219_n1790,
         DP_mult_219_n1789, DP_mult_219_n1788, DP_mult_219_n1787,
         DP_mult_219_n1786, DP_mult_219_n1785, DP_mult_219_n1784,
         DP_mult_219_n1783, DP_mult_219_n1782, DP_mult_219_n1781,
         DP_mult_219_n1780, DP_mult_219_n1779, DP_mult_219_n1778,
         DP_mult_219_n1777, DP_mult_219_n1776, DP_mult_219_n1775,
         DP_mult_219_n1774, DP_mult_219_n1773, DP_mult_219_n1772,
         DP_mult_219_n1771, DP_mult_219_n1770, DP_mult_219_n1769,
         DP_mult_219_n1768, DP_mult_219_n1767, DP_mult_219_n1766,
         DP_mult_219_n1765, DP_mult_219_n1764, DP_mult_219_n1763,
         DP_mult_219_n1762, DP_mult_219_n1761, DP_mult_219_n1760,
         DP_mult_219_n1759, DP_mult_219_n1758, DP_mult_219_n1757,
         DP_mult_219_n1756, DP_mult_219_n1755, DP_mult_219_n1754,
         DP_mult_219_n1753, DP_mult_219_n1752, DP_mult_219_n1751,
         DP_mult_219_n1750, DP_mult_219_n1749, DP_mult_219_n1748,
         DP_mult_219_n1747, DP_mult_219_n1746, DP_mult_219_n1745,
         DP_mult_219_n1744, DP_mult_219_n1743, DP_mult_219_n1742,
         DP_mult_219_n1741, DP_mult_219_n1740, DP_mult_219_n1739,
         DP_mult_219_n1738, DP_mult_219_n1737, DP_mult_219_n1736,
         DP_mult_219_n1735, DP_mult_219_n1734, DP_mult_219_n1733,
         DP_mult_219_n1732, DP_mult_219_n1731, DP_mult_219_n1730,
         DP_mult_219_n1729, DP_mult_219_n1728, DP_mult_219_n1727,
         DP_mult_219_n1726, DP_mult_219_n1725, DP_mult_219_n1724,
         DP_mult_219_n1723, DP_mult_219_n1722, DP_mult_219_n1721,
         DP_mult_219_n1720, DP_mult_219_n1719, DP_mult_219_n1718,
         DP_mult_219_n1717, DP_mult_219_n1716, DP_mult_219_n1715,
         DP_mult_219_n1714, DP_mult_219_n1713, DP_mult_219_n1712,
         DP_mult_219_n1711, DP_mult_219_n1710, DP_mult_219_n1709,
         DP_mult_219_n1708, DP_mult_219_n1707, DP_mult_219_n1706,
         DP_mult_219_n1705, DP_mult_219_n1704, DP_mult_219_n1703,
         DP_mult_219_n1702, DP_mult_219_n1701, DP_mult_219_n1700,
         DP_mult_219_n1699, DP_mult_219_n1698, DP_mult_219_n1697,
         DP_mult_219_n1696, DP_mult_219_n1695, DP_mult_219_n1694,
         DP_mult_219_n1693, DP_mult_219_n1692, DP_mult_219_n1691,
         DP_mult_219_n1690, DP_mult_219_n1689, DP_mult_219_n1688,
         DP_mult_219_n1687, DP_mult_219_n1686, DP_mult_219_n1685,
         DP_mult_219_n1684, DP_mult_219_n1683, DP_mult_219_n1682,
         DP_mult_219_n1681, DP_mult_219_n1680, DP_mult_219_n1679,
         DP_mult_219_n1678, DP_mult_219_n1677, DP_mult_219_n1676,
         DP_mult_219_n1675, DP_mult_219_n1674, DP_mult_219_n1673,
         DP_mult_219_n1672, DP_mult_219_n1671, DP_mult_219_n1670,
         DP_mult_219_n1669, DP_mult_219_n1668, DP_mult_219_n1667,
         DP_mult_219_n1666, DP_mult_219_n1665, DP_mult_219_n1664,
         DP_mult_219_n1663, DP_mult_219_n1662, DP_mult_219_n1661,
         DP_mult_219_n1660, DP_mult_219_n1659, DP_mult_219_n1658,
         DP_mult_219_n1657, DP_mult_219_n1656, DP_mult_219_n1655,
         DP_mult_219_n1654, DP_mult_219_n1653, DP_mult_219_n1652,
         DP_mult_219_n1651, DP_mult_219_n1650, DP_mult_219_n1649,
         DP_mult_219_n1648, DP_mult_219_n1647, DP_mult_219_n1646,
         DP_mult_219_n1645, DP_mult_219_n1644, DP_mult_219_n1643,
         DP_mult_219_n1642, DP_mult_219_n1641, DP_mult_219_n1640,
         DP_mult_219_n1639, DP_mult_219_n1638, DP_mult_219_n1637,
         DP_mult_219_n1636, DP_mult_219_n1635, DP_mult_219_n1634,
         DP_mult_219_n1633, DP_mult_219_n1632, DP_mult_219_n1631,
         DP_mult_219_n1630, DP_mult_219_n1629, DP_mult_219_n1628,
         DP_mult_219_n1627, DP_mult_219_n1626, DP_mult_219_n1625,
         DP_mult_219_n1624, DP_mult_219_n1623, DP_mult_219_n1622,
         DP_mult_219_n1621, DP_mult_219_n1620, DP_mult_219_n1619,
         DP_mult_219_n1618, DP_mult_219_n1617, DP_mult_219_n1616,
         DP_mult_219_n1615, DP_mult_219_n1614, DP_mult_219_n1613,
         DP_mult_219_n1612, DP_mult_219_n1611, DP_mult_219_n1610,
         DP_mult_219_n1609, DP_mult_219_n1608, DP_mult_219_n1607,
         DP_mult_219_n1606, DP_mult_219_n1605, DP_mult_219_n1604,
         DP_mult_219_n1603, DP_mult_219_n1602, DP_mult_219_n1601,
         DP_mult_219_n1600, DP_mult_219_n1599, DP_mult_219_n1598,
         DP_mult_219_n1597, DP_mult_219_n1596, DP_mult_219_n1595,
         DP_mult_219_n1594, DP_mult_219_n1593, DP_mult_219_n1592,
         DP_mult_219_n1591, DP_mult_219_n1590, DP_mult_219_n1589,
         DP_mult_219_n1588, DP_mult_219_n1587, DP_mult_219_n1586,
         DP_mult_219_n1585, DP_mult_219_n1584, DP_mult_219_n1583,
         DP_mult_219_n1582, DP_mult_219_n1581, DP_mult_219_n1580,
         DP_mult_219_n1579, DP_mult_219_n1578, DP_mult_219_n1577,
         DP_mult_219_n1576, DP_mult_219_n1575, DP_mult_219_n1574,
         DP_mult_219_n1573, DP_mult_219_n1572, DP_mult_219_n1571,
         DP_mult_219_n1570, DP_mult_219_n1569, DP_mult_219_n1568,
         DP_mult_219_n1567, DP_mult_219_n1566, DP_mult_219_n1565,
         DP_mult_219_n1564, DP_mult_219_n1563, DP_mult_219_n1562,
         DP_mult_219_n1561, DP_mult_219_n1560, DP_mult_219_n1559,
         DP_mult_219_n1558, DP_mult_219_n1557, DP_mult_219_n1556,
         DP_mult_219_n1555, DP_mult_219_n1554, DP_mult_219_n1553,
         DP_mult_219_n1552, DP_mult_219_n1551, DP_mult_219_n1550,
         DP_mult_219_n1549, DP_mult_219_n1548, DP_mult_219_n1547,
         DP_mult_219_n1546, DP_mult_219_n1545, DP_mult_219_n1544,
         DP_mult_219_n1543, DP_mult_219_n1542, DP_mult_219_n1541,
         DP_mult_219_n1540, DP_mult_219_n1539, DP_mult_219_n1538,
         DP_mult_219_n1537, DP_mult_219_n1536, DP_mult_219_n1535,
         DP_mult_219_n1534, DP_mult_219_n1533, DP_mult_219_n1397,
         DP_mult_219_n1396, DP_mult_219_n1395, DP_mult_219_n1394,
         DP_mult_219_n1393, DP_mult_219_n1392, DP_mult_219_n1391,
         DP_mult_219_n1390, DP_mult_219_n1389, DP_mult_219_n1388,
         DP_mult_219_n1387, DP_mult_219_n1386, DP_mult_219_n1385,
         DP_mult_219_n1384, DP_mult_219_n1383, DP_mult_219_n1382,
         DP_mult_219_n1381, DP_mult_219_n1380, DP_mult_219_n1379,
         DP_mult_219_n1378, DP_mult_219_n1377, DP_mult_219_n1376,
         DP_mult_219_n1375, DP_mult_219_n1374, DP_mult_219_n908,
         DP_mult_219_n907, DP_mult_219_n906, DP_mult_219_n904,
         DP_mult_219_n903, DP_mult_219_n902, DP_mult_219_n901,
         DP_mult_219_n900, DP_mult_219_n899, DP_mult_219_n898,
         DP_mult_219_n897, DP_mult_219_n896, DP_mult_219_n895,
         DP_mult_219_n894, DP_mult_219_n893, DP_mult_219_n892,
         DP_mult_219_n891, DP_mult_219_n890, DP_mult_219_n889,
         DP_mult_219_n888, DP_mult_219_n887, DP_mult_219_n886,
         DP_mult_219_n885, DP_mult_219_n884, DP_mult_219_n883,
         DP_mult_219_n882, DP_mult_219_n881, DP_mult_219_n880,
         DP_mult_219_n879, DP_mult_219_n878, DP_mult_219_n877,
         DP_mult_219_n876, DP_mult_219_n875, DP_mult_219_n874,
         DP_mult_219_n873, DP_mult_219_n872, DP_mult_219_n871,
         DP_mult_219_n870, DP_mult_219_n869, DP_mult_219_n868,
         DP_mult_219_n867, DP_mult_219_n866, DP_mult_219_n865,
         DP_mult_219_n864, DP_mult_219_n863, DP_mult_219_n862,
         DP_mult_219_n861, DP_mult_219_n860, DP_mult_219_n859,
         DP_mult_219_n858, DP_mult_219_n857, DP_mult_219_n856,
         DP_mult_219_n855, DP_mult_219_n854, DP_mult_219_n853,
         DP_mult_219_n852, DP_mult_219_n851, DP_mult_219_n850,
         DP_mult_219_n849, DP_mult_219_n848, DP_mult_219_n847,
         DP_mult_219_n846, DP_mult_219_n845, DP_mult_219_n844,
         DP_mult_219_n843, DP_mult_219_n842, DP_mult_219_n841,
         DP_mult_219_n840, DP_mult_219_n839, DP_mult_219_n838,
         DP_mult_219_n837, DP_mult_219_n836, DP_mult_219_n835,
         DP_mult_219_n834, DP_mult_219_n833, DP_mult_219_n832,
         DP_mult_219_n831, DP_mult_219_n830, DP_mult_219_n829,
         DP_mult_219_n828, DP_mult_219_n827, DP_mult_219_n826,
         DP_mult_219_n825, DP_mult_219_n824, DP_mult_219_n823,
         DP_mult_219_n822, DP_mult_219_n821, DP_mult_219_n820,
         DP_mult_219_n819, DP_mult_219_n818, DP_mult_219_n817,
         DP_mult_219_n816, DP_mult_219_n815, DP_mult_219_n814,
         DP_mult_219_n813, DP_mult_219_n812, DP_mult_219_n811,
         DP_mult_219_n810, DP_mult_219_n809, DP_mult_219_n808,
         DP_mult_219_n807, DP_mult_219_n806, DP_mult_219_n805,
         DP_mult_219_n804, DP_mult_219_n803, DP_mult_219_n802,
         DP_mult_219_n801, DP_mult_219_n800, DP_mult_219_n799,
         DP_mult_219_n798, DP_mult_219_n797, DP_mult_219_n796,
         DP_mult_219_n795, DP_mult_219_n794, DP_mult_219_n793,
         DP_mult_219_n792, DP_mult_219_n791, DP_mult_219_n790,
         DP_mult_219_n789, DP_mult_219_n788, DP_mult_219_n787,
         DP_mult_219_n786, DP_mult_219_n785, DP_mult_219_n784,
         DP_mult_219_n783, DP_mult_219_n782, DP_mult_219_n781,
         DP_mult_219_n780, DP_mult_219_n779, DP_mult_219_n778,
         DP_mult_219_n777, DP_mult_219_n776, DP_mult_219_n775,
         DP_mult_219_n774, DP_mult_219_n773, DP_mult_219_n772,
         DP_mult_219_n771, DP_mult_219_n770, DP_mult_219_n769,
         DP_mult_219_n768, DP_mult_219_n767, DP_mult_219_n766,
         DP_mult_219_n765, DP_mult_219_n764, DP_mult_219_n763,
         DP_mult_219_n762, DP_mult_219_n761, DP_mult_219_n760,
         DP_mult_219_n759, DP_mult_219_n758, DP_mult_219_n757,
         DP_mult_219_n756, DP_mult_219_n755, DP_mult_219_n754,
         DP_mult_219_n753, DP_mult_219_n752, DP_mult_219_n751,
         DP_mult_219_n750, DP_mult_219_n749, DP_mult_219_n748,
         DP_mult_219_n747, DP_mult_219_n746, DP_mult_219_n745,
         DP_mult_219_n744, DP_mult_219_n743, DP_mult_219_n742,
         DP_mult_219_n741, DP_mult_219_n740, DP_mult_219_n739,
         DP_mult_219_n738, DP_mult_219_n737, DP_mult_219_n736,
         DP_mult_219_n735, DP_mult_219_n734, DP_mult_219_n733,
         DP_mult_219_n732, DP_mult_219_n731, DP_mult_219_n730,
         DP_mult_219_n729, DP_mult_219_n727, DP_mult_219_n726,
         DP_mult_219_n725, DP_mult_219_n724, DP_mult_219_n723,
         DP_mult_219_n722, DP_mult_219_n721, DP_mult_219_n720,
         DP_mult_219_n719, DP_mult_219_n718, DP_mult_219_n717,
         DP_mult_219_n716, DP_mult_219_n715, DP_mult_219_n714,
         DP_mult_219_n713, DP_mult_219_n712, DP_mult_219_n711,
         DP_mult_219_n710, DP_mult_219_n709, DP_mult_219_n708,
         DP_mult_219_n707, DP_mult_219_n706, DP_mult_219_n688,
         DP_mult_219_n687, DP_mult_219_n686, DP_mult_219_n685,
         DP_mult_219_n684, DP_mult_219_n683, DP_mult_219_n682,
         DP_mult_219_n681, DP_mult_219_n680, DP_mult_219_n679,
         DP_mult_219_n678, DP_mult_219_n677, DP_mult_219_n676,
         DP_mult_219_n675, DP_mult_219_n674, DP_mult_219_n673,
         DP_mult_219_n672, DP_mult_219_n671, DP_mult_219_n670,
         DP_mult_219_n669, DP_mult_219_n668, DP_mult_219_n667,
         DP_mult_219_n666, DP_mult_219_n665, DP_mult_219_n664,
         DP_mult_219_n663, DP_mult_219_n662, DP_mult_219_n661,
         DP_mult_219_n660, DP_mult_219_n659, DP_mult_219_n658,
         DP_mult_219_n657, DP_mult_219_n656, DP_mult_219_n655,
         DP_mult_219_n654, DP_mult_219_n653, DP_mult_219_n652,
         DP_mult_219_n651, DP_mult_219_n650, DP_mult_219_n649,
         DP_mult_219_n648, DP_mult_219_n647, DP_mult_219_n646,
         DP_mult_219_n645, DP_mult_219_n644, DP_mult_219_n643,
         DP_mult_219_n642, DP_mult_219_n641, DP_mult_219_n640,
         DP_mult_219_n639, DP_mult_219_n638, DP_mult_219_n637,
         DP_mult_219_n636, DP_mult_219_n635, DP_mult_219_n634,
         DP_mult_219_n633, DP_mult_219_n632, DP_mult_219_n631,
         DP_mult_219_n630, DP_mult_219_n629, DP_mult_219_n628,
         DP_mult_219_n627, DP_mult_219_n626, DP_mult_219_n625,
         DP_mult_219_n624, DP_mult_219_n623, DP_mult_219_n622,
         DP_mult_219_n621, DP_mult_219_n620, DP_mult_219_n619,
         DP_mult_219_n618, DP_mult_219_n617, DP_mult_219_n616,
         DP_mult_219_n615, DP_mult_219_n614, DP_mult_219_n613,
         DP_mult_219_n612, DP_mult_219_n611, DP_mult_219_n610,
         DP_mult_219_n609, DP_mult_219_n608, DP_mult_219_n607,
         DP_mult_219_n606, DP_mult_219_n605, DP_mult_219_n604,
         DP_mult_219_n603, DP_mult_219_n602, DP_mult_219_n601,
         DP_mult_219_n600, DP_mult_219_n599, DP_mult_219_n598,
         DP_mult_219_n597, DP_mult_219_n596, DP_mult_219_n595,
         DP_mult_219_n594, DP_mult_219_n593, DP_mult_219_n592,
         DP_mult_219_n591, DP_mult_219_n590, DP_mult_219_n589,
         DP_mult_219_n588, DP_mult_219_n587, DP_mult_219_n586,
         DP_mult_219_n585, DP_mult_219_n584, DP_mult_219_n583,
         DP_mult_219_n582, DP_mult_219_n581, DP_mult_219_n580,
         DP_mult_219_n579, DP_mult_219_n578, DP_mult_219_n577,
         DP_mult_219_n576, DP_mult_219_n575, DP_mult_219_n574,
         DP_mult_219_n573, DP_mult_219_n572, DP_mult_219_n571,
         DP_mult_219_n570, DP_mult_219_n569, DP_mult_219_n568,
         DP_mult_219_n567, DP_mult_219_n566, DP_mult_219_n565,
         DP_mult_219_n564, DP_mult_219_n563, DP_mult_219_n562,
         DP_mult_219_n561, DP_mult_219_n560, DP_mult_219_n559,
         DP_mult_219_n558, DP_mult_219_n557, DP_mult_219_n556,
         DP_mult_219_n555, DP_mult_219_n554, DP_mult_219_n553,
         DP_mult_219_n552, DP_mult_219_n551, DP_mult_219_n550,
         DP_mult_219_n549, DP_mult_219_n548, DP_mult_219_n547,
         DP_mult_219_n546, DP_mult_219_n545, DP_mult_219_n544,
         DP_mult_219_n543, DP_mult_219_n542, DP_mult_219_n541,
         DP_mult_219_n540, DP_mult_219_n539, DP_mult_219_n538,
         DP_mult_219_n537, DP_mult_219_n536, DP_mult_219_n535,
         DP_mult_219_n534, DP_mult_219_n533, DP_mult_219_n532,
         DP_mult_219_n531, DP_mult_219_n530, DP_mult_219_n529,
         DP_mult_219_n528, DP_mult_219_n527, DP_mult_219_n526,
         DP_mult_219_n525, DP_mult_219_n524, DP_mult_219_n523,
         DP_mult_219_n522, DP_mult_219_n521, DP_mult_219_n520,
         DP_mult_219_n519, DP_mult_219_n518, DP_mult_219_n517,
         DP_mult_219_n516, DP_mult_219_n515, DP_mult_219_n514,
         DP_mult_219_n513, DP_mult_219_n512, DP_mult_219_n511,
         DP_mult_219_n510, DP_mult_219_n509, DP_mult_219_n508,
         DP_mult_219_n507, DP_mult_219_n506, DP_mult_219_n505,
         DP_mult_219_n504, DP_mult_219_n503, DP_mult_219_n502,
         DP_mult_219_n501, DP_mult_219_n500, DP_mult_219_n499,
         DP_mult_219_n498, DP_mult_219_n497, DP_mult_219_n496,
         DP_mult_219_n495, DP_mult_219_n494, DP_mult_219_n493,
         DP_mult_219_n492, DP_mult_219_n491, DP_mult_219_n490,
         DP_mult_219_n489, DP_mult_219_n488, DP_mult_219_n487,
         DP_mult_219_n486, DP_mult_219_n485, DP_mult_219_n484,
         DP_mult_219_n483, DP_mult_219_n482, DP_mult_219_n481,
         DP_mult_219_n479, DP_mult_219_n478, DP_mult_219_n477,
         DP_mult_219_n476, DP_mult_219_n475, DP_mult_219_n474,
         DP_mult_219_n473, DP_mult_219_n472, DP_mult_219_n471,
         DP_mult_219_n470, DP_mult_219_n469, DP_mult_219_n468,
         DP_mult_219_n467, DP_mult_219_n466, DP_mult_219_n465,
         DP_mult_219_n464, DP_mult_219_n463, DP_mult_219_n462,
         DP_mult_219_n461, DP_mult_219_n460, DP_mult_219_n459,
         DP_mult_219_n458, DP_mult_219_n457, DP_mult_219_n456,
         DP_mult_219_n455, DP_mult_219_n454, DP_mult_219_n453,
         DP_mult_219_n452, DP_mult_219_n451, DP_mult_219_n450,
         DP_mult_219_n449, DP_mult_219_n448, DP_mult_219_n447,
         DP_mult_219_n446, DP_mult_219_n445, DP_mult_219_n444,
         DP_mult_219_n442, DP_mult_219_n441, DP_mult_219_n440,
         DP_mult_219_n439, DP_mult_219_n438, DP_mult_219_n437,
         DP_mult_219_n436, DP_mult_219_n435, DP_mult_219_n434,
         DP_mult_219_n433, DP_mult_219_n432, DP_mult_219_n431,
         DP_mult_219_n430, DP_mult_219_n429, DP_mult_219_n428,
         DP_mult_219_n427, DP_mult_219_n426, DP_mult_219_n425,
         DP_mult_219_n424, DP_mult_219_n423, DP_mult_219_n422,
         DP_mult_219_n421, DP_mult_219_n420, DP_mult_219_n419,
         DP_mult_219_n418, DP_mult_219_n417, DP_mult_219_n416,
         DP_mult_219_n415, DP_mult_219_n414, DP_mult_219_n413,
         DP_mult_219_n411, DP_mult_219_n410, DP_mult_219_n409,
         DP_mult_219_n408, DP_mult_219_n407, DP_mult_219_n406,
         DP_mult_219_n405, DP_mult_219_n404, DP_mult_219_n403,
         DP_mult_219_n402, DP_mult_219_n401, DP_mult_219_n400,
         DP_mult_219_n399, DP_mult_219_n398, DP_mult_219_n397,
         DP_mult_219_n396, DP_mult_219_n395, DP_mult_219_n394,
         DP_mult_219_n393, DP_mult_219_n392, DP_mult_219_n391,
         DP_mult_219_n390, DP_mult_219_n389, DP_mult_219_n387,
         DP_mult_219_n386, DP_mult_219_n385, DP_mult_219_n384,
         DP_mult_219_n383, DP_mult_219_n382, DP_mult_219_n381,
         DP_mult_219_n380, DP_mult_219_n379, DP_mult_219_n378,
         DP_mult_219_n377, DP_mult_219_n376, DP_mult_219_n375,
         DP_mult_219_n374, DP_mult_219_n373, DP_mult_219_n372,
         DP_mult_219_n371, DP_mult_219_n370, DP_mult_219_n368,
         DP_mult_219_n367, DP_mult_219_n366, DP_mult_219_n365,
         DP_mult_219_n364, DP_mult_219_n363, DP_mult_219_n362,
         DP_mult_219_n361, DP_mult_219_n360, DP_mult_219_n359,
         DP_mult_219_n358, DP_mult_219_n356, DP_mult_219_n355,
         DP_mult_219_n354, DP_mult_219_n353, DP_mult_219_n352,
         DP_mult_219_n351, DP_mult_219_n326, DP_mult_219_n325,
         DP_mult_219_n324, DP_mult_219_n323, DP_mult_219_n322,
         DP_mult_219_n321, DP_mult_219_n320, DP_mult_219_n319,
         DP_mult_219_n318, DP_mult_219_n317, DP_mult_219_n316,
         DP_mult_219_n315, DP_mult_219_n314, DP_mult_219_n313,
         DP_mult_219_n312, DP_mult_219_n311, DP_mult_219_n310,
         DP_mult_219_n309, DP_mult_219_n308, DP_mult_219_n307,
         DP_mult_219_n306, DP_mult_219_n305, DP_mult_219_n304,
         DP_mult_219_n303, DP_mult_218_n2162, DP_mult_218_n2161,
         DP_mult_218_n2160, DP_mult_218_n2159, DP_mult_218_n2158,
         DP_mult_218_n2157, DP_mult_218_n2156, DP_mult_218_n2155,
         DP_mult_218_n2154, DP_mult_218_n2153, DP_mult_218_n2152,
         DP_mult_218_n2151, DP_mult_218_n2150, DP_mult_218_n2149,
         DP_mult_218_n2148, DP_mult_218_n2147, DP_mult_218_n2146,
         DP_mult_218_n2145, DP_mult_218_n2144, DP_mult_218_n2143,
         DP_mult_218_n2142, DP_mult_218_n2141, DP_mult_218_n2140,
         DP_mult_218_n2139, DP_mult_218_n2138, DP_mult_218_n2137,
         DP_mult_218_n2136, DP_mult_218_n2135, DP_mult_218_n2134,
         DP_mult_218_n2133, DP_mult_218_n2132, DP_mult_218_n2131,
         DP_mult_218_n2130, DP_mult_218_n2129, DP_mult_218_n2128,
         DP_mult_218_n2127, DP_mult_218_n2126, DP_mult_218_n2125,
         DP_mult_218_n2124, DP_mult_218_n2123, DP_mult_218_n2122,
         DP_mult_218_n2121, DP_mult_218_n2120, DP_mult_218_n2119,
         DP_mult_218_n2118, DP_mult_218_n2117, DP_mult_218_n2116,
         DP_mult_218_n2115, DP_mult_218_n2114, DP_mult_218_n2113,
         DP_mult_218_n2112, DP_mult_218_n2111, DP_mult_218_n2110,
         DP_mult_218_n2109, DP_mult_218_n2108, DP_mult_218_n2107,
         DP_mult_218_n2106, DP_mult_218_n2105, DP_mult_218_n2104,
         DP_mult_218_n2103, DP_mult_218_n2102, DP_mult_218_n2101,
         DP_mult_218_n2100, DP_mult_218_n2099, DP_mult_218_n2098,
         DP_mult_218_n2097, DP_mult_218_n2096, DP_mult_218_n2095,
         DP_mult_218_n2094, DP_mult_218_n2093, DP_mult_218_n2092,
         DP_mult_218_n2091, DP_mult_218_n2090, DP_mult_218_n2089,
         DP_mult_218_n2088, DP_mult_218_n2087, DP_mult_218_n2086,
         DP_mult_218_n2085, DP_mult_218_n2084, DP_mult_218_n2083,
         DP_mult_218_n2082, DP_mult_218_n2081, DP_mult_218_n2080,
         DP_mult_218_n2079, DP_mult_218_n2078, DP_mult_218_n2077,
         DP_mult_218_n2076, DP_mult_218_n2075, DP_mult_218_n2074,
         DP_mult_218_n2073, DP_mult_218_n2072, DP_mult_218_n2071,
         DP_mult_218_n2070, DP_mult_218_n2069, DP_mult_218_n2068,
         DP_mult_218_n2067, DP_mult_218_n2066, DP_mult_218_n2065,
         DP_mult_218_n2064, DP_mult_218_n2063, DP_mult_218_n2062,
         DP_mult_218_n2061, DP_mult_218_n2060, DP_mult_218_n2059,
         DP_mult_218_n2058, DP_mult_218_n2057, DP_mult_218_n2056,
         DP_mult_218_n2055, DP_mult_218_n2054, DP_mult_218_n2053,
         DP_mult_218_n2052, DP_mult_218_n2051, DP_mult_218_n2050,
         DP_mult_218_n2049, DP_mult_218_n2048, DP_mult_218_n2047,
         DP_mult_218_n2046, DP_mult_218_n2045, DP_mult_218_n2044,
         DP_mult_218_n2043, DP_mult_218_n2042, DP_mult_218_n2041,
         DP_mult_218_n2040, DP_mult_218_n2039, DP_mult_218_n2038,
         DP_mult_218_n2037, DP_mult_218_n2036, DP_mult_218_n2035,
         DP_mult_218_n2034, DP_mult_218_n2033, DP_mult_218_n2032,
         DP_mult_218_n2031, DP_mult_218_n2030, DP_mult_218_n2029,
         DP_mult_218_n2028, DP_mult_218_n2027, DP_mult_218_n2026,
         DP_mult_218_n2025, DP_mult_218_n2024, DP_mult_218_n2023,
         DP_mult_218_n2022, DP_mult_218_n2021, DP_mult_218_n2020,
         DP_mult_218_n2019, DP_mult_218_n2018, DP_mult_218_n2017,
         DP_mult_218_n2016, DP_mult_218_n2015, DP_mult_218_n2014,
         DP_mult_218_n2013, DP_mult_218_n2012, DP_mult_218_n2011,
         DP_mult_218_n2010, DP_mult_218_n2009, DP_mult_218_n2008,
         DP_mult_218_n2007, DP_mult_218_n2006, DP_mult_218_n2005,
         DP_mult_218_n2004, DP_mult_218_n2003, DP_mult_218_n2002,
         DP_mult_218_n2001, DP_mult_218_n2000, DP_mult_218_n1999,
         DP_mult_218_n1998, DP_mult_218_n1997, DP_mult_218_n1996,
         DP_mult_218_n1995, DP_mult_218_n1994, DP_mult_218_n1993,
         DP_mult_218_n1992, DP_mult_218_n1991, DP_mult_218_n1990,
         DP_mult_218_n1989, DP_mult_218_n1988, DP_mult_218_n1987,
         DP_mult_218_n1986, DP_mult_218_n1985, DP_mult_218_n1984,
         DP_mult_218_n1983, DP_mult_218_n1982, DP_mult_218_n1981,
         DP_mult_218_n1980, DP_mult_218_n1979, DP_mult_218_n1978,
         DP_mult_218_n1977, DP_mult_218_n1976, DP_mult_218_n1975,
         DP_mult_218_n1974, DP_mult_218_n1973, DP_mult_218_n1972,
         DP_mult_218_n1971, DP_mult_218_n1970, DP_mult_218_n1969,
         DP_mult_218_n1968, DP_mult_218_n1967, DP_mult_218_n1966,
         DP_mult_218_n1965, DP_mult_218_n1964, DP_mult_218_n1963,
         DP_mult_218_n1962, DP_mult_218_n1961, DP_mult_218_n1960,
         DP_mult_218_n1959, DP_mult_218_n1958, DP_mult_218_n1957,
         DP_mult_218_n1956, DP_mult_218_n1955, DP_mult_218_n1954,
         DP_mult_218_n1953, DP_mult_218_n1952, DP_mult_218_n1951,
         DP_mult_218_n1950, DP_mult_218_n1949, DP_mult_218_n1948,
         DP_mult_218_n1947, DP_mult_218_n1946, DP_mult_218_n1945,
         DP_mult_218_n1944, DP_mult_218_n1943, DP_mult_218_n1942,
         DP_mult_218_n1941, DP_mult_218_n1940, DP_mult_218_n1939,
         DP_mult_218_n1938, DP_mult_218_n1937, DP_mult_218_n1936,
         DP_mult_218_n1935, DP_mult_218_n1934, DP_mult_218_n1933,
         DP_mult_218_n1932, DP_mult_218_n1931, DP_mult_218_n1930,
         DP_mult_218_n1929, DP_mult_218_n1928, DP_mult_218_n1927,
         DP_mult_218_n1926, DP_mult_218_n1925, DP_mult_218_n1924,
         DP_mult_218_n1923, DP_mult_218_n1922, DP_mult_218_n1921,
         DP_mult_218_n1920, DP_mult_218_n1919, DP_mult_218_n1918,
         DP_mult_218_n1917, DP_mult_218_n1916, DP_mult_218_n1915,
         DP_mult_218_n1914, DP_mult_218_n1913, DP_mult_218_n1912,
         DP_mult_218_n1911, DP_mult_218_n1910, DP_mult_218_n1909,
         DP_mult_218_n1908, DP_mult_218_n1907, DP_mult_218_n1906,
         DP_mult_218_n1905, DP_mult_218_n1904, DP_mult_218_n1903,
         DP_mult_218_n1902, DP_mult_218_n1901, DP_mult_218_n1900,
         DP_mult_218_n1899, DP_mult_218_n1898, DP_mult_218_n1897,
         DP_mult_218_n1896, DP_mult_218_n1895, DP_mult_218_n1894,
         DP_mult_218_n1893, DP_mult_218_n1892, DP_mult_218_n1891,
         DP_mult_218_n1890, DP_mult_218_n1889, DP_mult_218_n1888,
         DP_mult_218_n1887, DP_mult_218_n1886, DP_mult_218_n1885,
         DP_mult_218_n1884, DP_mult_218_n1883, DP_mult_218_n1882,
         DP_mult_218_n1881, DP_mult_218_n1880, DP_mult_218_n1879,
         DP_mult_218_n1878, DP_mult_218_n1877, DP_mult_218_n1876,
         DP_mult_218_n1875, DP_mult_218_n1874, DP_mult_218_n1873,
         DP_mult_218_n1872, DP_mult_218_n1871, DP_mult_218_n1870,
         DP_mult_218_n1869, DP_mult_218_n1868, DP_mult_218_n1867,
         DP_mult_218_n1866, DP_mult_218_n1865, DP_mult_218_n1864,
         DP_mult_218_n1863, DP_mult_218_n1862, DP_mult_218_n1861,
         DP_mult_218_n1860, DP_mult_218_n1859, DP_mult_218_n1858,
         DP_mult_218_n1857, DP_mult_218_n1856, DP_mult_218_n1855,
         DP_mult_218_n1854, DP_mult_218_n1853, DP_mult_218_n1852,
         DP_mult_218_n1851, DP_mult_218_n1850, DP_mult_218_n1849,
         DP_mult_218_n1848, DP_mult_218_n1847, DP_mult_218_n1846,
         DP_mult_218_n1845, DP_mult_218_n1844, DP_mult_218_n1843,
         DP_mult_218_n1842, DP_mult_218_n1841, DP_mult_218_n1840,
         DP_mult_218_n1839, DP_mult_218_n1838, DP_mult_218_n1837,
         DP_mult_218_n1836, DP_mult_218_n1835, DP_mult_218_n1834,
         DP_mult_218_n1833, DP_mult_218_n1832, DP_mult_218_n1831,
         DP_mult_218_n1830, DP_mult_218_n1829, DP_mult_218_n1828,
         DP_mult_218_n1827, DP_mult_218_n1826, DP_mult_218_n1825,
         DP_mult_218_n1824, DP_mult_218_n1823, DP_mult_218_n1822,
         DP_mult_218_n1821, DP_mult_218_n1820, DP_mult_218_n1819,
         DP_mult_218_n1818, DP_mult_218_n1817, DP_mult_218_n1816,
         DP_mult_218_n1815, DP_mult_218_n1814, DP_mult_218_n1813,
         DP_mult_218_n1812, DP_mult_218_n1811, DP_mult_218_n1810,
         DP_mult_218_n1809, DP_mult_218_n1808, DP_mult_218_n1807,
         DP_mult_218_n1806, DP_mult_218_n1805, DP_mult_218_n1804,
         DP_mult_218_n1803, DP_mult_218_n1802, DP_mult_218_n1801,
         DP_mult_218_n1800, DP_mult_218_n1799, DP_mult_218_n1798,
         DP_mult_218_n1797, DP_mult_218_n1796, DP_mult_218_n1795,
         DP_mult_218_n1794, DP_mult_218_n1793, DP_mult_218_n1792,
         DP_mult_218_n1791, DP_mult_218_n1790, DP_mult_218_n1789,
         DP_mult_218_n1788, DP_mult_218_n1787, DP_mult_218_n1786,
         DP_mult_218_n1785, DP_mult_218_n1784, DP_mult_218_n1783,
         DP_mult_218_n1782, DP_mult_218_n1781, DP_mult_218_n1780,
         DP_mult_218_n1779, DP_mult_218_n1778, DP_mult_218_n1777,
         DP_mult_218_n1776, DP_mult_218_n1775, DP_mult_218_n1774,
         DP_mult_218_n1773, DP_mult_218_n1772, DP_mult_218_n1771,
         DP_mult_218_n1770, DP_mult_218_n1769, DP_mult_218_n1768,
         DP_mult_218_n1767, DP_mult_218_n1766, DP_mult_218_n1765,
         DP_mult_218_n1764, DP_mult_218_n1763, DP_mult_218_n1762,
         DP_mult_218_n1761, DP_mult_218_n1760, DP_mult_218_n1759,
         DP_mult_218_n1758, DP_mult_218_n1757, DP_mult_218_n1756,
         DP_mult_218_n1755, DP_mult_218_n1754, DP_mult_218_n1753,
         DP_mult_218_n1752, DP_mult_218_n1751, DP_mult_218_n1750,
         DP_mult_218_n1749, DP_mult_218_n1748, DP_mult_218_n1747,
         DP_mult_218_n1746, DP_mult_218_n1745, DP_mult_218_n1744,
         DP_mult_218_n1743, DP_mult_218_n1742, DP_mult_218_n1741,
         DP_mult_218_n1740, DP_mult_218_n1739, DP_mult_218_n1738,
         DP_mult_218_n1737, DP_mult_218_n1736, DP_mult_218_n1735,
         DP_mult_218_n1734, DP_mult_218_n1733, DP_mult_218_n1732,
         DP_mult_218_n1731, DP_mult_218_n1730, DP_mult_218_n1729,
         DP_mult_218_n1728, DP_mult_218_n1727, DP_mult_218_n1726,
         DP_mult_218_n1725, DP_mult_218_n1724, DP_mult_218_n1723,
         DP_mult_218_n1722, DP_mult_218_n1721, DP_mult_218_n1720,
         DP_mult_218_n1719, DP_mult_218_n1718, DP_mult_218_n1717,
         DP_mult_218_n1716, DP_mult_218_n1715, DP_mult_218_n1714,
         DP_mult_218_n1713, DP_mult_218_n1712, DP_mult_218_n1711,
         DP_mult_218_n1710, DP_mult_218_n1709, DP_mult_218_n1708,
         DP_mult_218_n1707, DP_mult_218_n1706, DP_mult_218_n1705,
         DP_mult_218_n1704, DP_mult_218_n1703, DP_mult_218_n1702,
         DP_mult_218_n1701, DP_mult_218_n1700, DP_mult_218_n1699,
         DP_mult_218_n1698, DP_mult_218_n1697, DP_mult_218_n1696,
         DP_mult_218_n1695, DP_mult_218_n1694, DP_mult_218_n1693,
         DP_mult_218_n1692, DP_mult_218_n1691, DP_mult_218_n1690,
         DP_mult_218_n1689, DP_mult_218_n1688, DP_mult_218_n1687,
         DP_mult_218_n1686, DP_mult_218_n1685, DP_mult_218_n1684,
         DP_mult_218_n1683, DP_mult_218_n1682, DP_mult_218_n1681,
         DP_mult_218_n1680, DP_mult_218_n1679, DP_mult_218_n1678,
         DP_mult_218_n1677, DP_mult_218_n1676, DP_mult_218_n1675,
         DP_mult_218_n1674, DP_mult_218_n1673, DP_mult_218_n1672,
         DP_mult_218_n1671, DP_mult_218_n1670, DP_mult_218_n1669,
         DP_mult_218_n1668, DP_mult_218_n1667, DP_mult_218_n1666,
         DP_mult_218_n1665, DP_mult_218_n1664, DP_mult_218_n1663,
         DP_mult_218_n1662, DP_mult_218_n1661, DP_mult_218_n1660,
         DP_mult_218_n1659, DP_mult_218_n1658, DP_mult_218_n1657,
         DP_mult_218_n1656, DP_mult_218_n1655, DP_mult_218_n1654,
         DP_mult_218_n1653, DP_mult_218_n1652, DP_mult_218_n1651,
         DP_mult_218_n1650, DP_mult_218_n1649, DP_mult_218_n1648,
         DP_mult_218_n1647, DP_mult_218_n1646, DP_mult_218_n1645,
         DP_mult_218_n1644, DP_mult_218_n1643, DP_mult_218_n1642,
         DP_mult_218_n1641, DP_mult_218_n1640, DP_mult_218_n1639,
         DP_mult_218_n1638, DP_mult_218_n1637, DP_mult_218_n1636,
         DP_mult_218_n1635, DP_mult_218_n1634, DP_mult_218_n1633,
         DP_mult_218_n1632, DP_mult_218_n1631, DP_mult_218_n1630,
         DP_mult_218_n1629, DP_mult_218_n1628, DP_mult_218_n1627,
         DP_mult_218_n1626, DP_mult_218_n1625, DP_mult_218_n1624,
         DP_mult_218_n1623, DP_mult_218_n1622, DP_mult_218_n1621,
         DP_mult_218_n1620, DP_mult_218_n1619, DP_mult_218_n1618,
         DP_mult_218_n1617, DP_mult_218_n1616, DP_mult_218_n1615,
         DP_mult_218_n1614, DP_mult_218_n1613, DP_mult_218_n1612,
         DP_mult_218_n1611, DP_mult_218_n1610, DP_mult_218_n1609,
         DP_mult_218_n1608, DP_mult_218_n1607, DP_mult_218_n1606,
         DP_mult_218_n1605, DP_mult_218_n1604, DP_mult_218_n1603,
         DP_mult_218_n1602, DP_mult_218_n1601, DP_mult_218_n1600,
         DP_mult_218_n1599, DP_mult_218_n1598, DP_mult_218_n1597,
         DP_mult_218_n1596, DP_mult_218_n1595, DP_mult_218_n1594,
         DP_mult_218_n1593, DP_mult_218_n1592, DP_mult_218_n1591,
         DP_mult_218_n1590, DP_mult_218_n1589, DP_mult_218_n1588,
         DP_mult_218_n1587, DP_mult_218_n1586, DP_mult_218_n1585,
         DP_mult_218_n1584, DP_mult_218_n1583, DP_mult_218_n1582,
         DP_mult_218_n1581, DP_mult_218_n1580, DP_mult_218_n1579,
         DP_mult_218_n1578, DP_mult_218_n1577, DP_mult_218_n1576,
         DP_mult_218_n1575, DP_mult_218_n1574, DP_mult_218_n1573,
         DP_mult_218_n1572, DP_mult_218_n1571, DP_mult_218_n1570,
         DP_mult_218_n1569, DP_mult_218_n1568, DP_mult_218_n1567,
         DP_mult_218_n1566, DP_mult_218_n1565, DP_mult_218_n1564,
         DP_mult_218_n1563, DP_mult_218_n1562, DP_mult_218_n1561,
         DP_mult_218_n1560, DP_mult_218_n1559, DP_mult_218_n1558,
         DP_mult_218_n1557, DP_mult_218_n1556, DP_mult_218_n1555,
         DP_mult_218_n1554, DP_mult_218_n1553, DP_mult_218_n1552,
         DP_mult_218_n1551, DP_mult_218_n1550, DP_mult_218_n1549,
         DP_mult_218_n1548, DP_mult_218_n1547, DP_mult_218_n1546,
         DP_mult_218_n1545, DP_mult_218_n1544, DP_mult_218_n1543,
         DP_mult_218_n1542, DP_mult_218_n1541, DP_mult_218_n1540,
         DP_mult_218_n1539, DP_mult_218_n1538, DP_mult_218_n1537,
         DP_mult_218_n1536, DP_mult_218_n1535, DP_mult_218_n1534,
         DP_mult_218_n1533, DP_mult_218_n1397, DP_mult_218_n1396,
         DP_mult_218_n1395, DP_mult_218_n1394, DP_mult_218_n1393,
         DP_mult_218_n1392, DP_mult_218_n1391, DP_mult_218_n1390,
         DP_mult_218_n1389, DP_mult_218_n1388, DP_mult_218_n1387,
         DP_mult_218_n1386, DP_mult_218_n1385, DP_mult_218_n1384,
         DP_mult_218_n1383, DP_mult_218_n1382, DP_mult_218_n1381,
         DP_mult_218_n1380, DP_mult_218_n1379, DP_mult_218_n1378,
         DP_mult_218_n1377, DP_mult_218_n1376, DP_mult_218_n1375,
         DP_mult_218_n1374, DP_mult_218_n908, DP_mult_218_n907,
         DP_mult_218_n906, DP_mult_218_n904, DP_mult_218_n903,
         DP_mult_218_n902, DP_mult_218_n901, DP_mult_218_n900,
         DP_mult_218_n899, DP_mult_218_n898, DP_mult_218_n897,
         DP_mult_218_n896, DP_mult_218_n895, DP_mult_218_n894,
         DP_mult_218_n893, DP_mult_218_n892, DP_mult_218_n891,
         DP_mult_218_n890, DP_mult_218_n889, DP_mult_218_n888,
         DP_mult_218_n887, DP_mult_218_n886, DP_mult_218_n885,
         DP_mult_218_n884, DP_mult_218_n883, DP_mult_218_n882,
         DP_mult_218_n881, DP_mult_218_n880, DP_mult_218_n879,
         DP_mult_218_n878, DP_mult_218_n877, DP_mult_218_n876,
         DP_mult_218_n875, DP_mult_218_n874, DP_mult_218_n873,
         DP_mult_218_n872, DP_mult_218_n871, DP_mult_218_n870,
         DP_mult_218_n869, DP_mult_218_n868, DP_mult_218_n867,
         DP_mult_218_n866, DP_mult_218_n865, DP_mult_218_n864,
         DP_mult_218_n863, DP_mult_218_n862, DP_mult_218_n861,
         DP_mult_218_n860, DP_mult_218_n859, DP_mult_218_n858,
         DP_mult_218_n857, DP_mult_218_n856, DP_mult_218_n855,
         DP_mult_218_n854, DP_mult_218_n853, DP_mult_218_n852,
         DP_mult_218_n851, DP_mult_218_n850, DP_mult_218_n849,
         DP_mult_218_n848, DP_mult_218_n847, DP_mult_218_n846,
         DP_mult_218_n845, DP_mult_218_n844, DP_mult_218_n843,
         DP_mult_218_n842, DP_mult_218_n841, DP_mult_218_n840,
         DP_mult_218_n839, DP_mult_218_n838, DP_mult_218_n837,
         DP_mult_218_n836, DP_mult_218_n835, DP_mult_218_n834,
         DP_mult_218_n833, DP_mult_218_n832, DP_mult_218_n831,
         DP_mult_218_n830, DP_mult_218_n829, DP_mult_218_n828,
         DP_mult_218_n827, DP_mult_218_n826, DP_mult_218_n825,
         DP_mult_218_n824, DP_mult_218_n823, DP_mult_218_n822,
         DP_mult_218_n821, DP_mult_218_n820, DP_mult_218_n819,
         DP_mult_218_n818, DP_mult_218_n817, DP_mult_218_n816,
         DP_mult_218_n815, DP_mult_218_n814, DP_mult_218_n813,
         DP_mult_218_n812, DP_mult_218_n811, DP_mult_218_n810,
         DP_mult_218_n809, DP_mult_218_n808, DP_mult_218_n807,
         DP_mult_218_n806, DP_mult_218_n805, DP_mult_218_n804,
         DP_mult_218_n803, DP_mult_218_n802, DP_mult_218_n801,
         DP_mult_218_n800, DP_mult_218_n799, DP_mult_218_n798,
         DP_mult_218_n797, DP_mult_218_n796, DP_mult_218_n795,
         DP_mult_218_n794, DP_mult_218_n793, DP_mult_218_n792,
         DP_mult_218_n791, DP_mult_218_n790, DP_mult_218_n789,
         DP_mult_218_n788, DP_mult_218_n787, DP_mult_218_n786,
         DP_mult_218_n785, DP_mult_218_n784, DP_mult_218_n783,
         DP_mult_218_n782, DP_mult_218_n781, DP_mult_218_n780,
         DP_mult_218_n779, DP_mult_218_n778, DP_mult_218_n777,
         DP_mult_218_n776, DP_mult_218_n775, DP_mult_218_n774,
         DP_mult_218_n773, DP_mult_218_n772, DP_mult_218_n771,
         DP_mult_218_n770, DP_mult_218_n769, DP_mult_218_n768,
         DP_mult_218_n767, DP_mult_218_n766, DP_mult_218_n765,
         DP_mult_218_n764, DP_mult_218_n763, DP_mult_218_n762,
         DP_mult_218_n761, DP_mult_218_n760, DP_mult_218_n759,
         DP_mult_218_n758, DP_mult_218_n757, DP_mult_218_n756,
         DP_mult_218_n755, DP_mult_218_n754, DP_mult_218_n753,
         DP_mult_218_n752, DP_mult_218_n751, DP_mult_218_n750,
         DP_mult_218_n749, DP_mult_218_n748, DP_mult_218_n747,
         DP_mult_218_n746, DP_mult_218_n745, DP_mult_218_n744,
         DP_mult_218_n743, DP_mult_218_n742, DP_mult_218_n741,
         DP_mult_218_n740, DP_mult_218_n739, DP_mult_218_n738,
         DP_mult_218_n737, DP_mult_218_n736, DP_mult_218_n735,
         DP_mult_218_n734, DP_mult_218_n733, DP_mult_218_n732,
         DP_mult_218_n731, DP_mult_218_n730, DP_mult_218_n729,
         DP_mult_218_n727, DP_mult_218_n726, DP_mult_218_n725,
         DP_mult_218_n724, DP_mult_218_n723, DP_mult_218_n722,
         DP_mult_218_n721, DP_mult_218_n720, DP_mult_218_n719,
         DP_mult_218_n718, DP_mult_218_n717, DP_mult_218_n716,
         DP_mult_218_n715, DP_mult_218_n714, DP_mult_218_n713,
         DP_mult_218_n712, DP_mult_218_n711, DP_mult_218_n710,
         DP_mult_218_n709, DP_mult_218_n708, DP_mult_218_n707,
         DP_mult_218_n706, DP_mult_218_n688, DP_mult_218_n687,
         DP_mult_218_n686, DP_mult_218_n685, DP_mult_218_n684,
         DP_mult_218_n683, DP_mult_218_n682, DP_mult_218_n681,
         DP_mult_218_n680, DP_mult_218_n679, DP_mult_218_n678,
         DP_mult_218_n677, DP_mult_218_n676, DP_mult_218_n675,
         DP_mult_218_n674, DP_mult_218_n673, DP_mult_218_n672,
         DP_mult_218_n671, DP_mult_218_n670, DP_mult_218_n669,
         DP_mult_218_n668, DP_mult_218_n667, DP_mult_218_n666,
         DP_mult_218_n665, DP_mult_218_n664, DP_mult_218_n663,
         DP_mult_218_n662, DP_mult_218_n661, DP_mult_218_n660,
         DP_mult_218_n659, DP_mult_218_n658, DP_mult_218_n657,
         DP_mult_218_n656, DP_mult_218_n655, DP_mult_218_n654,
         DP_mult_218_n653, DP_mult_218_n652, DP_mult_218_n651,
         DP_mult_218_n650, DP_mult_218_n649, DP_mult_218_n648,
         DP_mult_218_n647, DP_mult_218_n646, DP_mult_218_n645,
         DP_mult_218_n644, DP_mult_218_n643, DP_mult_218_n642,
         DP_mult_218_n641, DP_mult_218_n640, DP_mult_218_n639,
         DP_mult_218_n638, DP_mult_218_n637, DP_mult_218_n636,
         DP_mult_218_n635, DP_mult_218_n634, DP_mult_218_n633,
         DP_mult_218_n632, DP_mult_218_n631, DP_mult_218_n630,
         DP_mult_218_n629, DP_mult_218_n628, DP_mult_218_n627,
         DP_mult_218_n626, DP_mult_218_n625, DP_mult_218_n624,
         DP_mult_218_n623, DP_mult_218_n622, DP_mult_218_n621,
         DP_mult_218_n620, DP_mult_218_n619, DP_mult_218_n618,
         DP_mult_218_n617, DP_mult_218_n616, DP_mult_218_n615,
         DP_mult_218_n614, DP_mult_218_n613, DP_mult_218_n612,
         DP_mult_218_n611, DP_mult_218_n610, DP_mult_218_n609,
         DP_mult_218_n608, DP_mult_218_n607, DP_mult_218_n606,
         DP_mult_218_n605, DP_mult_218_n604, DP_mult_218_n603,
         DP_mult_218_n602, DP_mult_218_n601, DP_mult_218_n600,
         DP_mult_218_n599, DP_mult_218_n598, DP_mult_218_n597,
         DP_mult_218_n596, DP_mult_218_n595, DP_mult_218_n594,
         DP_mult_218_n593, DP_mult_218_n592, DP_mult_218_n591,
         DP_mult_218_n590, DP_mult_218_n589, DP_mult_218_n588,
         DP_mult_218_n587, DP_mult_218_n586, DP_mult_218_n585,
         DP_mult_218_n584, DP_mult_218_n583, DP_mult_218_n582,
         DP_mult_218_n581, DP_mult_218_n580, DP_mult_218_n579,
         DP_mult_218_n578, DP_mult_218_n577, DP_mult_218_n576,
         DP_mult_218_n575, DP_mult_218_n574, DP_mult_218_n573,
         DP_mult_218_n572, DP_mult_218_n571, DP_mult_218_n570,
         DP_mult_218_n569, DP_mult_218_n568, DP_mult_218_n567,
         DP_mult_218_n566, DP_mult_218_n565, DP_mult_218_n564,
         DP_mult_218_n563, DP_mult_218_n562, DP_mult_218_n561,
         DP_mult_218_n560, DP_mult_218_n559, DP_mult_218_n558,
         DP_mult_218_n557, DP_mult_218_n556, DP_mult_218_n555,
         DP_mult_218_n554, DP_mult_218_n553, DP_mult_218_n552,
         DP_mult_218_n551, DP_mult_218_n550, DP_mult_218_n549,
         DP_mult_218_n548, DP_mult_218_n547, DP_mult_218_n546,
         DP_mult_218_n545, DP_mult_218_n544, DP_mult_218_n543,
         DP_mult_218_n542, DP_mult_218_n541, DP_mult_218_n540,
         DP_mult_218_n539, DP_mult_218_n538, DP_mult_218_n537,
         DP_mult_218_n536, DP_mult_218_n535, DP_mult_218_n534,
         DP_mult_218_n533, DP_mult_218_n532, DP_mult_218_n531,
         DP_mult_218_n530, DP_mult_218_n529, DP_mult_218_n528,
         DP_mult_218_n527, DP_mult_218_n526, DP_mult_218_n525,
         DP_mult_218_n524, DP_mult_218_n523, DP_mult_218_n522,
         DP_mult_218_n521, DP_mult_218_n520, DP_mult_218_n519,
         DP_mult_218_n518, DP_mult_218_n517, DP_mult_218_n516,
         DP_mult_218_n515, DP_mult_218_n514, DP_mult_218_n513,
         DP_mult_218_n512, DP_mult_218_n511, DP_mult_218_n510,
         DP_mult_218_n509, DP_mult_218_n508, DP_mult_218_n507,
         DP_mult_218_n506, DP_mult_218_n505, DP_mult_218_n504,
         DP_mult_218_n503, DP_mult_218_n502, DP_mult_218_n501,
         DP_mult_218_n500, DP_mult_218_n499, DP_mult_218_n498,
         DP_mult_218_n497, DP_mult_218_n496, DP_mult_218_n495,
         DP_mult_218_n494, DP_mult_218_n493, DP_mult_218_n492,
         DP_mult_218_n491, DP_mult_218_n490, DP_mult_218_n489,
         DP_mult_218_n488, DP_mult_218_n487, DP_mult_218_n486,
         DP_mult_218_n485, DP_mult_218_n484, DP_mult_218_n483,
         DP_mult_218_n482, DP_mult_218_n481, DP_mult_218_n479,
         DP_mult_218_n478, DP_mult_218_n477, DP_mult_218_n476,
         DP_mult_218_n475, DP_mult_218_n474, DP_mult_218_n473,
         DP_mult_218_n472, DP_mult_218_n471, DP_mult_218_n470,
         DP_mult_218_n469, DP_mult_218_n468, DP_mult_218_n467,
         DP_mult_218_n466, DP_mult_218_n465, DP_mult_218_n464,
         DP_mult_218_n463, DP_mult_218_n462, DP_mult_218_n461,
         DP_mult_218_n460, DP_mult_218_n459, DP_mult_218_n458,
         DP_mult_218_n457, DP_mult_218_n456, DP_mult_218_n455,
         DP_mult_218_n454, DP_mult_218_n453, DP_mult_218_n452,
         DP_mult_218_n451, DP_mult_218_n450, DP_mult_218_n449,
         DP_mult_218_n448, DP_mult_218_n447, DP_mult_218_n446,
         DP_mult_218_n445, DP_mult_218_n444, DP_mult_218_n442,
         DP_mult_218_n441, DP_mult_218_n440, DP_mult_218_n439,
         DP_mult_218_n438, DP_mult_218_n437, DP_mult_218_n436,
         DP_mult_218_n435, DP_mult_218_n434, DP_mult_218_n433,
         DP_mult_218_n432, DP_mult_218_n431, DP_mult_218_n430,
         DP_mult_218_n429, DP_mult_218_n428, DP_mult_218_n427,
         DP_mult_218_n426, DP_mult_218_n425, DP_mult_218_n424,
         DP_mult_218_n423, DP_mult_218_n422, DP_mult_218_n421,
         DP_mult_218_n420, DP_mult_218_n419, DP_mult_218_n418,
         DP_mult_218_n417, DP_mult_218_n416, DP_mult_218_n415,
         DP_mult_218_n414, DP_mult_218_n413, DP_mult_218_n411,
         DP_mult_218_n410, DP_mult_218_n409, DP_mult_218_n408,
         DP_mult_218_n407, DP_mult_218_n406, DP_mult_218_n405,
         DP_mult_218_n404, DP_mult_218_n403, DP_mult_218_n402,
         DP_mult_218_n401, DP_mult_218_n400, DP_mult_218_n399,
         DP_mult_218_n398, DP_mult_218_n397, DP_mult_218_n396,
         DP_mult_218_n395, DP_mult_218_n394, DP_mult_218_n393,
         DP_mult_218_n392, DP_mult_218_n391, DP_mult_218_n390,
         DP_mult_218_n389, DP_mult_218_n387, DP_mult_218_n386,
         DP_mult_218_n385, DP_mult_218_n384, DP_mult_218_n383,
         DP_mult_218_n382, DP_mult_218_n381, DP_mult_218_n380,
         DP_mult_218_n379, DP_mult_218_n378, DP_mult_218_n377,
         DP_mult_218_n376, DP_mult_218_n375, DP_mult_218_n374,
         DP_mult_218_n373, DP_mult_218_n372, DP_mult_218_n371,
         DP_mult_218_n370, DP_mult_218_n368, DP_mult_218_n367,
         DP_mult_218_n366, DP_mult_218_n365, DP_mult_218_n364,
         DP_mult_218_n363, DP_mult_218_n362, DP_mult_218_n361,
         DP_mult_218_n360, DP_mult_218_n359, DP_mult_218_n358,
         DP_mult_218_n356, DP_mult_218_n355, DP_mult_218_n354,
         DP_mult_218_n353, DP_mult_218_n352, DP_mult_218_n351,
         DP_mult_218_n326, DP_mult_218_n325, DP_mult_218_n324,
         DP_mult_218_n323, DP_mult_218_n322, DP_mult_218_n321,
         DP_mult_218_n320, DP_mult_218_n319, DP_mult_218_n318,
         DP_mult_218_n317, DP_mult_218_n316, DP_mult_218_n315,
         DP_mult_218_n314, DP_mult_218_n313, DP_mult_218_n312,
         DP_mult_218_n311, DP_mult_218_n310, DP_mult_218_n309,
         DP_mult_218_n308, DP_mult_218_n307, DP_mult_218_n306,
         DP_mult_218_n305, DP_mult_218_n304, DP_mult_218_n303,
         DP_mult_217_n2162, DP_mult_217_n2161, DP_mult_217_n2160,
         DP_mult_217_n2159, DP_mult_217_n2158, DP_mult_217_n2157,
         DP_mult_217_n2156, DP_mult_217_n2155, DP_mult_217_n2154,
         DP_mult_217_n2153, DP_mult_217_n2152, DP_mult_217_n2151,
         DP_mult_217_n2150, DP_mult_217_n2149, DP_mult_217_n2148,
         DP_mult_217_n2147, DP_mult_217_n2146, DP_mult_217_n2145,
         DP_mult_217_n2144, DP_mult_217_n2143, DP_mult_217_n2142,
         DP_mult_217_n2141, DP_mult_217_n2140, DP_mult_217_n2139,
         DP_mult_217_n2138, DP_mult_217_n2137, DP_mult_217_n2136,
         DP_mult_217_n2135, DP_mult_217_n2134, DP_mult_217_n2133,
         DP_mult_217_n2132, DP_mult_217_n2131, DP_mult_217_n2130,
         DP_mult_217_n2129, DP_mult_217_n2128, DP_mult_217_n2127,
         DP_mult_217_n2126, DP_mult_217_n2125, DP_mult_217_n2124,
         DP_mult_217_n2123, DP_mult_217_n2122, DP_mult_217_n2121,
         DP_mult_217_n2120, DP_mult_217_n2119, DP_mult_217_n2118,
         DP_mult_217_n2117, DP_mult_217_n2116, DP_mult_217_n2115,
         DP_mult_217_n2114, DP_mult_217_n2113, DP_mult_217_n2112,
         DP_mult_217_n2111, DP_mult_217_n2110, DP_mult_217_n2109,
         DP_mult_217_n2108, DP_mult_217_n2107, DP_mult_217_n2106,
         DP_mult_217_n2105, DP_mult_217_n2104, DP_mult_217_n2103,
         DP_mult_217_n2102, DP_mult_217_n2101, DP_mult_217_n2100,
         DP_mult_217_n2099, DP_mult_217_n2098, DP_mult_217_n2097,
         DP_mult_217_n2096, DP_mult_217_n2095, DP_mult_217_n2094,
         DP_mult_217_n2093, DP_mult_217_n2092, DP_mult_217_n2091,
         DP_mult_217_n2090, DP_mult_217_n2089, DP_mult_217_n2088,
         DP_mult_217_n2087, DP_mult_217_n2086, DP_mult_217_n2085,
         DP_mult_217_n2084, DP_mult_217_n2083, DP_mult_217_n2082,
         DP_mult_217_n2081, DP_mult_217_n2080, DP_mult_217_n2079,
         DP_mult_217_n2078, DP_mult_217_n2077, DP_mult_217_n2076,
         DP_mult_217_n2075, DP_mult_217_n2074, DP_mult_217_n2073,
         DP_mult_217_n2072, DP_mult_217_n2071, DP_mult_217_n2070,
         DP_mult_217_n2069, DP_mult_217_n2068, DP_mult_217_n2067,
         DP_mult_217_n2066, DP_mult_217_n2065, DP_mult_217_n2064,
         DP_mult_217_n2063, DP_mult_217_n2062, DP_mult_217_n2061,
         DP_mult_217_n2060, DP_mult_217_n2059, DP_mult_217_n2058,
         DP_mult_217_n2057, DP_mult_217_n2056, DP_mult_217_n2055,
         DP_mult_217_n2054, DP_mult_217_n2053, DP_mult_217_n2052,
         DP_mult_217_n2051, DP_mult_217_n2050, DP_mult_217_n2049,
         DP_mult_217_n2048, DP_mult_217_n2047, DP_mult_217_n2046,
         DP_mult_217_n2045, DP_mult_217_n2044, DP_mult_217_n2043,
         DP_mult_217_n2042, DP_mult_217_n2041, DP_mult_217_n2040,
         DP_mult_217_n2039, DP_mult_217_n2038, DP_mult_217_n2037,
         DP_mult_217_n2036, DP_mult_217_n2035, DP_mult_217_n2034,
         DP_mult_217_n2033, DP_mult_217_n2032, DP_mult_217_n2031,
         DP_mult_217_n2030, DP_mult_217_n2029, DP_mult_217_n2028,
         DP_mult_217_n2027, DP_mult_217_n2026, DP_mult_217_n2025,
         DP_mult_217_n2024, DP_mult_217_n2023, DP_mult_217_n2022,
         DP_mult_217_n2021, DP_mult_217_n2020, DP_mult_217_n2019,
         DP_mult_217_n2018, DP_mult_217_n2017, DP_mult_217_n2016,
         DP_mult_217_n2015, DP_mult_217_n2014, DP_mult_217_n2013,
         DP_mult_217_n2012, DP_mult_217_n2011, DP_mult_217_n2010,
         DP_mult_217_n2009, DP_mult_217_n2008, DP_mult_217_n2007,
         DP_mult_217_n2006, DP_mult_217_n2005, DP_mult_217_n2004,
         DP_mult_217_n2003, DP_mult_217_n2002, DP_mult_217_n2001,
         DP_mult_217_n2000, DP_mult_217_n1999, DP_mult_217_n1998,
         DP_mult_217_n1997, DP_mult_217_n1996, DP_mult_217_n1995,
         DP_mult_217_n1994, DP_mult_217_n1993, DP_mult_217_n1992,
         DP_mult_217_n1991, DP_mult_217_n1990, DP_mult_217_n1989,
         DP_mult_217_n1988, DP_mult_217_n1987, DP_mult_217_n1986,
         DP_mult_217_n1985, DP_mult_217_n1984, DP_mult_217_n1983,
         DP_mult_217_n1982, DP_mult_217_n1981, DP_mult_217_n1980,
         DP_mult_217_n1979, DP_mult_217_n1978, DP_mult_217_n1977,
         DP_mult_217_n1976, DP_mult_217_n1975, DP_mult_217_n1974,
         DP_mult_217_n1973, DP_mult_217_n1972, DP_mult_217_n1971,
         DP_mult_217_n1970, DP_mult_217_n1969, DP_mult_217_n1968,
         DP_mult_217_n1967, DP_mult_217_n1966, DP_mult_217_n1965,
         DP_mult_217_n1964, DP_mult_217_n1963, DP_mult_217_n1962,
         DP_mult_217_n1961, DP_mult_217_n1960, DP_mult_217_n1959,
         DP_mult_217_n1958, DP_mult_217_n1957, DP_mult_217_n1956,
         DP_mult_217_n1955, DP_mult_217_n1954, DP_mult_217_n1953,
         DP_mult_217_n1952, DP_mult_217_n1951, DP_mult_217_n1950,
         DP_mult_217_n1949, DP_mult_217_n1948, DP_mult_217_n1947,
         DP_mult_217_n1946, DP_mult_217_n1945, DP_mult_217_n1944,
         DP_mult_217_n1943, DP_mult_217_n1942, DP_mult_217_n1941,
         DP_mult_217_n1940, DP_mult_217_n1939, DP_mult_217_n1938,
         DP_mult_217_n1937, DP_mult_217_n1936, DP_mult_217_n1935,
         DP_mult_217_n1934, DP_mult_217_n1933, DP_mult_217_n1932,
         DP_mult_217_n1931, DP_mult_217_n1930, DP_mult_217_n1929,
         DP_mult_217_n1928, DP_mult_217_n1927, DP_mult_217_n1926,
         DP_mult_217_n1925, DP_mult_217_n1924, DP_mult_217_n1923,
         DP_mult_217_n1922, DP_mult_217_n1921, DP_mult_217_n1920,
         DP_mult_217_n1919, DP_mult_217_n1918, DP_mult_217_n1917,
         DP_mult_217_n1916, DP_mult_217_n1915, DP_mult_217_n1914,
         DP_mult_217_n1913, DP_mult_217_n1912, DP_mult_217_n1911,
         DP_mult_217_n1910, DP_mult_217_n1909, DP_mult_217_n1908,
         DP_mult_217_n1907, DP_mult_217_n1906, DP_mult_217_n1905,
         DP_mult_217_n1904, DP_mult_217_n1903, DP_mult_217_n1902,
         DP_mult_217_n1901, DP_mult_217_n1900, DP_mult_217_n1899,
         DP_mult_217_n1898, DP_mult_217_n1897, DP_mult_217_n1896,
         DP_mult_217_n1895, DP_mult_217_n1894, DP_mult_217_n1893,
         DP_mult_217_n1892, DP_mult_217_n1891, DP_mult_217_n1890,
         DP_mult_217_n1889, DP_mult_217_n1888, DP_mult_217_n1887,
         DP_mult_217_n1886, DP_mult_217_n1885, DP_mult_217_n1884,
         DP_mult_217_n1883, DP_mult_217_n1882, DP_mult_217_n1881,
         DP_mult_217_n1880, DP_mult_217_n1879, DP_mult_217_n1878,
         DP_mult_217_n1877, DP_mult_217_n1876, DP_mult_217_n1875,
         DP_mult_217_n1874, DP_mult_217_n1873, DP_mult_217_n1872,
         DP_mult_217_n1871, DP_mult_217_n1870, DP_mult_217_n1869,
         DP_mult_217_n1868, DP_mult_217_n1867, DP_mult_217_n1866,
         DP_mult_217_n1865, DP_mult_217_n1864, DP_mult_217_n1863,
         DP_mult_217_n1862, DP_mult_217_n1861, DP_mult_217_n1860,
         DP_mult_217_n1859, DP_mult_217_n1858, DP_mult_217_n1857,
         DP_mult_217_n1856, DP_mult_217_n1855, DP_mult_217_n1854,
         DP_mult_217_n1853, DP_mult_217_n1852, DP_mult_217_n1851,
         DP_mult_217_n1850, DP_mult_217_n1849, DP_mult_217_n1848,
         DP_mult_217_n1847, DP_mult_217_n1846, DP_mult_217_n1845,
         DP_mult_217_n1844, DP_mult_217_n1843, DP_mult_217_n1842,
         DP_mult_217_n1841, DP_mult_217_n1840, DP_mult_217_n1839,
         DP_mult_217_n1838, DP_mult_217_n1837, DP_mult_217_n1836,
         DP_mult_217_n1835, DP_mult_217_n1834, DP_mult_217_n1833,
         DP_mult_217_n1832, DP_mult_217_n1831, DP_mult_217_n1830,
         DP_mult_217_n1829, DP_mult_217_n1828, DP_mult_217_n1827,
         DP_mult_217_n1826, DP_mult_217_n1825, DP_mult_217_n1824,
         DP_mult_217_n1823, DP_mult_217_n1822, DP_mult_217_n1821,
         DP_mult_217_n1820, DP_mult_217_n1819, DP_mult_217_n1818,
         DP_mult_217_n1817, DP_mult_217_n1816, DP_mult_217_n1815,
         DP_mult_217_n1814, DP_mult_217_n1813, DP_mult_217_n1812,
         DP_mult_217_n1811, DP_mult_217_n1810, DP_mult_217_n1809,
         DP_mult_217_n1808, DP_mult_217_n1807, DP_mult_217_n1806,
         DP_mult_217_n1805, DP_mult_217_n1804, DP_mult_217_n1803,
         DP_mult_217_n1802, DP_mult_217_n1801, DP_mult_217_n1800,
         DP_mult_217_n1799, DP_mult_217_n1798, DP_mult_217_n1797,
         DP_mult_217_n1796, DP_mult_217_n1795, DP_mult_217_n1794,
         DP_mult_217_n1793, DP_mult_217_n1792, DP_mult_217_n1791,
         DP_mult_217_n1790, DP_mult_217_n1789, DP_mult_217_n1788,
         DP_mult_217_n1787, DP_mult_217_n1786, DP_mult_217_n1785,
         DP_mult_217_n1784, DP_mult_217_n1783, DP_mult_217_n1782,
         DP_mult_217_n1781, DP_mult_217_n1780, DP_mult_217_n1779,
         DP_mult_217_n1778, DP_mult_217_n1777, DP_mult_217_n1776,
         DP_mult_217_n1775, DP_mult_217_n1774, DP_mult_217_n1773,
         DP_mult_217_n1772, DP_mult_217_n1771, DP_mult_217_n1770,
         DP_mult_217_n1769, DP_mult_217_n1768, DP_mult_217_n1767,
         DP_mult_217_n1766, DP_mult_217_n1765, DP_mult_217_n1764,
         DP_mult_217_n1763, DP_mult_217_n1762, DP_mult_217_n1761,
         DP_mult_217_n1760, DP_mult_217_n1759, DP_mult_217_n1758,
         DP_mult_217_n1757, DP_mult_217_n1756, DP_mult_217_n1755,
         DP_mult_217_n1754, DP_mult_217_n1753, DP_mult_217_n1752,
         DP_mult_217_n1751, DP_mult_217_n1750, DP_mult_217_n1749,
         DP_mult_217_n1748, DP_mult_217_n1747, DP_mult_217_n1746,
         DP_mult_217_n1745, DP_mult_217_n1744, DP_mult_217_n1743,
         DP_mult_217_n1742, DP_mult_217_n1741, DP_mult_217_n1740,
         DP_mult_217_n1739, DP_mult_217_n1738, DP_mult_217_n1737,
         DP_mult_217_n1736, DP_mult_217_n1735, DP_mult_217_n1734,
         DP_mult_217_n1733, DP_mult_217_n1732, DP_mult_217_n1731,
         DP_mult_217_n1730, DP_mult_217_n1729, DP_mult_217_n1728,
         DP_mult_217_n1727, DP_mult_217_n1726, DP_mult_217_n1725,
         DP_mult_217_n1724, DP_mult_217_n1723, DP_mult_217_n1722,
         DP_mult_217_n1721, DP_mult_217_n1720, DP_mult_217_n1719,
         DP_mult_217_n1718, DP_mult_217_n1717, DP_mult_217_n1716,
         DP_mult_217_n1715, DP_mult_217_n1714, DP_mult_217_n1713,
         DP_mult_217_n1712, DP_mult_217_n1711, DP_mult_217_n1710,
         DP_mult_217_n1709, DP_mult_217_n1708, DP_mult_217_n1707,
         DP_mult_217_n1706, DP_mult_217_n1705, DP_mult_217_n1704,
         DP_mult_217_n1703, DP_mult_217_n1702, DP_mult_217_n1701,
         DP_mult_217_n1700, DP_mult_217_n1699, DP_mult_217_n1698,
         DP_mult_217_n1697, DP_mult_217_n1696, DP_mult_217_n1695,
         DP_mult_217_n1694, DP_mult_217_n1693, DP_mult_217_n1692,
         DP_mult_217_n1691, DP_mult_217_n1690, DP_mult_217_n1689,
         DP_mult_217_n1688, DP_mult_217_n1687, DP_mult_217_n1686,
         DP_mult_217_n1685, DP_mult_217_n1684, DP_mult_217_n1683,
         DP_mult_217_n1682, DP_mult_217_n1681, DP_mult_217_n1680,
         DP_mult_217_n1679, DP_mult_217_n1678, DP_mult_217_n1677,
         DP_mult_217_n1676, DP_mult_217_n1675, DP_mult_217_n1674,
         DP_mult_217_n1673, DP_mult_217_n1672, DP_mult_217_n1671,
         DP_mult_217_n1670, DP_mult_217_n1669, DP_mult_217_n1668,
         DP_mult_217_n1667, DP_mult_217_n1666, DP_mult_217_n1665,
         DP_mult_217_n1664, DP_mult_217_n1663, DP_mult_217_n1662,
         DP_mult_217_n1661, DP_mult_217_n1660, DP_mult_217_n1659,
         DP_mult_217_n1658, DP_mult_217_n1657, DP_mult_217_n1656,
         DP_mult_217_n1655, DP_mult_217_n1654, DP_mult_217_n1653,
         DP_mult_217_n1652, DP_mult_217_n1651, DP_mult_217_n1650,
         DP_mult_217_n1649, DP_mult_217_n1648, DP_mult_217_n1647,
         DP_mult_217_n1646, DP_mult_217_n1645, DP_mult_217_n1644,
         DP_mult_217_n1643, DP_mult_217_n1642, DP_mult_217_n1641,
         DP_mult_217_n1640, DP_mult_217_n1639, DP_mult_217_n1638,
         DP_mult_217_n1637, DP_mult_217_n1636, DP_mult_217_n1635,
         DP_mult_217_n1634, DP_mult_217_n1633, DP_mult_217_n1632,
         DP_mult_217_n1631, DP_mult_217_n1630, DP_mult_217_n1629,
         DP_mult_217_n1628, DP_mult_217_n1627, DP_mult_217_n1626,
         DP_mult_217_n1625, DP_mult_217_n1624, DP_mult_217_n1623,
         DP_mult_217_n1622, DP_mult_217_n1621, DP_mult_217_n1620,
         DP_mult_217_n1619, DP_mult_217_n1618, DP_mult_217_n1617,
         DP_mult_217_n1616, DP_mult_217_n1615, DP_mult_217_n1614,
         DP_mult_217_n1613, DP_mult_217_n1612, DP_mult_217_n1611,
         DP_mult_217_n1610, DP_mult_217_n1609, DP_mult_217_n1608,
         DP_mult_217_n1607, DP_mult_217_n1606, DP_mult_217_n1605,
         DP_mult_217_n1604, DP_mult_217_n1603, DP_mult_217_n1602,
         DP_mult_217_n1601, DP_mult_217_n1600, DP_mult_217_n1599,
         DP_mult_217_n1598, DP_mult_217_n1597, DP_mult_217_n1596,
         DP_mult_217_n1595, DP_mult_217_n1594, DP_mult_217_n1593,
         DP_mult_217_n1592, DP_mult_217_n1591, DP_mult_217_n1590,
         DP_mult_217_n1589, DP_mult_217_n1588, DP_mult_217_n1587,
         DP_mult_217_n1586, DP_mult_217_n1585, DP_mult_217_n1584,
         DP_mult_217_n1583, DP_mult_217_n1582, DP_mult_217_n1581,
         DP_mult_217_n1580, DP_mult_217_n1579, DP_mult_217_n1578,
         DP_mult_217_n1577, DP_mult_217_n1576, DP_mult_217_n1575,
         DP_mult_217_n1574, DP_mult_217_n1573, DP_mult_217_n1572,
         DP_mult_217_n1571, DP_mult_217_n1570, DP_mult_217_n1569,
         DP_mult_217_n1568, DP_mult_217_n1567, DP_mult_217_n1566,
         DP_mult_217_n1565, DP_mult_217_n1564, DP_mult_217_n1563,
         DP_mult_217_n1562, DP_mult_217_n1561, DP_mult_217_n1560,
         DP_mult_217_n1559, DP_mult_217_n1558, DP_mult_217_n1557,
         DP_mult_217_n1556, DP_mult_217_n1555, DP_mult_217_n1554,
         DP_mult_217_n1553, DP_mult_217_n1552, DP_mult_217_n1551,
         DP_mult_217_n1550, DP_mult_217_n1549, DP_mult_217_n1548,
         DP_mult_217_n1547, DP_mult_217_n1546, DP_mult_217_n1545,
         DP_mult_217_n1544, DP_mult_217_n1543, DP_mult_217_n1542,
         DP_mult_217_n1541, DP_mult_217_n1540, DP_mult_217_n1539,
         DP_mult_217_n1538, DP_mult_217_n1537, DP_mult_217_n1536,
         DP_mult_217_n1535, DP_mult_217_n1534, DP_mult_217_n1533,
         DP_mult_217_n1397, DP_mult_217_n1396, DP_mult_217_n1395,
         DP_mult_217_n1394, DP_mult_217_n1393, DP_mult_217_n1392,
         DP_mult_217_n1391, DP_mult_217_n1390, DP_mult_217_n1389,
         DP_mult_217_n1388, DP_mult_217_n1387, DP_mult_217_n1386,
         DP_mult_217_n1385, DP_mult_217_n1384, DP_mult_217_n1383,
         DP_mult_217_n1382, DP_mult_217_n1381, DP_mult_217_n1380,
         DP_mult_217_n1379, DP_mult_217_n1378, DP_mult_217_n1377,
         DP_mult_217_n1376, DP_mult_217_n1375, DP_mult_217_n1374,
         DP_mult_217_n908, DP_mult_217_n907, DP_mult_217_n906,
         DP_mult_217_n904, DP_mult_217_n903, DP_mult_217_n902,
         DP_mult_217_n901, DP_mult_217_n900, DP_mult_217_n899,
         DP_mult_217_n898, DP_mult_217_n897, DP_mult_217_n896,
         DP_mult_217_n895, DP_mult_217_n894, DP_mult_217_n893,
         DP_mult_217_n892, DP_mult_217_n891, DP_mult_217_n890,
         DP_mult_217_n889, DP_mult_217_n888, DP_mult_217_n887,
         DP_mult_217_n886, DP_mult_217_n885, DP_mult_217_n884,
         DP_mult_217_n883, DP_mult_217_n882, DP_mult_217_n881,
         DP_mult_217_n880, DP_mult_217_n879, DP_mult_217_n878,
         DP_mult_217_n877, DP_mult_217_n876, DP_mult_217_n875,
         DP_mult_217_n874, DP_mult_217_n873, DP_mult_217_n872,
         DP_mult_217_n871, DP_mult_217_n870, DP_mult_217_n869,
         DP_mult_217_n868, DP_mult_217_n867, DP_mult_217_n866,
         DP_mult_217_n865, DP_mult_217_n864, DP_mult_217_n863,
         DP_mult_217_n862, DP_mult_217_n861, DP_mult_217_n860,
         DP_mult_217_n859, DP_mult_217_n858, DP_mult_217_n857,
         DP_mult_217_n856, DP_mult_217_n855, DP_mult_217_n854,
         DP_mult_217_n853, DP_mult_217_n852, DP_mult_217_n851,
         DP_mult_217_n850, DP_mult_217_n849, DP_mult_217_n848,
         DP_mult_217_n847, DP_mult_217_n846, DP_mult_217_n845,
         DP_mult_217_n844, DP_mult_217_n843, DP_mult_217_n842,
         DP_mult_217_n841, DP_mult_217_n840, DP_mult_217_n839,
         DP_mult_217_n838, DP_mult_217_n837, DP_mult_217_n836,
         DP_mult_217_n835, DP_mult_217_n834, DP_mult_217_n833,
         DP_mult_217_n832, DP_mult_217_n831, DP_mult_217_n830,
         DP_mult_217_n829, DP_mult_217_n828, DP_mult_217_n827,
         DP_mult_217_n826, DP_mult_217_n825, DP_mult_217_n824,
         DP_mult_217_n823, DP_mult_217_n822, DP_mult_217_n821,
         DP_mult_217_n820, DP_mult_217_n819, DP_mult_217_n818,
         DP_mult_217_n817, DP_mult_217_n816, DP_mult_217_n815,
         DP_mult_217_n814, DP_mult_217_n813, DP_mult_217_n812,
         DP_mult_217_n811, DP_mult_217_n810, DP_mult_217_n809,
         DP_mult_217_n808, DP_mult_217_n807, DP_mult_217_n806,
         DP_mult_217_n805, DP_mult_217_n804, DP_mult_217_n803,
         DP_mult_217_n802, DP_mult_217_n801, DP_mult_217_n800,
         DP_mult_217_n799, DP_mult_217_n798, DP_mult_217_n797,
         DP_mult_217_n796, DP_mult_217_n795, DP_mult_217_n794,
         DP_mult_217_n793, DP_mult_217_n792, DP_mult_217_n791,
         DP_mult_217_n790, DP_mult_217_n789, DP_mult_217_n788,
         DP_mult_217_n787, DP_mult_217_n786, DP_mult_217_n785,
         DP_mult_217_n784, DP_mult_217_n783, DP_mult_217_n782,
         DP_mult_217_n781, DP_mult_217_n780, DP_mult_217_n779,
         DP_mult_217_n778, DP_mult_217_n777, DP_mult_217_n776,
         DP_mult_217_n775, DP_mult_217_n774, DP_mult_217_n773,
         DP_mult_217_n772, DP_mult_217_n771, DP_mult_217_n770,
         DP_mult_217_n769, DP_mult_217_n768, DP_mult_217_n767,
         DP_mult_217_n766, DP_mult_217_n765, DP_mult_217_n764,
         DP_mult_217_n763, DP_mult_217_n762, DP_mult_217_n761,
         DP_mult_217_n760, DP_mult_217_n759, DP_mult_217_n758,
         DP_mult_217_n757, DP_mult_217_n756, DP_mult_217_n755,
         DP_mult_217_n754, DP_mult_217_n753, DP_mult_217_n752,
         DP_mult_217_n751, DP_mult_217_n750, DP_mult_217_n749,
         DP_mult_217_n748, DP_mult_217_n747, DP_mult_217_n746,
         DP_mult_217_n745, DP_mult_217_n744, DP_mult_217_n743,
         DP_mult_217_n742, DP_mult_217_n741, DP_mult_217_n740,
         DP_mult_217_n739, DP_mult_217_n738, DP_mult_217_n737,
         DP_mult_217_n736, DP_mult_217_n735, DP_mult_217_n734,
         DP_mult_217_n733, DP_mult_217_n732, DP_mult_217_n731,
         DP_mult_217_n730, DP_mult_217_n729, DP_mult_217_n727,
         DP_mult_217_n726, DP_mult_217_n725, DP_mult_217_n724,
         DP_mult_217_n723, DP_mult_217_n722, DP_mult_217_n721,
         DP_mult_217_n720, DP_mult_217_n719, DP_mult_217_n718,
         DP_mult_217_n717, DP_mult_217_n716, DP_mult_217_n715,
         DP_mult_217_n714, DP_mult_217_n713, DP_mult_217_n712,
         DP_mult_217_n711, DP_mult_217_n710, DP_mult_217_n709,
         DP_mult_217_n708, DP_mult_217_n707, DP_mult_217_n706,
         DP_mult_217_n688, DP_mult_217_n687, DP_mult_217_n686,
         DP_mult_217_n685, DP_mult_217_n684, DP_mult_217_n683,
         DP_mult_217_n682, DP_mult_217_n681, DP_mult_217_n680,
         DP_mult_217_n679, DP_mult_217_n678, DP_mult_217_n677,
         DP_mult_217_n676, DP_mult_217_n675, DP_mult_217_n674,
         DP_mult_217_n673, DP_mult_217_n672, DP_mult_217_n671,
         DP_mult_217_n670, DP_mult_217_n669, DP_mult_217_n668,
         DP_mult_217_n667, DP_mult_217_n666, DP_mult_217_n665,
         DP_mult_217_n664, DP_mult_217_n663, DP_mult_217_n662,
         DP_mult_217_n661, DP_mult_217_n660, DP_mult_217_n659,
         DP_mult_217_n658, DP_mult_217_n657, DP_mult_217_n656,
         DP_mult_217_n655, DP_mult_217_n654, DP_mult_217_n653,
         DP_mult_217_n652, DP_mult_217_n651, DP_mult_217_n650,
         DP_mult_217_n649, DP_mult_217_n648, DP_mult_217_n647,
         DP_mult_217_n646, DP_mult_217_n645, DP_mult_217_n644,
         DP_mult_217_n643, DP_mult_217_n642, DP_mult_217_n641,
         DP_mult_217_n640, DP_mult_217_n639, DP_mult_217_n638,
         DP_mult_217_n637, DP_mult_217_n636, DP_mult_217_n635,
         DP_mult_217_n634, DP_mult_217_n633, DP_mult_217_n632,
         DP_mult_217_n631, DP_mult_217_n630, DP_mult_217_n629,
         DP_mult_217_n628, DP_mult_217_n627, DP_mult_217_n626,
         DP_mult_217_n625, DP_mult_217_n624, DP_mult_217_n623,
         DP_mult_217_n622, DP_mult_217_n621, DP_mult_217_n620,
         DP_mult_217_n619, DP_mult_217_n618, DP_mult_217_n617,
         DP_mult_217_n616, DP_mult_217_n615, DP_mult_217_n614,
         DP_mult_217_n613, DP_mult_217_n612, DP_mult_217_n611,
         DP_mult_217_n610, DP_mult_217_n609, DP_mult_217_n608,
         DP_mult_217_n607, DP_mult_217_n606, DP_mult_217_n605,
         DP_mult_217_n604, DP_mult_217_n603, DP_mult_217_n602,
         DP_mult_217_n601, DP_mult_217_n600, DP_mult_217_n599,
         DP_mult_217_n598, DP_mult_217_n597, DP_mult_217_n596,
         DP_mult_217_n595, DP_mult_217_n594, DP_mult_217_n593,
         DP_mult_217_n592, DP_mult_217_n591, DP_mult_217_n590,
         DP_mult_217_n589, DP_mult_217_n588, DP_mult_217_n587,
         DP_mult_217_n586, DP_mult_217_n585, DP_mult_217_n584,
         DP_mult_217_n583, DP_mult_217_n582, DP_mult_217_n581,
         DP_mult_217_n580, DP_mult_217_n579, DP_mult_217_n578,
         DP_mult_217_n577, DP_mult_217_n576, DP_mult_217_n575,
         DP_mult_217_n574, DP_mult_217_n573, DP_mult_217_n572,
         DP_mult_217_n571, DP_mult_217_n570, DP_mult_217_n569,
         DP_mult_217_n568, DP_mult_217_n567, DP_mult_217_n566,
         DP_mult_217_n565, DP_mult_217_n564, DP_mult_217_n563,
         DP_mult_217_n562, DP_mult_217_n561, DP_mult_217_n560,
         DP_mult_217_n559, DP_mult_217_n558, DP_mult_217_n557,
         DP_mult_217_n556, DP_mult_217_n555, DP_mult_217_n554,
         DP_mult_217_n553, DP_mult_217_n552, DP_mult_217_n551,
         DP_mult_217_n550, DP_mult_217_n549, DP_mult_217_n548,
         DP_mult_217_n547, DP_mult_217_n546, DP_mult_217_n545,
         DP_mult_217_n544, DP_mult_217_n543, DP_mult_217_n542,
         DP_mult_217_n541, DP_mult_217_n540, DP_mult_217_n539,
         DP_mult_217_n538, DP_mult_217_n537, DP_mult_217_n536,
         DP_mult_217_n535, DP_mult_217_n534, DP_mult_217_n533,
         DP_mult_217_n532, DP_mult_217_n531, DP_mult_217_n530,
         DP_mult_217_n529, DP_mult_217_n528, DP_mult_217_n527,
         DP_mult_217_n526, DP_mult_217_n525, DP_mult_217_n524,
         DP_mult_217_n523, DP_mult_217_n522, DP_mult_217_n521,
         DP_mult_217_n520, DP_mult_217_n519, DP_mult_217_n518,
         DP_mult_217_n517, DP_mult_217_n516, DP_mult_217_n515,
         DP_mult_217_n514, DP_mult_217_n513, DP_mult_217_n512,
         DP_mult_217_n511, DP_mult_217_n510, DP_mult_217_n509,
         DP_mult_217_n508, DP_mult_217_n507, DP_mult_217_n506,
         DP_mult_217_n505, DP_mult_217_n504, DP_mult_217_n503,
         DP_mult_217_n502, DP_mult_217_n501, DP_mult_217_n500,
         DP_mult_217_n499, DP_mult_217_n498, DP_mult_217_n497,
         DP_mult_217_n496, DP_mult_217_n495, DP_mult_217_n494,
         DP_mult_217_n493, DP_mult_217_n492, DP_mult_217_n491,
         DP_mult_217_n490, DP_mult_217_n489, DP_mult_217_n488,
         DP_mult_217_n487, DP_mult_217_n486, DP_mult_217_n485,
         DP_mult_217_n484, DP_mult_217_n483, DP_mult_217_n482,
         DP_mult_217_n481, DP_mult_217_n479, DP_mult_217_n478,
         DP_mult_217_n477, DP_mult_217_n476, DP_mult_217_n475,
         DP_mult_217_n474, DP_mult_217_n473, DP_mult_217_n472,
         DP_mult_217_n471, DP_mult_217_n470, DP_mult_217_n469,
         DP_mult_217_n468, DP_mult_217_n467, DP_mult_217_n466,
         DP_mult_217_n465, DP_mult_217_n464, DP_mult_217_n463,
         DP_mult_217_n462, DP_mult_217_n461, DP_mult_217_n460,
         DP_mult_217_n459, DP_mult_217_n458, DP_mult_217_n457,
         DP_mult_217_n456, DP_mult_217_n455, DP_mult_217_n454,
         DP_mult_217_n453, DP_mult_217_n452, DP_mult_217_n451,
         DP_mult_217_n450, DP_mult_217_n449, DP_mult_217_n448,
         DP_mult_217_n447, DP_mult_217_n446, DP_mult_217_n445,
         DP_mult_217_n444, DP_mult_217_n442, DP_mult_217_n441,
         DP_mult_217_n440, DP_mult_217_n439, DP_mult_217_n438,
         DP_mult_217_n437, DP_mult_217_n436, DP_mult_217_n435,
         DP_mult_217_n434, DP_mult_217_n433, DP_mult_217_n432,
         DP_mult_217_n431, DP_mult_217_n430, DP_mult_217_n429,
         DP_mult_217_n428, DP_mult_217_n427, DP_mult_217_n426,
         DP_mult_217_n425, DP_mult_217_n424, DP_mult_217_n423,
         DP_mult_217_n422, DP_mult_217_n421, DP_mult_217_n420,
         DP_mult_217_n419, DP_mult_217_n418, DP_mult_217_n417,
         DP_mult_217_n416, DP_mult_217_n415, DP_mult_217_n414,
         DP_mult_217_n413, DP_mult_217_n411, DP_mult_217_n410,
         DP_mult_217_n409, DP_mult_217_n408, DP_mult_217_n407,
         DP_mult_217_n406, DP_mult_217_n405, DP_mult_217_n404,
         DP_mult_217_n403, DP_mult_217_n402, DP_mult_217_n401,
         DP_mult_217_n400, DP_mult_217_n399, DP_mult_217_n398,
         DP_mult_217_n397, DP_mult_217_n396, DP_mult_217_n395,
         DP_mult_217_n394, DP_mult_217_n393, DP_mult_217_n392,
         DP_mult_217_n391, DP_mult_217_n390, DP_mult_217_n389,
         DP_mult_217_n387, DP_mult_217_n386, DP_mult_217_n385,
         DP_mult_217_n384, DP_mult_217_n383, DP_mult_217_n382,
         DP_mult_217_n381, DP_mult_217_n380, DP_mult_217_n379,
         DP_mult_217_n378, DP_mult_217_n377, DP_mult_217_n376,
         DP_mult_217_n375, DP_mult_217_n374, DP_mult_217_n373,
         DP_mult_217_n372, DP_mult_217_n371, DP_mult_217_n370,
         DP_mult_217_n368, DP_mult_217_n367, DP_mult_217_n366,
         DP_mult_217_n365, DP_mult_217_n364, DP_mult_217_n363,
         DP_mult_217_n362, DP_mult_217_n361, DP_mult_217_n360,
         DP_mult_217_n359, DP_mult_217_n358, DP_mult_217_n356,
         DP_mult_217_n355, DP_mult_217_n354, DP_mult_217_n353,
         DP_mult_217_n352, DP_mult_217_n351, DP_mult_217_n326,
         DP_mult_217_n325, DP_mult_217_n324, DP_mult_217_n323,
         DP_mult_217_n322, DP_mult_217_n321, DP_mult_217_n320,
         DP_mult_217_n319, DP_mult_217_n318, DP_mult_217_n317,
         DP_mult_217_n316, DP_mult_217_n315, DP_mult_217_n314,
         DP_mult_217_n313, DP_mult_217_n312, DP_mult_217_n311,
         DP_mult_217_n310, DP_mult_217_n309, DP_mult_217_n308,
         DP_mult_217_n307, DP_mult_217_n306, DP_mult_217_n305,
         DP_mult_217_n304, DP_mult_217_n303, DP_mult_215_n2162,
         DP_mult_215_n2161, DP_mult_215_n2160, DP_mult_215_n2159,
         DP_mult_215_n2158, DP_mult_215_n2157, DP_mult_215_n2156,
         DP_mult_215_n2155, DP_mult_215_n2154, DP_mult_215_n2153,
         DP_mult_215_n2152, DP_mult_215_n2151, DP_mult_215_n2150,
         DP_mult_215_n2149, DP_mult_215_n2148, DP_mult_215_n2147,
         DP_mult_215_n2146, DP_mult_215_n2145, DP_mult_215_n2144,
         DP_mult_215_n2143, DP_mult_215_n2142, DP_mult_215_n2141,
         DP_mult_215_n2140, DP_mult_215_n2139, DP_mult_215_n2138,
         DP_mult_215_n2137, DP_mult_215_n2136, DP_mult_215_n2135,
         DP_mult_215_n2134, DP_mult_215_n2133, DP_mult_215_n2132,
         DP_mult_215_n2131, DP_mult_215_n2130, DP_mult_215_n2129,
         DP_mult_215_n2128, DP_mult_215_n2127, DP_mult_215_n2126,
         DP_mult_215_n2125, DP_mult_215_n2124, DP_mult_215_n2123,
         DP_mult_215_n2122, DP_mult_215_n2121, DP_mult_215_n2120,
         DP_mult_215_n2119, DP_mult_215_n2118, DP_mult_215_n2117,
         DP_mult_215_n2116, DP_mult_215_n2115, DP_mult_215_n2114,
         DP_mult_215_n2113, DP_mult_215_n2112, DP_mult_215_n2111,
         DP_mult_215_n2110, DP_mult_215_n2109, DP_mult_215_n2108,
         DP_mult_215_n2107, DP_mult_215_n2106, DP_mult_215_n2105,
         DP_mult_215_n2104, DP_mult_215_n2103, DP_mult_215_n2102,
         DP_mult_215_n2101, DP_mult_215_n2100, DP_mult_215_n2099,
         DP_mult_215_n2098, DP_mult_215_n2097, DP_mult_215_n2096,
         DP_mult_215_n2095, DP_mult_215_n2094, DP_mult_215_n2093,
         DP_mult_215_n2092, DP_mult_215_n2091, DP_mult_215_n2090,
         DP_mult_215_n2089, DP_mult_215_n2088, DP_mult_215_n2087,
         DP_mult_215_n2086, DP_mult_215_n2085, DP_mult_215_n2084,
         DP_mult_215_n2083, DP_mult_215_n2082, DP_mult_215_n2081,
         DP_mult_215_n2080, DP_mult_215_n2079, DP_mult_215_n2078,
         DP_mult_215_n2077, DP_mult_215_n2076, DP_mult_215_n2075,
         DP_mult_215_n2074, DP_mult_215_n2073, DP_mult_215_n2072,
         DP_mult_215_n2071, DP_mult_215_n2070, DP_mult_215_n2069,
         DP_mult_215_n2068, DP_mult_215_n2067, DP_mult_215_n2066,
         DP_mult_215_n2065, DP_mult_215_n2064, DP_mult_215_n2063,
         DP_mult_215_n2062, DP_mult_215_n2061, DP_mult_215_n2060,
         DP_mult_215_n2059, DP_mult_215_n2058, DP_mult_215_n2057,
         DP_mult_215_n2056, DP_mult_215_n2055, DP_mult_215_n2054,
         DP_mult_215_n2053, DP_mult_215_n2052, DP_mult_215_n2051,
         DP_mult_215_n2050, DP_mult_215_n2049, DP_mult_215_n2048,
         DP_mult_215_n2047, DP_mult_215_n2046, DP_mult_215_n2045,
         DP_mult_215_n2044, DP_mult_215_n2043, DP_mult_215_n2042,
         DP_mult_215_n2041, DP_mult_215_n2040, DP_mult_215_n2039,
         DP_mult_215_n2038, DP_mult_215_n2037, DP_mult_215_n2036,
         DP_mult_215_n2035, DP_mult_215_n2034, DP_mult_215_n2033,
         DP_mult_215_n2032, DP_mult_215_n2031, DP_mult_215_n2030,
         DP_mult_215_n2029, DP_mult_215_n2028, DP_mult_215_n2027,
         DP_mult_215_n2026, DP_mult_215_n2025, DP_mult_215_n2024,
         DP_mult_215_n2023, DP_mult_215_n2022, DP_mult_215_n2021,
         DP_mult_215_n2020, DP_mult_215_n2019, DP_mult_215_n2018,
         DP_mult_215_n2017, DP_mult_215_n2016, DP_mult_215_n2015,
         DP_mult_215_n2014, DP_mult_215_n2013, DP_mult_215_n2012,
         DP_mult_215_n2011, DP_mult_215_n2010, DP_mult_215_n2009,
         DP_mult_215_n2008, DP_mult_215_n2007, DP_mult_215_n2006,
         DP_mult_215_n2005, DP_mult_215_n2004, DP_mult_215_n2003,
         DP_mult_215_n2002, DP_mult_215_n2001, DP_mult_215_n2000,
         DP_mult_215_n1999, DP_mult_215_n1998, DP_mult_215_n1997,
         DP_mult_215_n1996, DP_mult_215_n1995, DP_mult_215_n1994,
         DP_mult_215_n1993, DP_mult_215_n1992, DP_mult_215_n1991,
         DP_mult_215_n1990, DP_mult_215_n1989, DP_mult_215_n1988,
         DP_mult_215_n1987, DP_mult_215_n1986, DP_mult_215_n1985,
         DP_mult_215_n1984, DP_mult_215_n1983, DP_mult_215_n1982,
         DP_mult_215_n1981, DP_mult_215_n1980, DP_mult_215_n1979,
         DP_mult_215_n1978, DP_mult_215_n1977, DP_mult_215_n1976,
         DP_mult_215_n1975, DP_mult_215_n1974, DP_mult_215_n1973,
         DP_mult_215_n1972, DP_mult_215_n1971, DP_mult_215_n1970,
         DP_mult_215_n1969, DP_mult_215_n1968, DP_mult_215_n1967,
         DP_mult_215_n1966, DP_mult_215_n1965, DP_mult_215_n1964,
         DP_mult_215_n1963, DP_mult_215_n1962, DP_mult_215_n1961,
         DP_mult_215_n1960, DP_mult_215_n1959, DP_mult_215_n1958,
         DP_mult_215_n1957, DP_mult_215_n1956, DP_mult_215_n1955,
         DP_mult_215_n1954, DP_mult_215_n1953, DP_mult_215_n1952,
         DP_mult_215_n1951, DP_mult_215_n1950, DP_mult_215_n1949,
         DP_mult_215_n1948, DP_mult_215_n1947, DP_mult_215_n1946,
         DP_mult_215_n1945, DP_mult_215_n1944, DP_mult_215_n1943,
         DP_mult_215_n1942, DP_mult_215_n1941, DP_mult_215_n1940,
         DP_mult_215_n1939, DP_mult_215_n1938, DP_mult_215_n1937,
         DP_mult_215_n1936, DP_mult_215_n1935, DP_mult_215_n1934,
         DP_mult_215_n1933, DP_mult_215_n1932, DP_mult_215_n1931,
         DP_mult_215_n1930, DP_mult_215_n1929, DP_mult_215_n1928,
         DP_mult_215_n1927, DP_mult_215_n1926, DP_mult_215_n1925,
         DP_mult_215_n1924, DP_mult_215_n1923, DP_mult_215_n1922,
         DP_mult_215_n1921, DP_mult_215_n1920, DP_mult_215_n1919,
         DP_mult_215_n1918, DP_mult_215_n1917, DP_mult_215_n1916,
         DP_mult_215_n1915, DP_mult_215_n1914, DP_mult_215_n1913,
         DP_mult_215_n1912, DP_mult_215_n1911, DP_mult_215_n1910,
         DP_mult_215_n1909, DP_mult_215_n1908, DP_mult_215_n1907,
         DP_mult_215_n1906, DP_mult_215_n1905, DP_mult_215_n1904,
         DP_mult_215_n1903, DP_mult_215_n1902, DP_mult_215_n1901,
         DP_mult_215_n1900, DP_mult_215_n1899, DP_mult_215_n1898,
         DP_mult_215_n1897, DP_mult_215_n1896, DP_mult_215_n1895,
         DP_mult_215_n1894, DP_mult_215_n1893, DP_mult_215_n1892,
         DP_mult_215_n1891, DP_mult_215_n1890, DP_mult_215_n1889,
         DP_mult_215_n1888, DP_mult_215_n1887, DP_mult_215_n1886,
         DP_mult_215_n1885, DP_mult_215_n1884, DP_mult_215_n1883,
         DP_mult_215_n1882, DP_mult_215_n1881, DP_mult_215_n1880,
         DP_mult_215_n1879, DP_mult_215_n1878, DP_mult_215_n1877,
         DP_mult_215_n1876, DP_mult_215_n1875, DP_mult_215_n1874,
         DP_mult_215_n1873, DP_mult_215_n1872, DP_mult_215_n1871,
         DP_mult_215_n1870, DP_mult_215_n1869, DP_mult_215_n1868,
         DP_mult_215_n1867, DP_mult_215_n1866, DP_mult_215_n1865,
         DP_mult_215_n1864, DP_mult_215_n1863, DP_mult_215_n1862,
         DP_mult_215_n1861, DP_mult_215_n1860, DP_mult_215_n1859,
         DP_mult_215_n1858, DP_mult_215_n1857, DP_mult_215_n1856,
         DP_mult_215_n1855, DP_mult_215_n1854, DP_mult_215_n1853,
         DP_mult_215_n1852, DP_mult_215_n1851, DP_mult_215_n1850,
         DP_mult_215_n1849, DP_mult_215_n1848, DP_mult_215_n1847,
         DP_mult_215_n1846, DP_mult_215_n1845, DP_mult_215_n1844,
         DP_mult_215_n1843, DP_mult_215_n1842, DP_mult_215_n1841,
         DP_mult_215_n1840, DP_mult_215_n1839, DP_mult_215_n1838,
         DP_mult_215_n1837, DP_mult_215_n1836, DP_mult_215_n1835,
         DP_mult_215_n1834, DP_mult_215_n1833, DP_mult_215_n1832,
         DP_mult_215_n1831, DP_mult_215_n1830, DP_mult_215_n1829,
         DP_mult_215_n1828, DP_mult_215_n1827, DP_mult_215_n1826,
         DP_mult_215_n1825, DP_mult_215_n1824, DP_mult_215_n1823,
         DP_mult_215_n1822, DP_mult_215_n1821, DP_mult_215_n1820,
         DP_mult_215_n1819, DP_mult_215_n1818, DP_mult_215_n1817,
         DP_mult_215_n1816, DP_mult_215_n1815, DP_mult_215_n1814,
         DP_mult_215_n1813, DP_mult_215_n1812, DP_mult_215_n1811,
         DP_mult_215_n1810, DP_mult_215_n1809, DP_mult_215_n1808,
         DP_mult_215_n1807, DP_mult_215_n1806, DP_mult_215_n1805,
         DP_mult_215_n1804, DP_mult_215_n1803, DP_mult_215_n1802,
         DP_mult_215_n1801, DP_mult_215_n1800, DP_mult_215_n1799,
         DP_mult_215_n1798, DP_mult_215_n1797, DP_mult_215_n1796,
         DP_mult_215_n1795, DP_mult_215_n1794, DP_mult_215_n1793,
         DP_mult_215_n1792, DP_mult_215_n1791, DP_mult_215_n1790,
         DP_mult_215_n1789, DP_mult_215_n1788, DP_mult_215_n1787,
         DP_mult_215_n1786, DP_mult_215_n1785, DP_mult_215_n1784,
         DP_mult_215_n1783, DP_mult_215_n1782, DP_mult_215_n1781,
         DP_mult_215_n1780, DP_mult_215_n1779, DP_mult_215_n1778,
         DP_mult_215_n1777, DP_mult_215_n1776, DP_mult_215_n1775,
         DP_mult_215_n1774, DP_mult_215_n1773, DP_mult_215_n1772,
         DP_mult_215_n1771, DP_mult_215_n1770, DP_mult_215_n1769,
         DP_mult_215_n1768, DP_mult_215_n1767, DP_mult_215_n1766,
         DP_mult_215_n1765, DP_mult_215_n1764, DP_mult_215_n1763,
         DP_mult_215_n1762, DP_mult_215_n1761, DP_mult_215_n1760,
         DP_mult_215_n1759, DP_mult_215_n1758, DP_mult_215_n1757,
         DP_mult_215_n1756, DP_mult_215_n1755, DP_mult_215_n1754,
         DP_mult_215_n1753, DP_mult_215_n1752, DP_mult_215_n1751,
         DP_mult_215_n1750, DP_mult_215_n1749, DP_mult_215_n1748,
         DP_mult_215_n1747, DP_mult_215_n1746, DP_mult_215_n1745,
         DP_mult_215_n1744, DP_mult_215_n1743, DP_mult_215_n1742,
         DP_mult_215_n1741, DP_mult_215_n1740, DP_mult_215_n1739,
         DP_mult_215_n1738, DP_mult_215_n1737, DP_mult_215_n1736,
         DP_mult_215_n1735, DP_mult_215_n1734, DP_mult_215_n1733,
         DP_mult_215_n1732, DP_mult_215_n1731, DP_mult_215_n1730,
         DP_mult_215_n1729, DP_mult_215_n1728, DP_mult_215_n1727,
         DP_mult_215_n1726, DP_mult_215_n1725, DP_mult_215_n1724,
         DP_mult_215_n1723, DP_mult_215_n1722, DP_mult_215_n1721,
         DP_mult_215_n1720, DP_mult_215_n1719, DP_mult_215_n1718,
         DP_mult_215_n1717, DP_mult_215_n1716, DP_mult_215_n1715,
         DP_mult_215_n1714, DP_mult_215_n1713, DP_mult_215_n1712,
         DP_mult_215_n1711, DP_mult_215_n1710, DP_mult_215_n1709,
         DP_mult_215_n1708, DP_mult_215_n1707, DP_mult_215_n1706,
         DP_mult_215_n1705, DP_mult_215_n1704, DP_mult_215_n1703,
         DP_mult_215_n1702, DP_mult_215_n1701, DP_mult_215_n1700,
         DP_mult_215_n1699, DP_mult_215_n1698, DP_mult_215_n1697,
         DP_mult_215_n1696, DP_mult_215_n1695, DP_mult_215_n1694,
         DP_mult_215_n1693, DP_mult_215_n1692, DP_mult_215_n1691,
         DP_mult_215_n1690, DP_mult_215_n1689, DP_mult_215_n1688,
         DP_mult_215_n1687, DP_mult_215_n1686, DP_mult_215_n1685,
         DP_mult_215_n1684, DP_mult_215_n1683, DP_mult_215_n1682,
         DP_mult_215_n1681, DP_mult_215_n1680, DP_mult_215_n1679,
         DP_mult_215_n1678, DP_mult_215_n1677, DP_mult_215_n1676,
         DP_mult_215_n1675, DP_mult_215_n1674, DP_mult_215_n1673,
         DP_mult_215_n1672, DP_mult_215_n1671, DP_mult_215_n1670,
         DP_mult_215_n1669, DP_mult_215_n1668, DP_mult_215_n1667,
         DP_mult_215_n1666, DP_mult_215_n1665, DP_mult_215_n1664,
         DP_mult_215_n1663, DP_mult_215_n1662, DP_mult_215_n1661,
         DP_mult_215_n1660, DP_mult_215_n1659, DP_mult_215_n1658,
         DP_mult_215_n1657, DP_mult_215_n1656, DP_mult_215_n1655,
         DP_mult_215_n1654, DP_mult_215_n1653, DP_mult_215_n1652,
         DP_mult_215_n1651, DP_mult_215_n1650, DP_mult_215_n1649,
         DP_mult_215_n1648, DP_mult_215_n1647, DP_mult_215_n1646,
         DP_mult_215_n1645, DP_mult_215_n1644, DP_mult_215_n1643,
         DP_mult_215_n1642, DP_mult_215_n1641, DP_mult_215_n1640,
         DP_mult_215_n1639, DP_mult_215_n1638, DP_mult_215_n1637,
         DP_mult_215_n1636, DP_mult_215_n1635, DP_mult_215_n1634,
         DP_mult_215_n1633, DP_mult_215_n1632, DP_mult_215_n1631,
         DP_mult_215_n1630, DP_mult_215_n1629, DP_mult_215_n1628,
         DP_mult_215_n1627, DP_mult_215_n1626, DP_mult_215_n1625,
         DP_mult_215_n1624, DP_mult_215_n1623, DP_mult_215_n1622,
         DP_mult_215_n1621, DP_mult_215_n1620, DP_mult_215_n1619,
         DP_mult_215_n1618, DP_mult_215_n1617, DP_mult_215_n1616,
         DP_mult_215_n1615, DP_mult_215_n1614, DP_mult_215_n1613,
         DP_mult_215_n1612, DP_mult_215_n1611, DP_mult_215_n1610,
         DP_mult_215_n1609, DP_mult_215_n1608, DP_mult_215_n1607,
         DP_mult_215_n1606, DP_mult_215_n1605, DP_mult_215_n1604,
         DP_mult_215_n1603, DP_mult_215_n1602, DP_mult_215_n1601,
         DP_mult_215_n1600, DP_mult_215_n1599, DP_mult_215_n1598,
         DP_mult_215_n1597, DP_mult_215_n1596, DP_mult_215_n1595,
         DP_mult_215_n1594, DP_mult_215_n1593, DP_mult_215_n1592,
         DP_mult_215_n1591, DP_mult_215_n1590, DP_mult_215_n1589,
         DP_mult_215_n1588, DP_mult_215_n1587, DP_mult_215_n1586,
         DP_mult_215_n1585, DP_mult_215_n1584, DP_mult_215_n1583,
         DP_mult_215_n1582, DP_mult_215_n1581, DP_mult_215_n1580,
         DP_mult_215_n1579, DP_mult_215_n1578, DP_mult_215_n1577,
         DP_mult_215_n1576, DP_mult_215_n1575, DP_mult_215_n1574,
         DP_mult_215_n1573, DP_mult_215_n1572, DP_mult_215_n1571,
         DP_mult_215_n1570, DP_mult_215_n1569, DP_mult_215_n1568,
         DP_mult_215_n1567, DP_mult_215_n1566, DP_mult_215_n1565,
         DP_mult_215_n1564, DP_mult_215_n1563, DP_mult_215_n1562,
         DP_mult_215_n1561, DP_mult_215_n1560, DP_mult_215_n1559,
         DP_mult_215_n1558, DP_mult_215_n1557, DP_mult_215_n1556,
         DP_mult_215_n1555, DP_mult_215_n1554, DP_mult_215_n1553,
         DP_mult_215_n1552, DP_mult_215_n1551, DP_mult_215_n1550,
         DP_mult_215_n1549, DP_mult_215_n1548, DP_mult_215_n1547,
         DP_mult_215_n1546, DP_mult_215_n1545, DP_mult_215_n1544,
         DP_mult_215_n1543, DP_mult_215_n1542, DP_mult_215_n1541,
         DP_mult_215_n1540, DP_mult_215_n1539, DP_mult_215_n1538,
         DP_mult_215_n1537, DP_mult_215_n1536, DP_mult_215_n1535,
         DP_mult_215_n1534, DP_mult_215_n1533, DP_mult_215_n1397,
         DP_mult_215_n1396, DP_mult_215_n1395, DP_mult_215_n1394,
         DP_mult_215_n1393, DP_mult_215_n1392, DP_mult_215_n1391,
         DP_mult_215_n1390, DP_mult_215_n1389, DP_mult_215_n1388,
         DP_mult_215_n1387, DP_mult_215_n1386, DP_mult_215_n1385,
         DP_mult_215_n1384, DP_mult_215_n1383, DP_mult_215_n1382,
         DP_mult_215_n1381, DP_mult_215_n1380, DP_mult_215_n1379,
         DP_mult_215_n1378, DP_mult_215_n1377, DP_mult_215_n1376,
         DP_mult_215_n1375, DP_mult_215_n1374, DP_mult_215_n908,
         DP_mult_215_n907, DP_mult_215_n906, DP_mult_215_n904,
         DP_mult_215_n903, DP_mult_215_n902, DP_mult_215_n901,
         DP_mult_215_n900, DP_mult_215_n899, DP_mult_215_n898,
         DP_mult_215_n897, DP_mult_215_n896, DP_mult_215_n895,
         DP_mult_215_n894, DP_mult_215_n893, DP_mult_215_n892,
         DP_mult_215_n891, DP_mult_215_n890, DP_mult_215_n889,
         DP_mult_215_n888, DP_mult_215_n887, DP_mult_215_n886,
         DP_mult_215_n885, DP_mult_215_n884, DP_mult_215_n883,
         DP_mult_215_n882, DP_mult_215_n881, DP_mult_215_n880,
         DP_mult_215_n879, DP_mult_215_n878, DP_mult_215_n877,
         DP_mult_215_n876, DP_mult_215_n875, DP_mult_215_n874,
         DP_mult_215_n873, DP_mult_215_n872, DP_mult_215_n871,
         DP_mult_215_n870, DP_mult_215_n869, DP_mult_215_n868,
         DP_mult_215_n867, DP_mult_215_n866, DP_mult_215_n865,
         DP_mult_215_n864, DP_mult_215_n863, DP_mult_215_n862,
         DP_mult_215_n861, DP_mult_215_n860, DP_mult_215_n859,
         DP_mult_215_n858, DP_mult_215_n857, DP_mult_215_n856,
         DP_mult_215_n855, DP_mult_215_n854, DP_mult_215_n853,
         DP_mult_215_n852, DP_mult_215_n851, DP_mult_215_n850,
         DP_mult_215_n849, DP_mult_215_n848, DP_mult_215_n847,
         DP_mult_215_n846, DP_mult_215_n845, DP_mult_215_n844,
         DP_mult_215_n843, DP_mult_215_n842, DP_mult_215_n841,
         DP_mult_215_n840, DP_mult_215_n839, DP_mult_215_n838,
         DP_mult_215_n837, DP_mult_215_n836, DP_mult_215_n835,
         DP_mult_215_n834, DP_mult_215_n833, DP_mult_215_n832,
         DP_mult_215_n831, DP_mult_215_n830, DP_mult_215_n829,
         DP_mult_215_n828, DP_mult_215_n827, DP_mult_215_n826,
         DP_mult_215_n825, DP_mult_215_n824, DP_mult_215_n823,
         DP_mult_215_n822, DP_mult_215_n821, DP_mult_215_n820,
         DP_mult_215_n819, DP_mult_215_n818, DP_mult_215_n817,
         DP_mult_215_n816, DP_mult_215_n815, DP_mult_215_n814,
         DP_mult_215_n813, DP_mult_215_n812, DP_mult_215_n811,
         DP_mult_215_n810, DP_mult_215_n809, DP_mult_215_n808,
         DP_mult_215_n807, DP_mult_215_n806, DP_mult_215_n805,
         DP_mult_215_n804, DP_mult_215_n803, DP_mult_215_n802,
         DP_mult_215_n801, DP_mult_215_n800, DP_mult_215_n799,
         DP_mult_215_n798, DP_mult_215_n797, DP_mult_215_n796,
         DP_mult_215_n795, DP_mult_215_n794, DP_mult_215_n793,
         DP_mult_215_n792, DP_mult_215_n791, DP_mult_215_n790,
         DP_mult_215_n789, DP_mult_215_n788, DP_mult_215_n787,
         DP_mult_215_n786, DP_mult_215_n785, DP_mult_215_n784,
         DP_mult_215_n783, DP_mult_215_n782, DP_mult_215_n781,
         DP_mult_215_n780, DP_mult_215_n779, DP_mult_215_n778,
         DP_mult_215_n777, DP_mult_215_n776, DP_mult_215_n775,
         DP_mult_215_n774, DP_mult_215_n773, DP_mult_215_n772,
         DP_mult_215_n771, DP_mult_215_n770, DP_mult_215_n769,
         DP_mult_215_n768, DP_mult_215_n767, DP_mult_215_n766,
         DP_mult_215_n765, DP_mult_215_n764, DP_mult_215_n763,
         DP_mult_215_n762, DP_mult_215_n761, DP_mult_215_n760,
         DP_mult_215_n759, DP_mult_215_n758, DP_mult_215_n757,
         DP_mult_215_n756, DP_mult_215_n755, DP_mult_215_n754,
         DP_mult_215_n753, DP_mult_215_n752, DP_mult_215_n751,
         DP_mult_215_n750, DP_mult_215_n749, DP_mult_215_n748,
         DP_mult_215_n747, DP_mult_215_n746, DP_mult_215_n745,
         DP_mult_215_n744, DP_mult_215_n743, DP_mult_215_n742,
         DP_mult_215_n741, DP_mult_215_n740, DP_mult_215_n739,
         DP_mult_215_n738, DP_mult_215_n737, DP_mult_215_n736,
         DP_mult_215_n735, DP_mult_215_n734, DP_mult_215_n733,
         DP_mult_215_n732, DP_mult_215_n731, DP_mult_215_n730,
         DP_mult_215_n729, DP_mult_215_n727, DP_mult_215_n726,
         DP_mult_215_n725, DP_mult_215_n724, DP_mult_215_n723,
         DP_mult_215_n722, DP_mult_215_n721, DP_mult_215_n720,
         DP_mult_215_n719, DP_mult_215_n718, DP_mult_215_n717,
         DP_mult_215_n716, DP_mult_215_n715, DP_mult_215_n714,
         DP_mult_215_n713, DP_mult_215_n712, DP_mult_215_n711,
         DP_mult_215_n710, DP_mult_215_n709, DP_mult_215_n708,
         DP_mult_215_n707, DP_mult_215_n706, DP_mult_215_n688,
         DP_mult_215_n687, DP_mult_215_n686, DP_mult_215_n685,
         DP_mult_215_n684, DP_mult_215_n683, DP_mult_215_n682,
         DP_mult_215_n681, DP_mult_215_n680, DP_mult_215_n679,
         DP_mult_215_n678, DP_mult_215_n677, DP_mult_215_n676,
         DP_mult_215_n675, DP_mult_215_n674, DP_mult_215_n673,
         DP_mult_215_n672, DP_mult_215_n671, DP_mult_215_n670,
         DP_mult_215_n669, DP_mult_215_n668, DP_mult_215_n667,
         DP_mult_215_n666, DP_mult_215_n665, DP_mult_215_n664,
         DP_mult_215_n663, DP_mult_215_n662, DP_mult_215_n661,
         DP_mult_215_n660, DP_mult_215_n659, DP_mult_215_n658,
         DP_mult_215_n657, DP_mult_215_n656, DP_mult_215_n655,
         DP_mult_215_n654, DP_mult_215_n653, DP_mult_215_n652,
         DP_mult_215_n651, DP_mult_215_n650, DP_mult_215_n649,
         DP_mult_215_n648, DP_mult_215_n647, DP_mult_215_n646,
         DP_mult_215_n645, DP_mult_215_n644, DP_mult_215_n643,
         DP_mult_215_n642, DP_mult_215_n641, DP_mult_215_n640,
         DP_mult_215_n639, DP_mult_215_n638, DP_mult_215_n637,
         DP_mult_215_n636, DP_mult_215_n635, DP_mult_215_n634,
         DP_mult_215_n633, DP_mult_215_n632, DP_mult_215_n631,
         DP_mult_215_n630, DP_mult_215_n629, DP_mult_215_n628,
         DP_mult_215_n627, DP_mult_215_n626, DP_mult_215_n625,
         DP_mult_215_n624, DP_mult_215_n623, DP_mult_215_n622,
         DP_mult_215_n621, DP_mult_215_n620, DP_mult_215_n619,
         DP_mult_215_n618, DP_mult_215_n617, DP_mult_215_n616,
         DP_mult_215_n615, DP_mult_215_n614, DP_mult_215_n613,
         DP_mult_215_n612, DP_mult_215_n611, DP_mult_215_n610,
         DP_mult_215_n609, DP_mult_215_n608, DP_mult_215_n607,
         DP_mult_215_n606, DP_mult_215_n605, DP_mult_215_n604,
         DP_mult_215_n603, DP_mult_215_n602, DP_mult_215_n601,
         DP_mult_215_n600, DP_mult_215_n599, DP_mult_215_n598,
         DP_mult_215_n597, DP_mult_215_n596, DP_mult_215_n595,
         DP_mult_215_n594, DP_mult_215_n593, DP_mult_215_n592,
         DP_mult_215_n591, DP_mult_215_n590, DP_mult_215_n589,
         DP_mult_215_n588, DP_mult_215_n587, DP_mult_215_n586,
         DP_mult_215_n585, DP_mult_215_n584, DP_mult_215_n583,
         DP_mult_215_n582, DP_mult_215_n581, DP_mult_215_n580,
         DP_mult_215_n579, DP_mult_215_n578, DP_mult_215_n577,
         DP_mult_215_n576, DP_mult_215_n575, DP_mult_215_n574,
         DP_mult_215_n573, DP_mult_215_n572, DP_mult_215_n571,
         DP_mult_215_n570, DP_mult_215_n569, DP_mult_215_n568,
         DP_mult_215_n567, DP_mult_215_n566, DP_mult_215_n565,
         DP_mult_215_n564, DP_mult_215_n563, DP_mult_215_n562,
         DP_mult_215_n561, DP_mult_215_n560, DP_mult_215_n559,
         DP_mult_215_n558, DP_mult_215_n557, DP_mult_215_n556,
         DP_mult_215_n555, DP_mult_215_n554, DP_mult_215_n553,
         DP_mult_215_n552, DP_mult_215_n551, DP_mult_215_n550,
         DP_mult_215_n549, DP_mult_215_n548, DP_mult_215_n547,
         DP_mult_215_n546, DP_mult_215_n545, DP_mult_215_n544,
         DP_mult_215_n543, DP_mult_215_n542, DP_mult_215_n541,
         DP_mult_215_n540, DP_mult_215_n539, DP_mult_215_n538,
         DP_mult_215_n537, DP_mult_215_n536, DP_mult_215_n535,
         DP_mult_215_n534, DP_mult_215_n533, DP_mult_215_n532,
         DP_mult_215_n531, DP_mult_215_n530, DP_mult_215_n529,
         DP_mult_215_n528, DP_mult_215_n527, DP_mult_215_n526,
         DP_mult_215_n525, DP_mult_215_n524, DP_mult_215_n523,
         DP_mult_215_n522, DP_mult_215_n521, DP_mult_215_n520,
         DP_mult_215_n519, DP_mult_215_n518, DP_mult_215_n517,
         DP_mult_215_n516, DP_mult_215_n515, DP_mult_215_n514,
         DP_mult_215_n513, DP_mult_215_n512, DP_mult_215_n511,
         DP_mult_215_n510, DP_mult_215_n509, DP_mult_215_n508,
         DP_mult_215_n507, DP_mult_215_n506, DP_mult_215_n505,
         DP_mult_215_n504, DP_mult_215_n503, DP_mult_215_n502,
         DP_mult_215_n501, DP_mult_215_n500, DP_mult_215_n499,
         DP_mult_215_n498, DP_mult_215_n497, DP_mult_215_n496,
         DP_mult_215_n495, DP_mult_215_n494, DP_mult_215_n493,
         DP_mult_215_n492, DP_mult_215_n491, DP_mult_215_n490,
         DP_mult_215_n489, DP_mult_215_n488, DP_mult_215_n487,
         DP_mult_215_n486, DP_mult_215_n485, DP_mult_215_n484,
         DP_mult_215_n483, DP_mult_215_n482, DP_mult_215_n481,
         DP_mult_215_n479, DP_mult_215_n478, DP_mult_215_n477,
         DP_mult_215_n476, DP_mult_215_n475, DP_mult_215_n474,
         DP_mult_215_n473, DP_mult_215_n472, DP_mult_215_n471,
         DP_mult_215_n470, DP_mult_215_n469, DP_mult_215_n468,
         DP_mult_215_n467, DP_mult_215_n466, DP_mult_215_n465,
         DP_mult_215_n464, DP_mult_215_n463, DP_mult_215_n462,
         DP_mult_215_n461, DP_mult_215_n460, DP_mult_215_n459,
         DP_mult_215_n458, DP_mult_215_n457, DP_mult_215_n456,
         DP_mult_215_n455, DP_mult_215_n454, DP_mult_215_n453,
         DP_mult_215_n452, DP_mult_215_n451, DP_mult_215_n450,
         DP_mult_215_n449, DP_mult_215_n448, DP_mult_215_n447,
         DP_mult_215_n446, DP_mult_215_n445, DP_mult_215_n444,
         DP_mult_215_n442, DP_mult_215_n441, DP_mult_215_n440,
         DP_mult_215_n439, DP_mult_215_n438, DP_mult_215_n437,
         DP_mult_215_n436, DP_mult_215_n435, DP_mult_215_n434,
         DP_mult_215_n433, DP_mult_215_n432, DP_mult_215_n431,
         DP_mult_215_n430, DP_mult_215_n429, DP_mult_215_n428,
         DP_mult_215_n427, DP_mult_215_n426, DP_mult_215_n425,
         DP_mult_215_n424, DP_mult_215_n423, DP_mult_215_n422,
         DP_mult_215_n421, DP_mult_215_n420, DP_mult_215_n419,
         DP_mult_215_n418, DP_mult_215_n417, DP_mult_215_n416,
         DP_mult_215_n415, DP_mult_215_n414, DP_mult_215_n413,
         DP_mult_215_n411, DP_mult_215_n410, DP_mult_215_n409,
         DP_mult_215_n408, DP_mult_215_n407, DP_mult_215_n406,
         DP_mult_215_n405, DP_mult_215_n404, DP_mult_215_n403,
         DP_mult_215_n402, DP_mult_215_n401, DP_mult_215_n400,
         DP_mult_215_n399, DP_mult_215_n398, DP_mult_215_n397,
         DP_mult_215_n396, DP_mult_215_n395, DP_mult_215_n394,
         DP_mult_215_n393, DP_mult_215_n392, DP_mult_215_n391,
         DP_mult_215_n390, DP_mult_215_n389, DP_mult_215_n387,
         DP_mult_215_n386, DP_mult_215_n385, DP_mult_215_n384,
         DP_mult_215_n383, DP_mult_215_n382, DP_mult_215_n381,
         DP_mult_215_n380, DP_mult_215_n379, DP_mult_215_n378,
         DP_mult_215_n377, DP_mult_215_n376, DP_mult_215_n375,
         DP_mult_215_n374, DP_mult_215_n373, DP_mult_215_n372,
         DP_mult_215_n371, DP_mult_215_n370, DP_mult_215_n368,
         DP_mult_215_n367, DP_mult_215_n366, DP_mult_215_n365,
         DP_mult_215_n364, DP_mult_215_n363, DP_mult_215_n362,
         DP_mult_215_n361, DP_mult_215_n360, DP_mult_215_n359,
         DP_mult_215_n358, DP_mult_215_n356, DP_mult_215_n355,
         DP_mult_215_n354, DP_mult_215_n353, DP_mult_215_n352,
         DP_mult_215_n351, DP_mult_215_n326, DP_mult_215_n325,
         DP_mult_215_n324, DP_mult_215_n323, DP_mult_215_n322,
         DP_mult_215_n321, DP_mult_215_n320, DP_mult_215_n319,
         DP_mult_215_n318, DP_mult_215_n317, DP_mult_215_n316,
         DP_mult_215_n315, DP_mult_215_n314, DP_mult_215_n313,
         DP_mult_215_n312, DP_mult_215_n311, DP_mult_215_n310,
         DP_mult_215_n309, DP_mult_215_n308, DP_mult_215_n307,
         DP_mult_215_n306, DP_mult_215_n305, DP_mult_215_n304,
         DP_mult_215_n303, DP_mult_216_n1266, DP_mult_216_n1265,
         DP_mult_216_n1264, DP_mult_216_n1263, DP_mult_216_n1262,
         DP_mult_216_n1261, DP_mult_216_n1260, DP_mult_216_n1259,
         DP_mult_216_n1258, DP_mult_216_n1257, DP_mult_216_n1256,
         DP_mult_216_n1255, DP_mult_216_n1254, DP_mult_216_n1253,
         DP_mult_216_n1252, DP_mult_216_n1251, DP_mult_216_n1250,
         DP_mult_216_n1249, DP_mult_216_n1248, DP_mult_216_n1247,
         DP_mult_216_n1246, DP_mult_216_n1245, DP_mult_216_n1244,
         DP_mult_216_n1243, DP_mult_216_n1242, DP_mult_216_n1241,
         DP_mult_216_n1240, DP_mult_216_n1239, DP_mult_216_n1238,
         DP_mult_216_n1237, DP_mult_216_n1236, DP_mult_216_n1235,
         DP_mult_216_n1234, DP_mult_216_n1233, DP_mult_216_n1232,
         DP_mult_216_n1231, DP_mult_216_n1230, DP_mult_216_n1229,
         DP_mult_216_n1228, DP_mult_216_n1227, DP_mult_216_n1226,
         DP_mult_216_n1225, DP_mult_216_n1224, DP_mult_216_n1223,
         DP_mult_216_n1222, DP_mult_216_n1221, DP_mult_216_n1220,
         DP_mult_216_n1219, DP_mult_216_n1218, DP_mult_216_n1217,
         DP_mult_216_n1216, DP_mult_216_n1215, DP_mult_216_n1214,
         DP_mult_216_n1213, DP_mult_216_n1212, DP_mult_216_n1211,
         DP_mult_216_n1210, DP_mult_216_n1209, DP_mult_216_n1208,
         DP_mult_216_n1207, DP_mult_216_n1206, DP_mult_216_n1205,
         DP_mult_216_n1204, DP_mult_216_n1203, DP_mult_216_n1202,
         DP_mult_216_n1201, DP_mult_216_n1200, DP_mult_216_n1199,
         DP_mult_216_n1198, DP_mult_216_n1197, DP_mult_216_n1196,
         DP_mult_216_n1195, DP_mult_216_n1194, DP_mult_216_n1193,
         DP_mult_216_n1192, DP_mult_216_n1191, DP_mult_216_n1190,
         DP_mult_216_n1189, DP_mult_216_n1188, DP_mult_216_n1187,
         DP_mult_216_n1186, DP_mult_216_n1185, DP_mult_216_n1184,
         DP_mult_216_n1183, DP_mult_216_n1182, DP_mult_216_n1181,
         DP_mult_216_n1180, DP_mult_216_n1179, DP_mult_216_n1178,
         DP_mult_216_n1177, DP_mult_216_n1176, DP_mult_216_n1175,
         DP_mult_216_n1174, DP_mult_216_n1173, DP_mult_216_n1172,
         DP_mult_216_n1171, DP_mult_216_n1170, DP_mult_216_n1169,
         DP_mult_216_n1168, DP_mult_216_n1167, DP_mult_216_n1166,
         DP_mult_216_n1165, DP_mult_216_n1164, DP_mult_216_n1163,
         DP_mult_216_n1162, DP_mult_216_n1161, DP_mult_216_n1160,
         DP_mult_216_n1159, DP_mult_216_n1158, DP_mult_216_n1157,
         DP_mult_216_n1156, DP_mult_216_n1155, DP_mult_216_n1154,
         DP_mult_216_n1153, DP_mult_216_n1152, DP_mult_216_n1151,
         DP_mult_216_n1150, DP_mult_216_n1149, DP_mult_216_n1148,
         DP_mult_216_n1147, DP_mult_216_n1146, DP_mult_216_n1145,
         DP_mult_216_n1144, DP_mult_216_n1143, DP_mult_216_n1142,
         DP_mult_216_n1141, DP_mult_216_n1140, DP_mult_216_n1139,
         DP_mult_216_n1138, DP_mult_216_n1137, DP_mult_216_n1136,
         DP_mult_216_n1135, DP_mult_216_n1134, DP_mult_216_n1133,
         DP_mult_216_n1132, DP_mult_216_n1131, DP_mult_216_n1130,
         DP_mult_216_n1129, DP_mult_216_n1128, DP_mult_216_n1127,
         DP_mult_216_n1126, DP_mult_216_n1125, DP_mult_216_n1124,
         DP_mult_216_n1123, DP_mult_216_n1122, DP_mult_216_n1121,
         DP_mult_216_n1120, DP_mult_216_n1119, DP_mult_216_n1118,
         DP_mult_216_n1117, DP_mult_216_n1116, DP_mult_216_n1115,
         DP_mult_216_n1114, DP_mult_216_n1113, DP_mult_216_n1112,
         DP_mult_216_n1111, DP_mult_216_n1110, DP_mult_216_n1109,
         DP_mult_216_n1108, DP_mult_216_n1107, DP_mult_216_n1106,
         DP_mult_216_n1105, DP_mult_216_n1104, DP_mult_216_n1103,
         DP_mult_216_n1102, DP_mult_216_n1101, DP_mult_216_n1100,
         DP_mult_216_n1099, DP_mult_216_n1098, DP_mult_216_n1097,
         DP_mult_216_n1096, DP_mult_216_n1095, DP_mult_216_n1094,
         DP_mult_216_n1093, DP_mult_216_n1092, DP_mult_216_n1091,
         DP_mult_216_n1090, DP_mult_216_n1089, DP_mult_216_n1088,
         DP_mult_216_n1087, DP_mult_216_n1086, DP_mult_216_n1085,
         DP_mult_216_n1084, DP_mult_216_n1083, DP_mult_216_n1082,
         DP_mult_216_n1081, DP_mult_216_n1080, DP_mult_216_n1079,
         DP_mult_216_n1078, DP_mult_216_n1077, DP_mult_216_n1076,
         DP_mult_216_n1075, DP_mult_216_n1074, DP_mult_216_n1073,
         DP_mult_216_n1072, DP_mult_216_n1071, DP_mult_216_n1070,
         DP_mult_216_n1069, DP_mult_216_n1068, DP_mult_216_n1067,
         DP_mult_216_n1066, DP_mult_216_n1065, DP_mult_216_n1064,
         DP_mult_216_n1063, DP_mult_216_n1062, DP_mult_216_n1061,
         DP_mult_216_n1060, DP_mult_216_n1059, DP_mult_216_n1058,
         DP_mult_216_n1057, DP_mult_216_n1056, DP_mult_216_n1055,
         DP_mult_216_n1054, DP_mult_216_n1053, DP_mult_216_n1052,
         DP_mult_216_n1051, DP_mult_216_n1050, DP_mult_216_n1049,
         DP_mult_216_n1048, DP_mult_216_n1047, DP_mult_216_n1046,
         DP_mult_216_n1045, DP_mult_216_n1044, DP_mult_216_n1043,
         DP_mult_216_n1042, DP_mult_216_n1041, DP_mult_216_n1040,
         DP_mult_216_n1039, DP_mult_216_n1038, DP_mult_216_n1037,
         DP_mult_216_n1036, DP_mult_216_n1035, DP_mult_216_n1034,
         DP_mult_216_n1033, DP_mult_216_n1032, DP_mult_216_n1031,
         DP_mult_216_n1030, DP_mult_216_n1029, DP_mult_216_n1028,
         DP_mult_216_n1027, DP_mult_216_n1026, DP_mult_216_n1025,
         DP_mult_216_n1024, DP_mult_216_n1023, DP_mult_216_n1022,
         DP_mult_216_n1021, DP_mult_216_n1020, DP_mult_216_n1019,
         DP_mult_216_n1018, DP_mult_216_n1017, DP_mult_216_n1016,
         DP_mult_216_n1015, DP_mult_216_n1014, DP_mult_216_n1013,
         DP_mult_216_n1012, DP_mult_216_n1011, DP_mult_216_n1010,
         DP_mult_216_n1009, DP_mult_216_n1008, DP_mult_216_n1007,
         DP_mult_216_n1006, DP_mult_216_n1005, DP_mult_216_n1004,
         DP_mult_216_n1003, DP_mult_216_n1002, DP_mult_216_n1001,
         DP_mult_216_n1000, DP_mult_216_n999, DP_mult_216_n998,
         DP_mult_216_n997, DP_mult_216_n996, DP_mult_216_n995,
         DP_mult_216_n994, DP_mult_216_n993, DP_mult_216_n992,
         DP_mult_216_n991, DP_mult_216_n990, DP_mult_216_n989,
         DP_mult_216_n988, DP_mult_216_n987, DP_mult_216_n986,
         DP_mult_216_n985, DP_mult_216_n984, DP_mult_216_n983,
         DP_mult_216_n982, DP_mult_216_n981, DP_mult_216_n980,
         DP_mult_216_n979, DP_mult_216_n978, DP_mult_216_n977,
         DP_mult_216_n976, DP_mult_216_n975, DP_mult_216_n974,
         DP_mult_216_n973, DP_mult_216_n972, DP_mult_216_n971,
         DP_mult_216_n970, DP_mult_216_n969, DP_mult_216_n968,
         DP_mult_216_n967, DP_mult_216_n966, DP_mult_216_n965,
         DP_mult_216_n964, DP_mult_216_n963, DP_mult_216_n962,
         DP_mult_216_n961, DP_mult_216_n960, DP_mult_216_n959,
         DP_mult_216_n958, DP_mult_216_n957, DP_mult_216_n825,
         DP_mult_216_n824, DP_mult_216_n823, DP_mult_216_n822,
         DP_mult_216_n821, DP_mult_216_n820, DP_mult_216_n819,
         DP_mult_216_n818, DP_mult_216_n817, DP_mult_216_n816,
         DP_mult_216_n815, DP_mult_216_n814, DP_mult_216_n813,
         DP_mult_216_n812, DP_mult_216_n811, DP_mult_216_n810,
         DP_mult_216_n809, DP_mult_216_n808, DP_mult_216_n807,
         DP_mult_216_n806, DP_mult_216_n805, DP_mult_216_n804,
         DP_mult_216_n803, DP_mult_216_n802, DP_mult_216_n518,
         DP_mult_216_n517, DP_mult_216_n516, DP_mult_216_n515,
         DP_mult_216_n514, DP_mult_216_n513, DP_mult_216_n512,
         DP_mult_216_n511, DP_mult_216_n510, DP_mult_216_n509,
         DP_mult_216_n508, DP_mult_216_n507, DP_mult_216_n506,
         DP_mult_216_n505, DP_mult_216_n504, DP_mult_216_n503,
         DP_mult_216_n502, DP_mult_216_n501, DP_mult_216_n500,
         DP_mult_216_n499, DP_mult_216_n498, DP_mult_216_n497,
         DP_mult_216_n485, DP_mult_216_n484, DP_mult_216_n483,
         DP_mult_216_n482, DP_mult_216_n481, DP_mult_216_n480,
         DP_mult_216_n479, DP_mult_216_n478, DP_mult_216_n477,
         DP_mult_216_n476, DP_mult_216_n475, DP_mult_216_n474,
         DP_mult_216_n473, DP_mult_216_n472, DP_mult_216_n471,
         DP_mult_216_n470, DP_mult_216_n469, DP_mult_216_n468,
         DP_mult_216_n467, DP_mult_216_n466, DP_mult_216_n465,
         DP_mult_216_n464, DP_mult_216_n463, DP_mult_216_n462,
         DP_mult_216_n461, DP_mult_216_n460, DP_mult_216_n459,
         DP_mult_216_n458, DP_mult_216_n457, DP_mult_216_n456,
         DP_mult_216_n455, DP_mult_216_n454, DP_mult_216_n453,
         DP_mult_216_n452, DP_mult_216_n451, DP_mult_216_n450,
         DP_mult_216_n449, DP_mult_216_n448, DP_mult_216_n447,
         DP_mult_216_n446, DP_mult_216_n445, DP_mult_216_n444,
         DP_mult_216_n443, DP_mult_216_n442, DP_mult_216_n441,
         DP_mult_216_n440, DP_mult_216_n439, DP_mult_216_n438,
         DP_mult_216_n437, DP_mult_216_n436, DP_mult_216_n435,
         DP_mult_216_n434, DP_mult_216_n433, DP_mult_216_n432,
         DP_mult_216_n431, DP_mult_216_n430, DP_mult_216_n429,
         DP_mult_216_n428, DP_mult_216_n427, DP_mult_216_n426,
         DP_mult_216_n425, DP_mult_216_n424, DP_mult_216_n423,
         DP_mult_216_n422, DP_mult_216_n421, DP_mult_216_n420,
         DP_mult_216_n419, DP_mult_216_n418, DP_mult_216_n417,
         DP_mult_216_n416, DP_mult_216_n415, DP_mult_216_n414,
         DP_mult_216_n413, DP_mult_216_n412, DP_mult_216_n411,
         DP_mult_216_n410, DP_mult_216_n409, DP_mult_216_n408,
         DP_mult_216_n407, DP_mult_216_n406, DP_mult_216_n405,
         DP_mult_216_n404, DP_mult_216_n403, DP_mult_216_n402,
         DP_mult_216_n401, DP_mult_216_n400, DP_mult_216_n399,
         DP_mult_216_n398, DP_mult_216_n397, DP_mult_216_n396,
         DP_mult_216_n394, DP_mult_216_n393, DP_mult_216_n392,
         DP_mult_216_n391, DP_mult_216_n390, DP_mult_216_n389,
         DP_mult_216_n388, DP_mult_216_n387, DP_mult_216_n386,
         DP_mult_216_n385, DP_mult_216_n384, DP_mult_216_n383,
         DP_mult_216_n382, DP_mult_216_n381, DP_mult_216_n380,
         DP_mult_216_n379, DP_mult_216_n378, DP_mult_216_n377,
         DP_mult_216_n376, DP_mult_216_n375, DP_mult_216_n374,
         DP_mult_216_n373, DP_mult_216_n363, DP_mult_216_n362,
         DP_mult_216_n361, DP_mult_216_n360, DP_mult_216_n359,
         DP_mult_216_n358, DP_mult_216_n357, DP_mult_216_n356,
         DP_mult_216_n355, DP_mult_216_n354, DP_mult_216_n353,
         DP_mult_216_n352, DP_mult_216_n351, DP_mult_216_n350,
         DP_mult_216_n349, DP_mult_216_n348, DP_mult_216_n347,
         DP_mult_216_n346, DP_mult_216_n345, DP_mult_216_n344,
         DP_mult_216_n343, DP_mult_216_n342, DP_mult_216_n341,
         DP_mult_216_n340, DP_mult_216_n339, DP_mult_216_n338,
         DP_mult_216_n337, DP_mult_216_n336, DP_mult_216_n335,
         DP_mult_216_n334, DP_mult_216_n333, DP_mult_216_n332,
         DP_mult_216_n331, DP_mult_216_n330, DP_mult_216_n329,
         DP_mult_216_n328, DP_mult_216_n327, DP_mult_216_n326,
         DP_mult_216_n325, DP_mult_216_n324, DP_mult_216_n323,
         DP_mult_216_n322, DP_mult_216_n321, DP_mult_216_n320,
         DP_mult_216_n319, DP_mult_216_n318, DP_mult_216_n317,
         DP_mult_216_n316, DP_mult_216_n315, DP_mult_216_n314,
         DP_mult_216_n313, DP_mult_216_n312, DP_mult_216_n311,
         DP_mult_216_n310, DP_mult_216_n309, DP_mult_216_n308,
         DP_mult_216_n307, DP_mult_216_n306, DP_mult_216_n305,
         DP_mult_216_n304, DP_mult_216_n303, DP_mult_216_n302,
         DP_mult_216_n301, DP_mult_216_n300, DP_mult_216_n299,
         DP_mult_216_n298, DP_mult_216_n297, DP_mult_216_n296,
         DP_mult_216_n295, DP_mult_216_n294, DP_mult_216_n293,
         DP_mult_216_n292, DP_mult_216_n291, DP_mult_216_n290,
         DP_mult_216_n289, DP_mult_216_n288, DP_mult_216_n287,
         DP_mult_216_n286, DP_mult_216_n285, DP_mult_216_n284,
         DP_mult_216_n283, DP_mult_216_n282, DP_mult_216_n281,
         DP_mult_216_n280, DP_mult_216_n279, DP_mult_216_n278,
         DP_mult_216_n277, DP_mult_216_n276, DP_mult_216_n275,
         DP_mult_216_n274, DP_mult_216_n273, DP_mult_216_n272,
         DP_mult_216_n271, DP_mult_216_n270, DP_mult_216_n269,
         DP_mult_216_n268, DP_mult_216_n267, DP_mult_216_n266,
         DP_mult_216_n265, DP_mult_216_n264, DP_mult_216_n263,
         DP_mult_216_n262, DP_mult_216_n261, DP_mult_216_n260,
         DP_mult_216_n259, DP_mult_216_n258, DP_mult_216_n257,
         DP_mult_216_n256, DP_mult_216_n255, DP_mult_216_n254,
         DP_mult_216_n253, DP_mult_216_n252, DP_mult_216_n251,
         DP_mult_216_n250, DP_mult_216_n249, DP_mult_216_n248,
         DP_mult_216_n247, DP_mult_216_n246, DP_mult_216_n245,
         DP_mult_216_n244, DP_mult_216_n243, DP_mult_216_n242,
         DP_mult_216_n241, DP_mult_216_n240, DP_mult_216_n239,
         DP_mult_216_n238, DP_mult_216_n237, DP_mult_216_n236,
         DP_mult_216_n235, DP_mult_216_n234, DP_mult_216_n233,
         DP_mult_216_n232, DP_mult_216_n231, DP_mult_216_n230,
         DP_mult_216_n229, DP_mult_216_n228, DP_mult_216_n227,
         DP_mult_216_n226, DP_mult_216_n225, DP_mult_216_n224,
         DP_mult_216_n223, DP_mult_216_n222, DP_mult_216_n221,
         DP_mult_216_n220, DP_mult_216_n219, DP_mult_216_n218,
         DP_mult_216_n217, DP_mult_216_n216, DP_mult_216_n215,
         DP_mult_216_n214, DP_mult_216_n213, DP_mult_216_n212,
         DP_mult_216_n211, DP_mult_216_n210, DP_mult_216_n208,
         DP_mult_216_n207, DP_mult_216_n206, DP_mult_216_n205,
         DP_mult_216_n204, DP_mult_216_n203, DP_mult_216_n202,
         DP_mult_216_n201, DP_mult_216_n200, DP_mult_216_n199,
         DP_mult_216_n198, DP_mult_216_n197, DP_mult_216_n196,
         DP_mult_216_n195, DP_mult_216_n194, DP_mult_216_n193,
         DP_mult_216_n192, DP_mult_216_n191, DP_mult_216_n189,
         DP_mult_216_n188, DP_mult_216_n187, DP_mult_216_n186,
         DP_mult_216_n185, DP_mult_216_n184, DP_mult_216_n183,
         DP_mult_216_n182, DP_mult_216_n181, DP_mult_216_n180,
         DP_mult_216_n179, DP_mult_216_n177, DP_mult_216_n176,
         DP_mult_216_n175, DP_mult_216_n174, DP_mult_216_n173,
         DP_mult_216_n172, DP_mult_216_n158, DP_mult_216_n157,
         DP_mult_216_n156, DP_mult_216_n155, DP_mult_216_n154,
         DP_mult_216_n153, DP_mult_216_n152, DP_mult_216_n151,
         DP_mult_216_n150, DP_mult_216_n149, DP_mult_216_n148,
         DP_mult_216_n147, DP_mult_216_n146, DP_mult_216_n145,
         DP_mult_216_n144, DP_mult_216_n143, DP_mult_216_n142,
         DP_mult_216_n141, DP_mult_216_n140, DP_mult_216_n139,
         DP_mult_216_n138, DP_mult_216_n137, DP_mult_216_n136,
         DP_mult_216_n135, DP_mult_214_n2161, DP_mult_214_n2160,
         DP_mult_214_n2159, DP_mult_214_n2158, DP_mult_214_n2157,
         DP_mult_214_n2156, DP_mult_214_n2155, DP_mult_214_n2154,
         DP_mult_214_n2153, DP_mult_214_n2152, DP_mult_214_n2151,
         DP_mult_214_n2150, DP_mult_214_n2149, DP_mult_214_n2148,
         DP_mult_214_n2147, DP_mult_214_n2146, DP_mult_214_n2145,
         DP_mult_214_n2144, DP_mult_214_n2143, DP_mult_214_n2142,
         DP_mult_214_n2141, DP_mult_214_n2140, DP_mult_214_n2139,
         DP_mult_214_n2138, DP_mult_214_n2137, DP_mult_214_n2136,
         DP_mult_214_n2135, DP_mult_214_n2134, DP_mult_214_n2133,
         DP_mult_214_n2132, DP_mult_214_n2131, DP_mult_214_n2130,
         DP_mult_214_n2129, DP_mult_214_n2128, DP_mult_214_n2127,
         DP_mult_214_n2126, DP_mult_214_n2125, DP_mult_214_n2124,
         DP_mult_214_n2123, DP_mult_214_n2122, DP_mult_214_n2121,
         DP_mult_214_n2120, DP_mult_214_n2119, DP_mult_214_n2118,
         DP_mult_214_n2117, DP_mult_214_n2116, DP_mult_214_n2115,
         DP_mult_214_n2114, DP_mult_214_n2113, DP_mult_214_n2112,
         DP_mult_214_n2111, DP_mult_214_n2110, DP_mult_214_n2109,
         DP_mult_214_n2108, DP_mult_214_n2107, DP_mult_214_n2106,
         DP_mult_214_n2105, DP_mult_214_n2104, DP_mult_214_n2103,
         DP_mult_214_n2102, DP_mult_214_n2101, DP_mult_214_n2100,
         DP_mult_214_n2099, DP_mult_214_n2098, DP_mult_214_n2097,
         DP_mult_214_n2096, DP_mult_214_n2095, DP_mult_214_n2094,
         DP_mult_214_n2093, DP_mult_214_n2092, DP_mult_214_n2091,
         DP_mult_214_n2090, DP_mult_214_n2089, DP_mult_214_n2088,
         DP_mult_214_n2087, DP_mult_214_n2086, DP_mult_214_n2085,
         DP_mult_214_n2084, DP_mult_214_n2083, DP_mult_214_n2082,
         DP_mult_214_n2081, DP_mult_214_n2080, DP_mult_214_n2079,
         DP_mult_214_n2078, DP_mult_214_n2077, DP_mult_214_n2076,
         DP_mult_214_n2075, DP_mult_214_n2074, DP_mult_214_n2073,
         DP_mult_214_n2072, DP_mult_214_n2071, DP_mult_214_n2070,
         DP_mult_214_n2069, DP_mult_214_n2068, DP_mult_214_n2067,
         DP_mult_214_n2066, DP_mult_214_n2065, DP_mult_214_n2064,
         DP_mult_214_n2063, DP_mult_214_n2062, DP_mult_214_n2061,
         DP_mult_214_n2060, DP_mult_214_n2059, DP_mult_214_n2058,
         DP_mult_214_n2057, DP_mult_214_n2056, DP_mult_214_n2055,
         DP_mult_214_n2054, DP_mult_214_n2053, DP_mult_214_n2052,
         DP_mult_214_n2051, DP_mult_214_n2050, DP_mult_214_n2049,
         DP_mult_214_n2048, DP_mult_214_n2047, DP_mult_214_n2046,
         DP_mult_214_n2045, DP_mult_214_n2044, DP_mult_214_n2043,
         DP_mult_214_n2042, DP_mult_214_n2041, DP_mult_214_n2040,
         DP_mult_214_n2039, DP_mult_214_n2038, DP_mult_214_n2037,
         DP_mult_214_n2036, DP_mult_214_n2035, DP_mult_214_n2034,
         DP_mult_214_n2033, DP_mult_214_n2032, DP_mult_214_n2031,
         DP_mult_214_n2030, DP_mult_214_n2029, DP_mult_214_n2028,
         DP_mult_214_n2027, DP_mult_214_n2026, DP_mult_214_n2025,
         DP_mult_214_n2024, DP_mult_214_n2023, DP_mult_214_n2022,
         DP_mult_214_n2021, DP_mult_214_n2020, DP_mult_214_n2019,
         DP_mult_214_n2018, DP_mult_214_n2017, DP_mult_214_n2016,
         DP_mult_214_n2015, DP_mult_214_n2014, DP_mult_214_n2013,
         DP_mult_214_n2012, DP_mult_214_n2011, DP_mult_214_n2010,
         DP_mult_214_n2009, DP_mult_214_n2008, DP_mult_214_n2007,
         DP_mult_214_n2006, DP_mult_214_n2005, DP_mult_214_n2004,
         DP_mult_214_n2003, DP_mult_214_n2002, DP_mult_214_n2001,
         DP_mult_214_n2000, DP_mult_214_n1999, DP_mult_214_n1998,
         DP_mult_214_n1997, DP_mult_214_n1996, DP_mult_214_n1995,
         DP_mult_214_n1994, DP_mult_214_n1993, DP_mult_214_n1992,
         DP_mult_214_n1991, DP_mult_214_n1990, DP_mult_214_n1989,
         DP_mult_214_n1988, DP_mult_214_n1987, DP_mult_214_n1986,
         DP_mult_214_n1985, DP_mult_214_n1984, DP_mult_214_n1983,
         DP_mult_214_n1982, DP_mult_214_n1981, DP_mult_214_n1980,
         DP_mult_214_n1979, DP_mult_214_n1978, DP_mult_214_n1977,
         DP_mult_214_n1976, DP_mult_214_n1975, DP_mult_214_n1974,
         DP_mult_214_n1973, DP_mult_214_n1972, DP_mult_214_n1971,
         DP_mult_214_n1970, DP_mult_214_n1969, DP_mult_214_n1968,
         DP_mult_214_n1967, DP_mult_214_n1966, DP_mult_214_n1965,
         DP_mult_214_n1964, DP_mult_214_n1963, DP_mult_214_n1962,
         DP_mult_214_n1961, DP_mult_214_n1960, DP_mult_214_n1959,
         DP_mult_214_n1958, DP_mult_214_n1957, DP_mult_214_n1956,
         DP_mult_214_n1955, DP_mult_214_n1954, DP_mult_214_n1953,
         DP_mult_214_n1952, DP_mult_214_n1951, DP_mult_214_n1950,
         DP_mult_214_n1949, DP_mult_214_n1948, DP_mult_214_n1947,
         DP_mult_214_n1946, DP_mult_214_n1945, DP_mult_214_n1944,
         DP_mult_214_n1943, DP_mult_214_n1942, DP_mult_214_n1941,
         DP_mult_214_n1940, DP_mult_214_n1939, DP_mult_214_n1938,
         DP_mult_214_n1937, DP_mult_214_n1936, DP_mult_214_n1935,
         DP_mult_214_n1934, DP_mult_214_n1933, DP_mult_214_n1932,
         DP_mult_214_n1931, DP_mult_214_n1930, DP_mult_214_n1929,
         DP_mult_214_n1928, DP_mult_214_n1927, DP_mult_214_n1926,
         DP_mult_214_n1925, DP_mult_214_n1924, DP_mult_214_n1923,
         DP_mult_214_n1922, DP_mult_214_n1921, DP_mult_214_n1920,
         DP_mult_214_n1919, DP_mult_214_n1918, DP_mult_214_n1917,
         DP_mult_214_n1916, DP_mult_214_n1915, DP_mult_214_n1914,
         DP_mult_214_n1913, DP_mult_214_n1912, DP_mult_214_n1911,
         DP_mult_214_n1910, DP_mult_214_n1909, DP_mult_214_n1908,
         DP_mult_214_n1907, DP_mult_214_n1906, DP_mult_214_n1905,
         DP_mult_214_n1904, DP_mult_214_n1903, DP_mult_214_n1902,
         DP_mult_214_n1901, DP_mult_214_n1900, DP_mult_214_n1899,
         DP_mult_214_n1898, DP_mult_214_n1897, DP_mult_214_n1896,
         DP_mult_214_n1895, DP_mult_214_n1894, DP_mult_214_n1893,
         DP_mult_214_n1892, DP_mult_214_n1891, DP_mult_214_n1890,
         DP_mult_214_n1889, DP_mult_214_n1888, DP_mult_214_n1887,
         DP_mult_214_n1886, DP_mult_214_n1885, DP_mult_214_n1884,
         DP_mult_214_n1883, DP_mult_214_n1882, DP_mult_214_n1881,
         DP_mult_214_n1880, DP_mult_214_n1879, DP_mult_214_n1878,
         DP_mult_214_n1877, DP_mult_214_n1876, DP_mult_214_n1875,
         DP_mult_214_n1874, DP_mult_214_n1873, DP_mult_214_n1872,
         DP_mult_214_n1871, DP_mult_214_n1870, DP_mult_214_n1869,
         DP_mult_214_n1868, DP_mult_214_n1867, DP_mult_214_n1866,
         DP_mult_214_n1865, DP_mult_214_n1864, DP_mult_214_n1863,
         DP_mult_214_n1862, DP_mult_214_n1861, DP_mult_214_n1860,
         DP_mult_214_n1859, DP_mult_214_n1858, DP_mult_214_n1857,
         DP_mult_214_n1856, DP_mult_214_n1855, DP_mult_214_n1854,
         DP_mult_214_n1853, DP_mult_214_n1852, DP_mult_214_n1851,
         DP_mult_214_n1850, DP_mult_214_n1849, DP_mult_214_n1848,
         DP_mult_214_n1847, DP_mult_214_n1846, DP_mult_214_n1845,
         DP_mult_214_n1844, DP_mult_214_n1843, DP_mult_214_n1842,
         DP_mult_214_n1841, DP_mult_214_n1840, DP_mult_214_n1839,
         DP_mult_214_n1838, DP_mult_214_n1837, DP_mult_214_n1836,
         DP_mult_214_n1835, DP_mult_214_n1834, DP_mult_214_n1833,
         DP_mult_214_n1832, DP_mult_214_n1831, DP_mult_214_n1830,
         DP_mult_214_n1829, DP_mult_214_n1828, DP_mult_214_n1827,
         DP_mult_214_n1826, DP_mult_214_n1825, DP_mult_214_n1824,
         DP_mult_214_n1823, DP_mult_214_n1822, DP_mult_214_n1821,
         DP_mult_214_n1820, DP_mult_214_n1819, DP_mult_214_n1818,
         DP_mult_214_n1817, DP_mult_214_n1816, DP_mult_214_n1815,
         DP_mult_214_n1814, DP_mult_214_n1813, DP_mult_214_n1812,
         DP_mult_214_n1811, DP_mult_214_n1810, DP_mult_214_n1809,
         DP_mult_214_n1808, DP_mult_214_n1807, DP_mult_214_n1806,
         DP_mult_214_n1805, DP_mult_214_n1804, DP_mult_214_n1803,
         DP_mult_214_n1802, DP_mult_214_n1801, DP_mult_214_n1800,
         DP_mult_214_n1799, DP_mult_214_n1798, DP_mult_214_n1797,
         DP_mult_214_n1796, DP_mult_214_n1795, DP_mult_214_n1794,
         DP_mult_214_n1793, DP_mult_214_n1792, DP_mult_214_n1791,
         DP_mult_214_n1790, DP_mult_214_n1789, DP_mult_214_n1788,
         DP_mult_214_n1787, DP_mult_214_n1786, DP_mult_214_n1785,
         DP_mult_214_n1784, DP_mult_214_n1783, DP_mult_214_n1782,
         DP_mult_214_n1781, DP_mult_214_n1780, DP_mult_214_n1779,
         DP_mult_214_n1778, DP_mult_214_n1777, DP_mult_214_n1776,
         DP_mult_214_n1775, DP_mult_214_n1774, DP_mult_214_n1773,
         DP_mult_214_n1772, DP_mult_214_n1771, DP_mult_214_n1770,
         DP_mult_214_n1769, DP_mult_214_n1768, DP_mult_214_n1767,
         DP_mult_214_n1766, DP_mult_214_n1765, DP_mult_214_n1764,
         DP_mult_214_n1763, DP_mult_214_n1762, DP_mult_214_n1761,
         DP_mult_214_n1760, DP_mult_214_n1759, DP_mult_214_n1758,
         DP_mult_214_n1757, DP_mult_214_n1756, DP_mult_214_n1755,
         DP_mult_214_n1754, DP_mult_214_n1753, DP_mult_214_n1752,
         DP_mult_214_n1751, DP_mult_214_n1750, DP_mult_214_n1749,
         DP_mult_214_n1748, DP_mult_214_n1747, DP_mult_214_n1746,
         DP_mult_214_n1745, DP_mult_214_n1744, DP_mult_214_n1743,
         DP_mult_214_n1742, DP_mult_214_n1741, DP_mult_214_n1740,
         DP_mult_214_n1739, DP_mult_214_n1738, DP_mult_214_n1737,
         DP_mult_214_n1736, DP_mult_214_n1735, DP_mult_214_n1734,
         DP_mult_214_n1733, DP_mult_214_n1732, DP_mult_214_n1731,
         DP_mult_214_n1730, DP_mult_214_n1729, DP_mult_214_n1728,
         DP_mult_214_n1727, DP_mult_214_n1726, DP_mult_214_n1725,
         DP_mult_214_n1724, DP_mult_214_n1723, DP_mult_214_n1722,
         DP_mult_214_n1721, DP_mult_214_n1720, DP_mult_214_n1719,
         DP_mult_214_n1718, DP_mult_214_n1717, DP_mult_214_n1716,
         DP_mult_214_n1715, DP_mult_214_n1714, DP_mult_214_n1713,
         DP_mult_214_n1712, DP_mult_214_n1711, DP_mult_214_n1710,
         DP_mult_214_n1709, DP_mult_214_n1708, DP_mult_214_n1707,
         DP_mult_214_n1706, DP_mult_214_n1705, DP_mult_214_n1704,
         DP_mult_214_n1703, DP_mult_214_n1702, DP_mult_214_n1701,
         DP_mult_214_n1700, DP_mult_214_n1699, DP_mult_214_n1698,
         DP_mult_214_n1697, DP_mult_214_n1696, DP_mult_214_n1695,
         DP_mult_214_n1694, DP_mult_214_n1693, DP_mult_214_n1692,
         DP_mult_214_n1691, DP_mult_214_n1690, DP_mult_214_n1689,
         DP_mult_214_n1688, DP_mult_214_n1687, DP_mult_214_n1686,
         DP_mult_214_n1685, DP_mult_214_n1684, DP_mult_214_n1683,
         DP_mult_214_n1682, DP_mult_214_n1681, DP_mult_214_n1680,
         DP_mult_214_n1679, DP_mult_214_n1678, DP_mult_214_n1677,
         DP_mult_214_n1676, DP_mult_214_n1675, DP_mult_214_n1674,
         DP_mult_214_n1673, DP_mult_214_n1672, DP_mult_214_n1671,
         DP_mult_214_n1670, DP_mult_214_n1669, DP_mult_214_n1668,
         DP_mult_214_n1667, DP_mult_214_n1666, DP_mult_214_n1665,
         DP_mult_214_n1664, DP_mult_214_n1663, DP_mult_214_n1662,
         DP_mult_214_n1661, DP_mult_214_n1660, DP_mult_214_n1659,
         DP_mult_214_n1658, DP_mult_214_n1657, DP_mult_214_n1656,
         DP_mult_214_n1655, DP_mult_214_n1654, DP_mult_214_n1653,
         DP_mult_214_n1652, DP_mult_214_n1651, DP_mult_214_n1650,
         DP_mult_214_n1649, DP_mult_214_n1648, DP_mult_214_n1647,
         DP_mult_214_n1646, DP_mult_214_n1645, DP_mult_214_n1644,
         DP_mult_214_n1643, DP_mult_214_n1642, DP_mult_214_n1641,
         DP_mult_214_n1640, DP_mult_214_n1639, DP_mult_214_n1638,
         DP_mult_214_n1637, DP_mult_214_n1636, DP_mult_214_n1635,
         DP_mult_214_n1634, DP_mult_214_n1633, DP_mult_214_n1632,
         DP_mult_214_n1631, DP_mult_214_n1630, DP_mult_214_n1629,
         DP_mult_214_n1628, DP_mult_214_n1627, DP_mult_214_n1626,
         DP_mult_214_n1625, DP_mult_214_n1624, DP_mult_214_n1623,
         DP_mult_214_n1622, DP_mult_214_n1621, DP_mult_214_n1620,
         DP_mult_214_n1619, DP_mult_214_n1618, DP_mult_214_n1617,
         DP_mult_214_n1616, DP_mult_214_n1615, DP_mult_214_n1614,
         DP_mult_214_n1613, DP_mult_214_n1612, DP_mult_214_n1611,
         DP_mult_214_n1610, DP_mult_214_n1609, DP_mult_214_n1608,
         DP_mult_214_n1607, DP_mult_214_n1606, DP_mult_214_n1605,
         DP_mult_214_n1604, DP_mult_214_n1603, DP_mult_214_n1602,
         DP_mult_214_n1601, DP_mult_214_n1600, DP_mult_214_n1599,
         DP_mult_214_n1598, DP_mult_214_n1597, DP_mult_214_n1596,
         DP_mult_214_n1595, DP_mult_214_n1594, DP_mult_214_n1593,
         DP_mult_214_n1592, DP_mult_214_n1591, DP_mult_214_n1590,
         DP_mult_214_n1589, DP_mult_214_n1588, DP_mult_214_n1587,
         DP_mult_214_n1586, DP_mult_214_n1585, DP_mult_214_n1584,
         DP_mult_214_n1583, DP_mult_214_n1582, DP_mult_214_n1581,
         DP_mult_214_n1580, DP_mult_214_n1579, DP_mult_214_n1578,
         DP_mult_214_n1577, DP_mult_214_n1576, DP_mult_214_n1575,
         DP_mult_214_n1574, DP_mult_214_n1573, DP_mult_214_n1572,
         DP_mult_214_n1571, DP_mult_214_n1570, DP_mult_214_n1569,
         DP_mult_214_n1568, DP_mult_214_n1567, DP_mult_214_n1566,
         DP_mult_214_n1565, DP_mult_214_n1564, DP_mult_214_n1563,
         DP_mult_214_n1562, DP_mult_214_n1561, DP_mult_214_n1560,
         DP_mult_214_n1559, DP_mult_214_n1558, DP_mult_214_n1557,
         DP_mult_214_n1556, DP_mult_214_n1555, DP_mult_214_n1554,
         DP_mult_214_n1553, DP_mult_214_n1552, DP_mult_214_n1551,
         DP_mult_214_n1550, DP_mult_214_n1549, DP_mult_214_n1548,
         DP_mult_214_n1547, DP_mult_214_n1546, DP_mult_214_n1545,
         DP_mult_214_n1544, DP_mult_214_n1543, DP_mult_214_n1542,
         DP_mult_214_n1541, DP_mult_214_n1540, DP_mult_214_n1539,
         DP_mult_214_n1538, DP_mult_214_n1537, DP_mult_214_n1536,
         DP_mult_214_n1535, DP_mult_214_n1534, DP_mult_214_n1533,
         DP_mult_214_n1397, DP_mult_214_n1396, DP_mult_214_n1395,
         DP_mult_214_n1394, DP_mult_214_n1393, DP_mult_214_n1392,
         DP_mult_214_n1391, DP_mult_214_n1390, DP_mult_214_n1389,
         DP_mult_214_n1388, DP_mult_214_n1387, DP_mult_214_n1386,
         DP_mult_214_n1385, DP_mult_214_n1384, DP_mult_214_n1383,
         DP_mult_214_n1382, DP_mult_214_n1381, DP_mult_214_n1380,
         DP_mult_214_n1379, DP_mult_214_n1378, DP_mult_214_n1377,
         DP_mult_214_n1376, DP_mult_214_n1375, DP_mult_214_n1374,
         DP_mult_214_n908, DP_mult_214_n907, DP_mult_214_n906,
         DP_mult_214_n904, DP_mult_214_n903, DP_mult_214_n902,
         DP_mult_214_n901, DP_mult_214_n900, DP_mult_214_n899,
         DP_mult_214_n898, DP_mult_214_n897, DP_mult_214_n896,
         DP_mult_214_n895, DP_mult_214_n894, DP_mult_214_n893,
         DP_mult_214_n892, DP_mult_214_n891, DP_mult_214_n890,
         DP_mult_214_n889, DP_mult_214_n888, DP_mult_214_n887,
         DP_mult_214_n886, DP_mult_214_n885, DP_mult_214_n884,
         DP_mult_214_n883, DP_mult_214_n882, DP_mult_214_n881,
         DP_mult_214_n880, DP_mult_214_n879, DP_mult_214_n878,
         DP_mult_214_n877, DP_mult_214_n876, DP_mult_214_n875,
         DP_mult_214_n874, DP_mult_214_n873, DP_mult_214_n872,
         DP_mult_214_n871, DP_mult_214_n870, DP_mult_214_n869,
         DP_mult_214_n868, DP_mult_214_n867, DP_mult_214_n866,
         DP_mult_214_n865, DP_mult_214_n864, DP_mult_214_n863,
         DP_mult_214_n862, DP_mult_214_n861, DP_mult_214_n860,
         DP_mult_214_n859, DP_mult_214_n858, DP_mult_214_n857,
         DP_mult_214_n856, DP_mult_214_n855, DP_mult_214_n854,
         DP_mult_214_n853, DP_mult_214_n852, DP_mult_214_n851,
         DP_mult_214_n850, DP_mult_214_n849, DP_mult_214_n848,
         DP_mult_214_n847, DP_mult_214_n846, DP_mult_214_n845,
         DP_mult_214_n844, DP_mult_214_n843, DP_mult_214_n842,
         DP_mult_214_n841, DP_mult_214_n840, DP_mult_214_n839,
         DP_mult_214_n838, DP_mult_214_n837, DP_mult_214_n836,
         DP_mult_214_n835, DP_mult_214_n834, DP_mult_214_n833,
         DP_mult_214_n832, DP_mult_214_n831, DP_mult_214_n830,
         DP_mult_214_n829, DP_mult_214_n828, DP_mult_214_n827,
         DP_mult_214_n826, DP_mult_214_n825, DP_mult_214_n824,
         DP_mult_214_n823, DP_mult_214_n822, DP_mult_214_n821,
         DP_mult_214_n820, DP_mult_214_n819, DP_mult_214_n818,
         DP_mult_214_n817, DP_mult_214_n816, DP_mult_214_n815,
         DP_mult_214_n814, DP_mult_214_n813, DP_mult_214_n812,
         DP_mult_214_n811, DP_mult_214_n810, DP_mult_214_n809,
         DP_mult_214_n808, DP_mult_214_n807, DP_mult_214_n806,
         DP_mult_214_n805, DP_mult_214_n804, DP_mult_214_n803,
         DP_mult_214_n802, DP_mult_214_n801, DP_mult_214_n800,
         DP_mult_214_n799, DP_mult_214_n798, DP_mult_214_n797,
         DP_mult_214_n796, DP_mult_214_n795, DP_mult_214_n794,
         DP_mult_214_n793, DP_mult_214_n792, DP_mult_214_n791,
         DP_mult_214_n790, DP_mult_214_n789, DP_mult_214_n788,
         DP_mult_214_n787, DP_mult_214_n786, DP_mult_214_n785,
         DP_mult_214_n784, DP_mult_214_n783, DP_mult_214_n782,
         DP_mult_214_n781, DP_mult_214_n780, DP_mult_214_n779,
         DP_mult_214_n778, DP_mult_214_n777, DP_mult_214_n776,
         DP_mult_214_n775, DP_mult_214_n774, DP_mult_214_n773,
         DP_mult_214_n772, DP_mult_214_n771, DP_mult_214_n770,
         DP_mult_214_n769, DP_mult_214_n768, DP_mult_214_n767,
         DP_mult_214_n766, DP_mult_214_n765, DP_mult_214_n764,
         DP_mult_214_n763, DP_mult_214_n762, DP_mult_214_n761,
         DP_mult_214_n760, DP_mult_214_n759, DP_mult_214_n758,
         DP_mult_214_n757, DP_mult_214_n756, DP_mult_214_n755,
         DP_mult_214_n754, DP_mult_214_n753, DP_mult_214_n752,
         DP_mult_214_n751, DP_mult_214_n750, DP_mult_214_n749,
         DP_mult_214_n748, DP_mult_214_n747, DP_mult_214_n746,
         DP_mult_214_n745, DP_mult_214_n744, DP_mult_214_n743,
         DP_mult_214_n742, DP_mult_214_n741, DP_mult_214_n740,
         DP_mult_214_n739, DP_mult_214_n738, DP_mult_214_n737,
         DP_mult_214_n736, DP_mult_214_n735, DP_mult_214_n734,
         DP_mult_214_n733, DP_mult_214_n732, DP_mult_214_n731,
         DP_mult_214_n730, DP_mult_214_n729, DP_mult_214_n727,
         DP_mult_214_n726, DP_mult_214_n725, DP_mult_214_n724,
         DP_mult_214_n723, DP_mult_214_n722, DP_mult_214_n721,
         DP_mult_214_n720, DP_mult_214_n719, DP_mult_214_n718,
         DP_mult_214_n717, DP_mult_214_n716, DP_mult_214_n715,
         DP_mult_214_n714, DP_mult_214_n713, DP_mult_214_n712,
         DP_mult_214_n711, DP_mult_214_n710, DP_mult_214_n709,
         DP_mult_214_n708, DP_mult_214_n707, DP_mult_214_n706,
         DP_mult_214_n688, DP_mult_214_n687, DP_mult_214_n686,
         DP_mult_214_n685, DP_mult_214_n684, DP_mult_214_n683,
         DP_mult_214_n682, DP_mult_214_n681, DP_mult_214_n680,
         DP_mult_214_n679, DP_mult_214_n678, DP_mult_214_n677,
         DP_mult_214_n676, DP_mult_214_n675, DP_mult_214_n674,
         DP_mult_214_n673, DP_mult_214_n672, DP_mult_214_n671,
         DP_mult_214_n670, DP_mult_214_n669, DP_mult_214_n668,
         DP_mult_214_n667, DP_mult_214_n666, DP_mult_214_n665,
         DP_mult_214_n664, DP_mult_214_n663, DP_mult_214_n662,
         DP_mult_214_n661, DP_mult_214_n660, DP_mult_214_n659,
         DP_mult_214_n658, DP_mult_214_n657, DP_mult_214_n656,
         DP_mult_214_n655, DP_mult_214_n654, DP_mult_214_n653,
         DP_mult_214_n652, DP_mult_214_n651, DP_mult_214_n650,
         DP_mult_214_n649, DP_mult_214_n648, DP_mult_214_n647,
         DP_mult_214_n646, DP_mult_214_n645, DP_mult_214_n644,
         DP_mult_214_n643, DP_mult_214_n642, DP_mult_214_n641,
         DP_mult_214_n640, DP_mult_214_n639, DP_mult_214_n638,
         DP_mult_214_n637, DP_mult_214_n636, DP_mult_214_n635,
         DP_mult_214_n634, DP_mult_214_n633, DP_mult_214_n632,
         DP_mult_214_n631, DP_mult_214_n630, DP_mult_214_n629,
         DP_mult_214_n628, DP_mult_214_n627, DP_mult_214_n626,
         DP_mult_214_n625, DP_mult_214_n624, DP_mult_214_n623,
         DP_mult_214_n622, DP_mult_214_n621, DP_mult_214_n620,
         DP_mult_214_n619, DP_mult_214_n618, DP_mult_214_n617,
         DP_mult_214_n616, DP_mult_214_n615, DP_mult_214_n614,
         DP_mult_214_n613, DP_mult_214_n612, DP_mult_214_n611,
         DP_mult_214_n610, DP_mult_214_n609, DP_mult_214_n608,
         DP_mult_214_n607, DP_mult_214_n606, DP_mult_214_n605,
         DP_mult_214_n604, DP_mult_214_n603, DP_mult_214_n602,
         DP_mult_214_n601, DP_mult_214_n600, DP_mult_214_n599,
         DP_mult_214_n598, DP_mult_214_n597, DP_mult_214_n596,
         DP_mult_214_n595, DP_mult_214_n594, DP_mult_214_n593,
         DP_mult_214_n592, DP_mult_214_n591, DP_mult_214_n590,
         DP_mult_214_n589, DP_mult_214_n588, DP_mult_214_n587,
         DP_mult_214_n586, DP_mult_214_n585, DP_mult_214_n584,
         DP_mult_214_n583, DP_mult_214_n582, DP_mult_214_n581,
         DP_mult_214_n580, DP_mult_214_n579, DP_mult_214_n578,
         DP_mult_214_n577, DP_mult_214_n576, DP_mult_214_n575,
         DP_mult_214_n574, DP_mult_214_n573, DP_mult_214_n572,
         DP_mult_214_n571, DP_mult_214_n570, DP_mult_214_n569,
         DP_mult_214_n568, DP_mult_214_n567, DP_mult_214_n566,
         DP_mult_214_n565, DP_mult_214_n564, DP_mult_214_n563,
         DP_mult_214_n562, DP_mult_214_n561, DP_mult_214_n560,
         DP_mult_214_n559, DP_mult_214_n558, DP_mult_214_n557,
         DP_mult_214_n556, DP_mult_214_n555, DP_mult_214_n554,
         DP_mult_214_n553, DP_mult_214_n552, DP_mult_214_n551,
         DP_mult_214_n550, DP_mult_214_n549, DP_mult_214_n548,
         DP_mult_214_n547, DP_mult_214_n546, DP_mult_214_n545,
         DP_mult_214_n544, DP_mult_214_n543, DP_mult_214_n542,
         DP_mult_214_n541, DP_mult_214_n540, DP_mult_214_n539,
         DP_mult_214_n538, DP_mult_214_n537, DP_mult_214_n536,
         DP_mult_214_n535, DP_mult_214_n534, DP_mult_214_n533,
         DP_mult_214_n532, DP_mult_214_n531, DP_mult_214_n530,
         DP_mult_214_n529, DP_mult_214_n528, DP_mult_214_n527,
         DP_mult_214_n526, DP_mult_214_n525, DP_mult_214_n524,
         DP_mult_214_n523, DP_mult_214_n522, DP_mult_214_n521,
         DP_mult_214_n520, DP_mult_214_n519, DP_mult_214_n518,
         DP_mult_214_n517, DP_mult_214_n516, DP_mult_214_n515,
         DP_mult_214_n514, DP_mult_214_n513, DP_mult_214_n512,
         DP_mult_214_n511, DP_mult_214_n510, DP_mult_214_n509,
         DP_mult_214_n508, DP_mult_214_n507, DP_mult_214_n506,
         DP_mult_214_n505, DP_mult_214_n504, DP_mult_214_n503,
         DP_mult_214_n502, DP_mult_214_n501, DP_mult_214_n500,
         DP_mult_214_n499, DP_mult_214_n498, DP_mult_214_n497,
         DP_mult_214_n496, DP_mult_214_n495, DP_mult_214_n494,
         DP_mult_214_n493, DP_mult_214_n492, DP_mult_214_n491,
         DP_mult_214_n490, DP_mult_214_n489, DP_mult_214_n488,
         DP_mult_214_n487, DP_mult_214_n486, DP_mult_214_n485,
         DP_mult_214_n484, DP_mult_214_n483, DP_mult_214_n482,
         DP_mult_214_n481, DP_mult_214_n479, DP_mult_214_n478,
         DP_mult_214_n477, DP_mult_214_n476, DP_mult_214_n475,
         DP_mult_214_n474, DP_mult_214_n473, DP_mult_214_n472,
         DP_mult_214_n471, DP_mult_214_n470, DP_mult_214_n469,
         DP_mult_214_n468, DP_mult_214_n467, DP_mult_214_n466,
         DP_mult_214_n465, DP_mult_214_n464, DP_mult_214_n463,
         DP_mult_214_n462, DP_mult_214_n461, DP_mult_214_n460,
         DP_mult_214_n459, DP_mult_214_n458, DP_mult_214_n457,
         DP_mult_214_n456, DP_mult_214_n455, DP_mult_214_n454,
         DP_mult_214_n453, DP_mult_214_n452, DP_mult_214_n451,
         DP_mult_214_n450, DP_mult_214_n449, DP_mult_214_n448,
         DP_mult_214_n447, DP_mult_214_n446, DP_mult_214_n445,
         DP_mult_214_n444, DP_mult_214_n442, DP_mult_214_n441,
         DP_mult_214_n440, DP_mult_214_n439, DP_mult_214_n438,
         DP_mult_214_n437, DP_mult_214_n436, DP_mult_214_n435,
         DP_mult_214_n434, DP_mult_214_n433, DP_mult_214_n432,
         DP_mult_214_n431, DP_mult_214_n430, DP_mult_214_n429,
         DP_mult_214_n428, DP_mult_214_n427, DP_mult_214_n426,
         DP_mult_214_n425, DP_mult_214_n424, DP_mult_214_n423,
         DP_mult_214_n422, DP_mult_214_n421, DP_mult_214_n420,
         DP_mult_214_n419, DP_mult_214_n418, DP_mult_214_n417,
         DP_mult_214_n416, DP_mult_214_n415, DP_mult_214_n414,
         DP_mult_214_n413, DP_mult_214_n411, DP_mult_214_n410,
         DP_mult_214_n409, DP_mult_214_n408, DP_mult_214_n407,
         DP_mult_214_n406, DP_mult_214_n405, DP_mult_214_n404,
         DP_mult_214_n403, DP_mult_214_n402, DP_mult_214_n401,
         DP_mult_214_n400, DP_mult_214_n399, DP_mult_214_n398,
         DP_mult_214_n397, DP_mult_214_n396, DP_mult_214_n395,
         DP_mult_214_n394, DP_mult_214_n393, DP_mult_214_n392,
         DP_mult_214_n391, DP_mult_214_n390, DP_mult_214_n389,
         DP_mult_214_n387, DP_mult_214_n386, DP_mult_214_n385,
         DP_mult_214_n384, DP_mult_214_n383, DP_mult_214_n382,
         DP_mult_214_n381, DP_mult_214_n380, DP_mult_214_n379,
         DP_mult_214_n378, DP_mult_214_n377, DP_mult_214_n376,
         DP_mult_214_n375, DP_mult_214_n374, DP_mult_214_n373,
         DP_mult_214_n372, DP_mult_214_n371, DP_mult_214_n370,
         DP_mult_214_n368, DP_mult_214_n367, DP_mult_214_n366,
         DP_mult_214_n365, DP_mult_214_n364, DP_mult_214_n363,
         DP_mult_214_n362, DP_mult_214_n361, DP_mult_214_n360,
         DP_mult_214_n359, DP_mult_214_n358, DP_mult_214_n356,
         DP_mult_214_n355, DP_mult_214_n354, DP_mult_214_n353,
         DP_mult_214_n352, DP_mult_214_n351, DP_mult_214_n326,
         DP_mult_214_n325, DP_mult_214_n324, DP_mult_214_n323,
         DP_mult_214_n322, DP_mult_214_n321, DP_mult_214_n320,
         DP_mult_214_n319, DP_mult_214_n318, DP_mult_214_n317,
         DP_mult_214_n316, DP_mult_214_n315, DP_mult_214_n314,
         DP_mult_214_n313, DP_mult_214_n312, DP_mult_214_n311,
         DP_mult_214_n310, DP_mult_214_n309, DP_mult_214_n308,
         DP_mult_214_n307, DP_mult_214_n306, DP_mult_214_n305,
         DP_mult_214_n304, DP_mult_214_n303, DP_mult_207_n249,
         DP_mult_207_n248, DP_mult_207_n247, DP_mult_207_n246,
         DP_mult_207_n245, DP_mult_207_n244, DP_mult_207_n243,
         DP_mult_207_n242, DP_mult_207_n241, DP_mult_207_n240,
         DP_mult_207_n239, DP_mult_207_n10, DP_mult_207_n100, DP_mult_207_n101,
         DP_mult_207_n102, DP_mult_207_n103, DP_mult_207_n104,
         DP_mult_207_n105, DP_mult_207_n106, DP_mult_207_n107,
         DP_mult_207_n108, DP_mult_207_n109, DP_mult_207_n11, DP_mult_207_n110,
         DP_mult_207_n111, DP_mult_207_n112, DP_mult_207_n113,
         DP_mult_207_n114, DP_mult_207_n115, DP_mult_207_n116,
         DP_mult_207_n117, DP_mult_207_n118, DP_mult_207_n119, DP_mult_207_n12,
         DP_mult_207_n120, DP_mult_207_n121, DP_mult_207_n122,
         DP_mult_207_n123, DP_mult_207_n124, DP_mult_207_n125,
         DP_mult_207_n126, DP_mult_207_n127, DP_mult_207_n128,
         DP_mult_207_n129, DP_mult_207_n13, DP_mult_207_n130, DP_mult_207_n131,
         DP_mult_207_n132, DP_mult_207_n133, DP_mult_207_n134,
         DP_mult_207_n135, DP_mult_207_n136, DP_mult_207_n137,
         DP_mult_207_n138, DP_mult_207_n139, DP_mult_207_n14, DP_mult_207_n140,
         DP_mult_207_n141, DP_mult_207_n142, DP_mult_207_n143,
         DP_mult_207_n144, DP_mult_207_n145, DP_mult_207_n146,
         DP_mult_207_n147, DP_mult_207_n148, DP_mult_207_n149, DP_mult_207_n15,
         DP_mult_207_n150, DP_mult_207_n151, DP_mult_207_n152,
         DP_mult_207_n153, DP_mult_207_n154, DP_mult_207_n155,
         DP_mult_207_n156, DP_mult_207_n158, DP_mult_207_n159, DP_mult_207_n16,
         DP_mult_207_n160, DP_mult_207_n161, DP_mult_207_n162,
         DP_mult_207_n163, DP_mult_207_n164, DP_mult_207_n165,
         DP_mult_207_n166, DP_mult_207_n167, DP_mult_207_n168,
         DP_mult_207_n169, DP_mult_207_n17, DP_mult_207_n170, DP_mult_207_n171,
         DP_mult_207_n172, DP_mult_207_n173, DP_mult_207_n174,
         DP_mult_207_n175, DP_mult_207_n176, DP_mult_207_n177, DP_mult_207_n18,
         DP_mult_207_n19, DP_mult_207_n2, DP_mult_207_n20, DP_mult_207_n21,
         DP_mult_207_n22, DP_mult_207_n23, DP_mult_207_n24, DP_mult_207_n25,
         DP_mult_207_n26, DP_mult_207_n27, DP_mult_207_n28, DP_mult_207_n29,
         DP_mult_207_n3, DP_mult_207_n30, DP_mult_207_n31, DP_mult_207_n32,
         DP_mult_207_n33, DP_mult_207_n34, DP_mult_207_n35, DP_mult_207_n36,
         DP_mult_207_n37, DP_mult_207_n38, DP_mult_207_n39, DP_mult_207_n4,
         DP_mult_207_n40, DP_mult_207_n41, DP_mult_207_n42, DP_mult_207_n43,
         DP_mult_207_n44, DP_mult_207_n45, DP_mult_207_n46, DP_mult_207_n47,
         DP_mult_207_n48, DP_mult_207_n49, DP_mult_207_n5, DP_mult_207_n50,
         DP_mult_207_n51, DP_mult_207_n52, DP_mult_207_n53, DP_mult_207_n54,
         DP_mult_207_n55, DP_mult_207_n56, DP_mult_207_n57, DP_mult_207_n58,
         DP_mult_207_n59, DP_mult_207_n6, DP_mult_207_n60, DP_mult_207_n61,
         DP_mult_207_n62, DP_mult_207_n63, DP_mult_207_n64, DP_mult_207_n65,
         DP_mult_207_n66, DP_mult_207_n67, DP_mult_207_n68, DP_mult_207_n69,
         DP_mult_207_n7, DP_mult_207_n71, DP_mult_207_n72, DP_mult_207_n73,
         DP_mult_207_n74, DP_mult_207_n75, DP_mult_207_n76, DP_mult_207_n77,
         DP_mult_207_n78, DP_mult_207_n79, DP_mult_207_n8, DP_mult_207_n80,
         DP_mult_207_n81, DP_mult_207_n82, DP_mult_207_n83, DP_mult_207_n84,
         DP_mult_207_n85, DP_mult_207_n86, DP_mult_207_n87, DP_mult_207_n88,
         DP_mult_207_n89, DP_mult_207_n9, DP_mult_207_n90, DP_mult_207_n91,
         DP_mult_207_n92, DP_mult_207_n93, DP_mult_207_n94, DP_mult_207_n95,
         DP_mult_207_n96, DP_mult_207_n97, DP_mult_207_n98, DP_mult_207_n99,
         DP_mult_207_n1, DP_sub_0_root_add_0_root_add_207_B_not_2_,
         DP_sub_0_root_add_0_root_add_207_B_not_3_,
         DP_sub_0_root_add_0_root_add_207_B_not_4_,
         DP_sub_0_root_add_0_root_add_207_B_not_5_,
         DP_sub_0_root_add_0_root_add_207_B_not_6_,
         DP_sub_0_root_add_0_root_add_207_B_not_7_,
         DP_sub_0_root_add_0_root_add_207_B_not_8_,
         DP_sub_0_root_add_0_root_add_207_B_not_9_,
         DP_sub_0_root_add_0_root_add_207_B_not_10_,
         DP_sub_0_root_add_0_root_add_207_B_not_11_,
         DP_sub_0_root_add_0_root_add_207_B_not_12_,
         DP_sub_0_root_add_0_root_add_207_B_not_13_,
         DP_sub_0_root_add_0_root_add_207_B_not_14_,
         DP_sub_0_root_add_0_root_add_207_B_not_15_,
         DP_sub_0_root_add_0_root_add_207_B_not_16_,
         DP_sub_0_root_add_0_root_add_207_B_not_17_,
         DP_sub_0_root_add_0_root_add_207_B_not_18_,
         DP_sub_0_root_add_0_root_add_207_B_not_19_,
         DP_sub_0_root_add_0_root_add_207_B_not_20_,
         DP_sub_0_root_add_0_root_add_207_B_not_21_,
         DP_sub_0_root_add_0_root_add_207_B_not_22_,
         DP_sub_0_root_add_0_root_add_207_B_not_23_,
         DP_sub_0_root_add_0_root_add_207_carry_2_,
         DP_sub_0_root_add_0_root_add_207_carry_3_,
         DP_sub_0_root_add_0_root_add_207_carry_4_,
         DP_sub_0_root_add_0_root_add_207_carry_5_,
         DP_sub_0_root_add_0_root_add_207_carry_6_,
         DP_sub_0_root_add_0_root_add_207_carry_7_,
         DP_sub_0_root_add_0_root_add_207_carry_8_,
         DP_sub_0_root_add_0_root_add_207_carry_9_,
         DP_sub_0_root_add_0_root_add_207_carry_10_,
         DP_sub_0_root_add_0_root_add_207_carry_11_,
         DP_sub_0_root_add_0_root_add_207_carry_12_,
         DP_sub_0_root_add_0_root_add_207_carry_13_,
         DP_sub_0_root_add_0_root_add_207_carry_14_,
         DP_sub_0_root_add_0_root_add_207_carry_15_,
         DP_sub_0_root_add_0_root_add_207_carry_16_,
         DP_sub_0_root_add_0_root_add_207_carry_17_,
         DP_sub_0_root_add_0_root_add_207_carry_18_,
         DP_sub_0_root_add_0_root_add_207_carry_19_,
         DP_sub_0_root_add_0_root_add_207_carry_20_,
         DP_sub_0_root_add_0_root_add_207_carry_21_,
         DP_sub_0_root_add_0_root_add_207_carry_22_,
         DP_sub_0_root_add_0_root_add_207_carry_23_, DP_mult_208_n626,
         DP_mult_208_n625, DP_mult_208_n624, DP_mult_208_n623,
         DP_mult_208_n622, DP_mult_208_n621, DP_mult_208_n620,
         DP_mult_208_n619, DP_mult_208_n618, DP_mult_208_n617,
         DP_mult_208_n616, DP_mult_208_n615, DP_mult_208_n614,
         DP_mult_208_n613, DP_mult_208_n612, DP_mult_208_n611,
         DP_mult_208_n610, DP_mult_208_n609, DP_mult_208_n608,
         DP_mult_208_n607, DP_mult_208_n606, DP_mult_208_n605,
         DP_mult_208_n604, DP_mult_208_n603, DP_mult_208_n602,
         DP_mult_208_n601, DP_mult_208_n600, DP_mult_208_n599,
         DP_mult_208_n598, DP_mult_208_n597, DP_mult_208_n596,
         DP_mult_208_n595, DP_mult_208_n594, DP_mult_208_n593,
         DP_mult_208_n592, DP_mult_208_n591, DP_mult_208_n590,
         DP_mult_208_n589, DP_mult_208_n588, DP_mult_208_n587,
         DP_mult_208_n586, DP_mult_208_n585, DP_mult_208_n584,
         DP_mult_208_n583, DP_mult_208_n582, DP_mult_208_n581,
         DP_mult_208_n580, DP_mult_208_n579, DP_mult_208_n578,
         DP_mult_208_n577, DP_mult_208_n576, DP_mult_208_n575,
         DP_mult_208_n574, DP_mult_208_n573, DP_mult_208_n572,
         DP_mult_208_n571, DP_mult_208_n570, DP_mult_208_n569,
         DP_mult_208_n568, DP_mult_208_n567, DP_mult_208_n566,
         DP_mult_208_n565, DP_mult_208_n564, DP_mult_208_n563,
         DP_mult_208_n562, DP_mult_208_n561, DP_mult_208_n560,
         DP_mult_208_n559, DP_mult_208_n558, DP_mult_208_n557,
         DP_mult_208_n556, DP_mult_208_n555, DP_mult_208_n554,
         DP_mult_208_n553, DP_mult_208_n552, DP_mult_208_n551,
         DP_mult_208_n550, DP_mult_208_n549, DP_mult_208_n548,
         DP_mult_208_n547, DP_mult_208_n546, DP_mult_208_n545,
         DP_mult_208_n544, DP_mult_208_n543, DP_mult_208_n542,
         DP_mult_208_n541, DP_mult_208_n540, DP_mult_208_n539,
         DP_mult_208_n538, DP_mult_208_n537, DP_mult_208_n536,
         DP_mult_208_n535, DP_mult_208_n534, DP_mult_208_n533,
         DP_mult_208_n532, DP_mult_208_n531, DP_mult_208_n530,
         DP_mult_208_n529, DP_mult_208_n528, DP_mult_208_n527,
         DP_mult_208_n526, DP_mult_208_n525, DP_mult_208_n524,
         DP_mult_208_n523, DP_mult_208_n522, DP_mult_208_n521,
         DP_mult_208_n520, DP_mult_208_n519, DP_mult_208_n518,
         DP_mult_208_n517, DP_mult_208_n516, DP_mult_208_n515,
         DP_mult_208_n514, DP_mult_208_n513, DP_mult_208_n329,
         DP_mult_208_n328, DP_mult_208_n327, DP_mult_208_n326,
         DP_mult_208_n325, DP_mult_208_n324, DP_mult_208_n323,
         DP_mult_208_n322, DP_mult_208_n321, DP_mult_208_n320,
         DP_mult_208_n319, DP_mult_208_n318, DP_mult_208_n317,
         DP_mult_208_n316, DP_mult_208_n315, DP_mult_208_n314,
         DP_mult_208_n313, DP_mult_208_n312, DP_mult_208_n311,
         DP_mult_208_n310, DP_mult_208_n309, DP_mult_208_n308,
         DP_mult_208_n307, DP_mult_208_n306, DP_mult_208_n305,
         DP_mult_208_n304, DP_mult_208_n303, DP_mult_208_n302,
         DP_mult_208_n301, DP_mult_208_n300, DP_mult_208_n299,
         DP_mult_208_n298, DP_mult_208_n296, DP_mult_208_n295,
         DP_mult_208_n294, DP_mult_208_n293, DP_mult_208_n292,
         DP_mult_208_n291, DP_mult_208_n290, DP_mult_208_n289,
         DP_mult_208_n288, DP_mult_208_n287, DP_mult_208_n286,
         DP_mult_208_n285, DP_mult_208_n284, DP_mult_208_n283,
         DP_mult_208_n282, DP_mult_208_n281, DP_mult_208_n280,
         DP_mult_208_n279, DP_mult_208_n278, DP_mult_208_n276,
         DP_mult_208_n275, DP_mult_208_n274, DP_mult_208_n273,
         DP_mult_208_n272, DP_mult_208_n271, DP_mult_208_n270,
         DP_mult_208_n269, DP_mult_208_n268, DP_mult_208_n267,
         DP_mult_208_n266, DP_mult_208_n265, DP_mult_208_n264,
         DP_mult_208_n263, DP_mult_208_n262, DP_mult_208_n261,
         DP_mult_208_n260, DP_mult_208_n259, DP_mult_208_n258,
         DP_mult_208_n257, DP_mult_208_n256, DP_mult_208_n255,
         DP_mult_208_n254, DP_mult_208_n253, DP_mult_208_n252,
         DP_mult_208_n251, DP_mult_208_n250, DP_mult_208_n249,
         DP_mult_208_n248, DP_mult_208_n247, DP_mult_208_n246,
         DP_mult_208_n245, DP_mult_208_n244, DP_mult_208_n243,
         DP_mult_208_n242, DP_mult_208_n241, DP_mult_208_n240,
         DP_mult_208_n239, DP_mult_208_n238, DP_mult_208_n237,
         DP_mult_208_n236, DP_mult_208_n235, DP_mult_208_n234,
         DP_mult_208_n233, DP_mult_208_n232, DP_mult_208_n231,
         DP_mult_208_n230, DP_mult_208_n229, DP_mult_208_n228,
         DP_mult_208_n227, DP_mult_208_n226, DP_mult_208_n225,
         DP_mult_208_n224, DP_mult_208_n223, DP_mult_208_n222,
         DP_mult_208_n221, DP_mult_208_n220, DP_mult_208_n219,
         DP_mult_208_n218, DP_mult_208_n217, DP_mult_208_n216,
         DP_mult_208_n215, DP_mult_208_n214, DP_mult_208_n213,
         DP_mult_208_n212, DP_mult_208_n211, DP_mult_208_n210,
         DP_mult_208_n209, DP_mult_208_n208, DP_mult_208_n207,
         DP_mult_208_n206, DP_mult_208_n205, DP_mult_208_n204,
         DP_mult_208_n203, DP_mult_208_n202, DP_mult_208_n201,
         DP_mult_208_n200, DP_mult_208_n199, DP_mult_208_n198,
         DP_mult_208_n197, DP_mult_208_n196, DP_mult_208_n195,
         DP_mult_208_n194, DP_mult_208_n193, DP_mult_208_n192,
         DP_mult_208_n191, DP_mult_208_n190, DP_mult_208_n189,
         DP_mult_208_n188, DP_mult_208_n187, DP_mult_208_n186,
         DP_mult_208_n185, DP_mult_208_n184, DP_mult_208_n183,
         DP_mult_208_n182, DP_mult_208_n181, DP_mult_208_n180,
         DP_mult_208_n179, DP_mult_208_n178, DP_mult_208_n177,
         DP_mult_208_n176, DP_mult_208_n175, DP_mult_208_n174,
         DP_mult_208_n173, DP_mult_208_n172, DP_mult_208_n171,
         DP_mult_208_n170, DP_mult_208_n169, DP_mult_208_n168,
         DP_mult_208_n167, DP_mult_208_n166, DP_mult_208_n165,
         DP_mult_208_n164, DP_mult_208_n163, DP_mult_208_n162,
         DP_mult_208_n161, DP_mult_208_n160, DP_mult_208_n159,
         DP_mult_208_n158, DP_mult_208_n157, DP_mult_208_n156,
         DP_mult_208_n155, DP_mult_208_n154, DP_mult_208_n153,
         DP_mult_208_n152, DP_mult_208_n151, DP_mult_208_n150,
         DP_mult_208_n149, DP_mult_208_n148, DP_mult_208_n147,
         DP_mult_208_n146, DP_mult_208_n145, DP_mult_208_n144,
         DP_mult_208_n143, DP_mult_208_n142, DP_mult_208_n141,
         DP_mult_208_n140, DP_mult_208_n139, DP_mult_208_n138,
         DP_mult_208_n137, DP_mult_208_n136, DP_mult_208_n135,
         DP_mult_208_n134, DP_mult_208_n133, DP_mult_208_n132,
         DP_mult_208_n131, DP_mult_208_n130, DP_mult_208_n129,
         DP_mult_208_n128, DP_mult_208_n127, DP_mult_208_n126,
         DP_mult_208_n125, DP_mult_208_n124, DP_mult_208_n123,
         DP_mult_208_n122, DP_mult_208_n121, DP_mult_208_n120,
         DP_sub_208_B_not_1_, DP_sub_208_B_not_2_, DP_sub_208_B_not_3_,
         DP_sub_208_B_not_4_, DP_sub_208_B_not_5_, DP_sub_208_B_not_6_,
         DP_sub_208_B_not_7_, DP_sub_208_B_not_8_, DP_sub_208_B_not_9_,
         DP_sub_208_B_not_10_, DP_sub_208_B_not_11_, DP_sub_208_B_not_12_,
         DP_sub_208_B_not_13_, DP_sub_208_B_not_14_, DP_sub_208_B_not_15_,
         DP_sub_208_B_not_16_, DP_sub_208_B_not_17_, DP_sub_208_B_not_18_,
         DP_sub_208_B_not_19_, DP_sub_208_B_not_20_, DP_sub_208_B_not_21_,
         DP_sub_208_B_not_22_, DP_sub_208_B_not_23_, DP_sub_208_carry_1_,
         DP_sub_208_carry_2_, DP_sub_208_carry_3_, DP_sub_208_carry_4_,
         DP_sub_208_carry_5_, DP_sub_208_carry_6_, DP_sub_208_carry_7_,
         DP_sub_208_carry_8_, DP_sub_208_carry_9_, DP_sub_208_carry_10_,
         DP_sub_208_carry_11_, DP_sub_208_carry_12_, DP_sub_208_carry_13_,
         DP_sub_208_carry_14_, DP_sub_208_carry_15_, DP_sub_208_carry_16_,
         DP_sub_208_carry_17_, DP_sub_208_carry_18_, DP_sub_208_carry_19_,
         DP_sub_208_carry_20_, DP_sub_208_carry_21_, DP_sub_208_carry_22_,
         DP_sub_208_carry_23_, DP_mult_209_n626, DP_mult_209_n625,
         DP_mult_209_n624, DP_mult_209_n623, DP_mult_209_n622,
         DP_mult_209_n621, DP_mult_209_n620, DP_mult_209_n619,
         DP_mult_209_n618, DP_mult_209_n617, DP_mult_209_n616,
         DP_mult_209_n615, DP_mult_209_n614, DP_mult_209_n613,
         DP_mult_209_n612, DP_mult_209_n611, DP_mult_209_n610,
         DP_mult_209_n609, DP_mult_209_n608, DP_mult_209_n607,
         DP_mult_209_n606, DP_mult_209_n605, DP_mult_209_n604,
         DP_mult_209_n603, DP_mult_209_n602, DP_mult_209_n601,
         DP_mult_209_n600, DP_mult_209_n599, DP_mult_209_n598,
         DP_mult_209_n597, DP_mult_209_n596, DP_mult_209_n595,
         DP_mult_209_n594, DP_mult_209_n593, DP_mult_209_n592,
         DP_mult_209_n591, DP_mult_209_n590, DP_mult_209_n589,
         DP_mult_209_n588, DP_mult_209_n587, DP_mult_209_n586,
         DP_mult_209_n585, DP_mult_209_n584, DP_mult_209_n583,
         DP_mult_209_n582, DP_mult_209_n581, DP_mult_209_n580,
         DP_mult_209_n579, DP_mult_209_n578, DP_mult_209_n577,
         DP_mult_209_n576, DP_mult_209_n575, DP_mult_209_n574,
         DP_mult_209_n573, DP_mult_209_n572, DP_mult_209_n571,
         DP_mult_209_n570, DP_mult_209_n569, DP_mult_209_n568,
         DP_mult_209_n567, DP_mult_209_n566, DP_mult_209_n565,
         DP_mult_209_n564, DP_mult_209_n563, DP_mult_209_n562,
         DP_mult_209_n561, DP_mult_209_n560, DP_mult_209_n559,
         DP_mult_209_n558, DP_mult_209_n557, DP_mult_209_n556,
         DP_mult_209_n555, DP_mult_209_n554, DP_mult_209_n553,
         DP_mult_209_n552, DP_mult_209_n551, DP_mult_209_n550,
         DP_mult_209_n549, DP_mult_209_n548, DP_mult_209_n547,
         DP_mult_209_n546, DP_mult_209_n545, DP_mult_209_n544,
         DP_mult_209_n543, DP_mult_209_n542, DP_mult_209_n541,
         DP_mult_209_n540, DP_mult_209_n539, DP_mult_209_n538,
         DP_mult_209_n537, DP_mult_209_n536, DP_mult_209_n535,
         DP_mult_209_n534, DP_mult_209_n533, DP_mult_209_n532,
         DP_mult_209_n531, DP_mult_209_n530, DP_mult_209_n529,
         DP_mult_209_n528, DP_mult_209_n527, DP_mult_209_n526,
         DP_mult_209_n525, DP_mult_209_n524, DP_mult_209_n523,
         DP_mult_209_n522, DP_mult_209_n521, DP_mult_209_n520,
         DP_mult_209_n519, DP_mult_209_n518, DP_mult_209_n517,
         DP_mult_209_n516, DP_mult_209_n515, DP_mult_209_n514,
         DP_mult_209_n513, DP_mult_209_n329, DP_mult_209_n328,
         DP_mult_209_n327, DP_mult_209_n326, DP_mult_209_n325,
         DP_mult_209_n324, DP_mult_209_n323, DP_mult_209_n322,
         DP_mult_209_n321, DP_mult_209_n320, DP_mult_209_n319,
         DP_mult_209_n318, DP_mult_209_n317, DP_mult_209_n316,
         DP_mult_209_n315, DP_mult_209_n314, DP_mult_209_n313,
         DP_mult_209_n312, DP_mult_209_n311, DP_mult_209_n310,
         DP_mult_209_n309, DP_mult_209_n308, DP_mult_209_n307,
         DP_mult_209_n306, DP_mult_209_n305, DP_mult_209_n304,
         DP_mult_209_n303, DP_mult_209_n302, DP_mult_209_n301,
         DP_mult_209_n300, DP_mult_209_n299, DP_mult_209_n298,
         DP_mult_209_n296, DP_mult_209_n295, DP_mult_209_n294,
         DP_mult_209_n293, DP_mult_209_n292, DP_mult_209_n291,
         DP_mult_209_n290, DP_mult_209_n289, DP_mult_209_n288,
         DP_mult_209_n287, DP_mult_209_n286, DP_mult_209_n285,
         DP_mult_209_n284, DP_mult_209_n283, DP_mult_209_n282,
         DP_mult_209_n281, DP_mult_209_n280, DP_mult_209_n279,
         DP_mult_209_n278, DP_mult_209_n276, DP_mult_209_n275,
         DP_mult_209_n274, DP_mult_209_n273, DP_mult_209_n272,
         DP_mult_209_n271, DP_mult_209_n270, DP_mult_209_n269,
         DP_mult_209_n268, DP_mult_209_n267, DP_mult_209_n266,
         DP_mult_209_n265, DP_mult_209_n264, DP_mult_209_n263,
         DP_mult_209_n262, DP_mult_209_n261, DP_mult_209_n260,
         DP_mult_209_n259, DP_mult_209_n258, DP_mult_209_n257,
         DP_mult_209_n256, DP_mult_209_n255, DP_mult_209_n254,
         DP_mult_209_n253, DP_mult_209_n252, DP_mult_209_n251,
         DP_mult_209_n250, DP_mult_209_n249, DP_mult_209_n248,
         DP_mult_209_n247, DP_mult_209_n246, DP_mult_209_n245,
         DP_mult_209_n244, DP_mult_209_n243, DP_mult_209_n242,
         DP_mult_209_n241, DP_mult_209_n240, DP_mult_209_n239,
         DP_mult_209_n238, DP_mult_209_n237, DP_mult_209_n236,
         DP_mult_209_n235, DP_mult_209_n234, DP_mult_209_n233,
         DP_mult_209_n232, DP_mult_209_n231, DP_mult_209_n230,
         DP_mult_209_n229, DP_mult_209_n228, DP_mult_209_n227,
         DP_mult_209_n226, DP_mult_209_n225, DP_mult_209_n224,
         DP_mult_209_n223, DP_mult_209_n222, DP_mult_209_n221,
         DP_mult_209_n220, DP_mult_209_n219, DP_mult_209_n218,
         DP_mult_209_n217, DP_mult_209_n216, DP_mult_209_n215,
         DP_mult_209_n214, DP_mult_209_n213, DP_mult_209_n212,
         DP_mult_209_n211, DP_mult_209_n210, DP_mult_209_n209,
         DP_mult_209_n208, DP_mult_209_n207, DP_mult_209_n206,
         DP_mult_209_n205, DP_mult_209_n204, DP_mult_209_n203,
         DP_mult_209_n202, DP_mult_209_n201, DP_mult_209_n200,
         DP_mult_209_n199, DP_mult_209_n198, DP_mult_209_n197,
         DP_mult_209_n196, DP_mult_209_n195, DP_mult_209_n194,
         DP_mult_209_n193, DP_mult_209_n192, DP_mult_209_n191,
         DP_mult_209_n190, DP_mult_209_n189, DP_mult_209_n188,
         DP_mult_209_n187, DP_mult_209_n186, DP_mult_209_n185,
         DP_mult_209_n184, DP_mult_209_n183, DP_mult_209_n182,
         DP_mult_209_n181, DP_mult_209_n180, DP_mult_209_n179,
         DP_mult_209_n178, DP_mult_209_n177, DP_mult_209_n176,
         DP_mult_209_n175, DP_mult_209_n174, DP_mult_209_n173,
         DP_mult_209_n172, DP_mult_209_n171, DP_mult_209_n170,
         DP_mult_209_n169, DP_mult_209_n168, DP_mult_209_n167,
         DP_mult_209_n166, DP_mult_209_n165, DP_mult_209_n164,
         DP_mult_209_n163, DP_mult_209_n162, DP_mult_209_n161,
         DP_mult_209_n160, DP_mult_209_n159, DP_mult_209_n158,
         DP_mult_209_n157, DP_mult_209_n156, DP_mult_209_n155,
         DP_mult_209_n154, DP_mult_209_n153, DP_mult_209_n152,
         DP_mult_209_n151, DP_mult_209_n150, DP_mult_209_n149,
         DP_mult_209_n148, DP_mult_209_n147, DP_mult_209_n146,
         DP_mult_209_n145, DP_mult_209_n144, DP_mult_209_n143,
         DP_mult_209_n142, DP_mult_209_n141, DP_mult_209_n140,
         DP_mult_209_n139, DP_mult_209_n138, DP_mult_209_n137,
         DP_mult_209_n136, DP_mult_209_n135, DP_mult_209_n134,
         DP_mult_209_n133, DP_mult_209_n132, DP_mult_209_n131,
         DP_mult_209_n130, DP_mult_209_n129, DP_mult_209_n128,
         DP_mult_209_n127, DP_mult_209_n126, DP_mult_209_n125,
         DP_mult_209_n124, DP_mult_209_n123, DP_mult_209_n122,
         DP_mult_209_n121, DP_mult_209_n120, DP_sub_209_B_not_1_,
         DP_sub_209_B_not_2_, DP_sub_209_B_not_3_, DP_sub_209_B_not_4_,
         DP_sub_209_B_not_5_, DP_sub_209_B_not_6_, DP_sub_209_B_not_7_,
         DP_sub_209_B_not_8_, DP_sub_209_B_not_9_, DP_sub_209_B_not_10_,
         DP_sub_209_B_not_11_, DP_sub_209_B_not_12_, DP_sub_209_B_not_13_,
         DP_sub_209_B_not_14_, DP_sub_209_B_not_15_, DP_sub_209_B_not_16_,
         DP_sub_209_B_not_17_, DP_sub_209_B_not_18_, DP_sub_209_B_not_19_,
         DP_sub_209_B_not_20_, DP_sub_209_B_not_21_, DP_sub_209_B_not_22_,
         DP_sub_209_B_not_23_, DP_sub_209_carry_1_, DP_sub_209_carry_2_,
         DP_sub_209_carry_3_, DP_sub_209_carry_4_, DP_sub_209_carry_5_,
         DP_sub_209_carry_6_, DP_sub_209_carry_7_, DP_sub_209_carry_8_,
         DP_sub_209_carry_9_, DP_sub_209_carry_10_, DP_sub_209_carry_11_,
         DP_sub_209_carry_12_, DP_sub_209_carry_13_, DP_sub_209_carry_14_,
         DP_sub_209_carry_15_, DP_sub_209_carry_16_, DP_sub_209_carry_17_,
         DP_sub_209_carry_18_, DP_sub_209_carry_19_, DP_sub_209_carry_20_,
         DP_sub_209_carry_21_, DP_sub_209_carry_22_, DP_sub_209_carry_23_,
         DP_mult_210_n626, DP_mult_210_n625, DP_mult_210_n624,
         DP_mult_210_n623, DP_mult_210_n622, DP_mult_210_n621,
         DP_mult_210_n620, DP_mult_210_n619, DP_mult_210_n618,
         DP_mult_210_n617, DP_mult_210_n616, DP_mult_210_n615,
         DP_mult_210_n614, DP_mult_210_n613, DP_mult_210_n612,
         DP_mult_210_n611, DP_mult_210_n610, DP_mult_210_n609,
         DP_mult_210_n608, DP_mult_210_n607, DP_mult_210_n606,
         DP_mult_210_n605, DP_mult_210_n604, DP_mult_210_n603,
         DP_mult_210_n602, DP_mult_210_n601, DP_mult_210_n600,
         DP_mult_210_n599, DP_mult_210_n598, DP_mult_210_n597,
         DP_mult_210_n596, DP_mult_210_n595, DP_mult_210_n594,
         DP_mult_210_n593, DP_mult_210_n592, DP_mult_210_n591,
         DP_mult_210_n590, DP_mult_210_n589, DP_mult_210_n588,
         DP_mult_210_n587, DP_mult_210_n586, DP_mult_210_n585,
         DP_mult_210_n584, DP_mult_210_n583, DP_mult_210_n582,
         DP_mult_210_n581, DP_mult_210_n580, DP_mult_210_n579,
         DP_mult_210_n578, DP_mult_210_n577, DP_mult_210_n576,
         DP_mult_210_n575, DP_mult_210_n574, DP_mult_210_n573,
         DP_mult_210_n572, DP_mult_210_n571, DP_mult_210_n570,
         DP_mult_210_n569, DP_mult_210_n568, DP_mult_210_n567,
         DP_mult_210_n566, DP_mult_210_n565, DP_mult_210_n564,
         DP_mult_210_n563, DP_mult_210_n562, DP_mult_210_n561,
         DP_mult_210_n560, DP_mult_210_n559, DP_mult_210_n558,
         DP_mult_210_n557, DP_mult_210_n556, DP_mult_210_n555,
         DP_mult_210_n554, DP_mult_210_n553, DP_mult_210_n552,
         DP_mult_210_n551, DP_mult_210_n550, DP_mult_210_n549,
         DP_mult_210_n548, DP_mult_210_n547, DP_mult_210_n546,
         DP_mult_210_n545, DP_mult_210_n544, DP_mult_210_n543,
         DP_mult_210_n542, DP_mult_210_n541, DP_mult_210_n540,
         DP_mult_210_n539, DP_mult_210_n538, DP_mult_210_n537,
         DP_mult_210_n536, DP_mult_210_n535, DP_mult_210_n534,
         DP_mult_210_n533, DP_mult_210_n532, DP_mult_210_n531,
         DP_mult_210_n530, DP_mult_210_n529, DP_mult_210_n528,
         DP_mult_210_n527, DP_mult_210_n526, DP_mult_210_n525,
         DP_mult_210_n524, DP_mult_210_n523, DP_mult_210_n522,
         DP_mult_210_n521, DP_mult_210_n520, DP_mult_210_n519,
         DP_mult_210_n518, DP_mult_210_n517, DP_mult_210_n516,
         DP_mult_210_n515, DP_mult_210_n514, DP_mult_210_n513,
         DP_mult_210_n329, DP_mult_210_n328, DP_mult_210_n327,
         DP_mult_210_n326, DP_mult_210_n325, DP_mult_210_n324,
         DP_mult_210_n323, DP_mult_210_n322, DP_mult_210_n321,
         DP_mult_210_n320, DP_mult_210_n319, DP_mult_210_n318,
         DP_mult_210_n317, DP_mult_210_n316, DP_mult_210_n315,
         DP_mult_210_n314, DP_mult_210_n313, DP_mult_210_n312,
         DP_mult_210_n311, DP_mult_210_n310, DP_mult_210_n309,
         DP_mult_210_n308, DP_mult_210_n307, DP_mult_210_n306,
         DP_mult_210_n305, DP_mult_210_n304, DP_mult_210_n303,
         DP_mult_210_n302, DP_mult_210_n301, DP_mult_210_n300,
         DP_mult_210_n299, DP_mult_210_n298, DP_mult_210_n296,
         DP_mult_210_n295, DP_mult_210_n294, DP_mult_210_n293,
         DP_mult_210_n292, DP_mult_210_n291, DP_mult_210_n290,
         DP_mult_210_n289, DP_mult_210_n288, DP_mult_210_n287,
         DP_mult_210_n286, DP_mult_210_n285, DP_mult_210_n284,
         DP_mult_210_n283, DP_mult_210_n282, DP_mult_210_n281,
         DP_mult_210_n280, DP_mult_210_n279, DP_mult_210_n278,
         DP_mult_210_n276, DP_mult_210_n275, DP_mult_210_n274,
         DP_mult_210_n273, DP_mult_210_n272, DP_mult_210_n271,
         DP_mult_210_n270, DP_mult_210_n269, DP_mult_210_n268,
         DP_mult_210_n267, DP_mult_210_n266, DP_mult_210_n265,
         DP_mult_210_n264, DP_mult_210_n263, DP_mult_210_n262,
         DP_mult_210_n261, DP_mult_210_n260, DP_mult_210_n259,
         DP_mult_210_n258, DP_mult_210_n257, DP_mult_210_n256,
         DP_mult_210_n255, DP_mult_210_n254, DP_mult_210_n253,
         DP_mult_210_n252, DP_mult_210_n251, DP_mult_210_n250,
         DP_mult_210_n249, DP_mult_210_n248, DP_mult_210_n247,
         DP_mult_210_n246, DP_mult_210_n245, DP_mult_210_n244,
         DP_mult_210_n243, DP_mult_210_n242, DP_mult_210_n241,
         DP_mult_210_n240, DP_mult_210_n239, DP_mult_210_n238,
         DP_mult_210_n237, DP_mult_210_n236, DP_mult_210_n235,
         DP_mult_210_n234, DP_mult_210_n233, DP_mult_210_n232,
         DP_mult_210_n231, DP_mult_210_n230, DP_mult_210_n229,
         DP_mult_210_n228, DP_mult_210_n227, DP_mult_210_n226,
         DP_mult_210_n225, DP_mult_210_n224, DP_mult_210_n223,
         DP_mult_210_n222, DP_mult_210_n221, DP_mult_210_n220,
         DP_mult_210_n219, DP_mult_210_n218, DP_mult_210_n217,
         DP_mult_210_n216, DP_mult_210_n215, DP_mult_210_n214,
         DP_mult_210_n213, DP_mult_210_n212, DP_mult_210_n211,
         DP_mult_210_n210, DP_mult_210_n209, DP_mult_210_n208,
         DP_mult_210_n207, DP_mult_210_n206, DP_mult_210_n205,
         DP_mult_210_n204, DP_mult_210_n203, DP_mult_210_n202,
         DP_mult_210_n201, DP_mult_210_n200, DP_mult_210_n199,
         DP_mult_210_n198, DP_mult_210_n197, DP_mult_210_n196,
         DP_mult_210_n195, DP_mult_210_n194, DP_mult_210_n193,
         DP_mult_210_n192, DP_mult_210_n191, DP_mult_210_n190,
         DP_mult_210_n189, DP_mult_210_n188, DP_mult_210_n187,
         DP_mult_210_n186, DP_mult_210_n185, DP_mult_210_n184,
         DP_mult_210_n183, DP_mult_210_n182, DP_mult_210_n181,
         DP_mult_210_n180, DP_mult_210_n179, DP_mult_210_n178,
         DP_mult_210_n177, DP_mult_210_n176, DP_mult_210_n175,
         DP_mult_210_n174, DP_mult_210_n173, DP_mult_210_n172,
         DP_mult_210_n171, DP_mult_210_n170, DP_mult_210_n169,
         DP_mult_210_n168, DP_mult_210_n167, DP_mult_210_n166,
         DP_mult_210_n165, DP_mult_210_n164, DP_mult_210_n163,
         DP_mult_210_n162, DP_mult_210_n161, DP_mult_210_n160,
         DP_mult_210_n159, DP_mult_210_n158, DP_mult_210_n157,
         DP_mult_210_n156, DP_mult_210_n155, DP_mult_210_n154,
         DP_mult_210_n153, DP_mult_210_n152, DP_mult_210_n151,
         DP_mult_210_n150, DP_mult_210_n149, DP_mult_210_n148,
         DP_mult_210_n147, DP_mult_210_n146, DP_mult_210_n145,
         DP_mult_210_n144, DP_mult_210_n143, DP_mult_210_n142,
         DP_mult_210_n141, DP_mult_210_n140, DP_mult_210_n139,
         DP_mult_210_n138, DP_mult_210_n137, DP_mult_210_n136,
         DP_mult_210_n135, DP_mult_210_n134, DP_mult_210_n133,
         DP_mult_210_n132, DP_mult_210_n131, DP_mult_210_n130,
         DP_mult_210_n129, DP_mult_210_n128, DP_mult_210_n127,
         DP_mult_210_n126, DP_mult_210_n125, DP_mult_210_n124,
         DP_mult_210_n123, DP_mult_210_n122, DP_mult_210_n121,
         DP_mult_210_n120, DP_sub_210_B_not_1_, DP_sub_210_B_not_2_,
         DP_sub_210_B_not_3_, DP_sub_210_B_not_4_, DP_sub_210_B_not_5_,
         DP_sub_210_B_not_6_, DP_sub_210_B_not_7_, DP_sub_210_B_not_8_,
         DP_sub_210_B_not_9_, DP_sub_210_B_not_10_, DP_sub_210_B_not_11_,
         DP_sub_210_B_not_12_, DP_sub_210_B_not_13_, DP_sub_210_B_not_14_,
         DP_sub_210_B_not_15_, DP_sub_210_B_not_16_, DP_sub_210_B_not_17_,
         DP_sub_210_B_not_18_, DP_sub_210_B_not_19_, DP_sub_210_B_not_20_,
         DP_sub_210_B_not_21_, DP_sub_210_B_not_22_, DP_sub_210_B_not_23_,
         DP_sub_210_carry_1_, DP_sub_210_carry_2_, DP_sub_210_carry_3_,
         DP_sub_210_carry_4_, DP_sub_210_carry_5_, DP_sub_210_carry_6_,
         DP_sub_210_carry_7_, DP_sub_210_carry_8_, DP_sub_210_carry_9_,
         DP_sub_210_carry_10_, DP_sub_210_carry_11_, DP_sub_210_carry_12_,
         DP_sub_210_carry_13_, DP_sub_210_carry_14_, DP_sub_210_carry_15_,
         DP_sub_210_carry_16_, DP_sub_210_carry_17_, DP_sub_210_carry_18_,
         DP_sub_210_carry_19_, DP_sub_210_carry_20_, DP_sub_210_carry_21_,
         DP_sub_210_carry_22_, DP_sub_210_carry_23_, DP_mult_211_n621,
         DP_mult_211_n620, DP_mult_211_n619, DP_mult_211_n618,
         DP_mult_211_n617, DP_mult_211_n616, DP_mult_211_n615,
         DP_mult_211_n614, DP_mult_211_n613, DP_mult_211_n612,
         DP_mult_211_n611, DP_mult_211_n610, DP_mult_211_n609,
         DP_mult_211_n608, DP_mult_211_n607, DP_mult_211_n606,
         DP_mult_211_n605, DP_mult_211_n604, DP_mult_211_n603,
         DP_mult_211_n602, DP_mult_211_n601, DP_mult_211_n600,
         DP_mult_211_n599, DP_mult_211_n598, DP_mult_211_n597,
         DP_mult_211_n596, DP_mult_211_n595, DP_mult_211_n594,
         DP_mult_211_n593, DP_mult_211_n592, DP_mult_211_n591,
         DP_mult_211_n590, DP_mult_211_n589, DP_mult_211_n588,
         DP_mult_211_n587, DP_mult_211_n586, DP_mult_211_n585,
         DP_mult_211_n584, DP_mult_211_n583, DP_mult_211_n582,
         DP_mult_211_n581, DP_mult_211_n580, DP_mult_211_n579,
         DP_mult_211_n578, DP_mult_211_n577, DP_mult_211_n576,
         DP_mult_211_n575, DP_mult_211_n574, DP_mult_211_n573,
         DP_mult_211_n572, DP_mult_211_n571, DP_mult_211_n570,
         DP_mult_211_n569, DP_mult_211_n568, DP_mult_211_n567,
         DP_mult_211_n566, DP_mult_211_n565, DP_mult_211_n564,
         DP_mult_211_n563, DP_mult_211_n562, DP_mult_211_n561,
         DP_mult_211_n560, DP_mult_211_n559, DP_mult_211_n558,
         DP_mult_211_n557, DP_mult_211_n556, DP_mult_211_n555,
         DP_mult_211_n554, DP_mult_211_n553, DP_mult_211_n552,
         DP_mult_211_n551, DP_mult_211_n550, DP_mult_211_n549,
         DP_mult_211_n548, DP_mult_211_n547, DP_mult_211_n546,
         DP_mult_211_n545, DP_mult_211_n544, DP_mult_211_n543,
         DP_mult_211_n542, DP_mult_211_n541, DP_mult_211_n540,
         DP_mult_211_n539, DP_mult_211_n538, DP_mult_211_n537,
         DP_mult_211_n536, DP_mult_211_n535, DP_mult_211_n534,
         DP_mult_211_n533, DP_mult_211_n532, DP_mult_211_n531,
         DP_mult_211_n530, DP_mult_211_n529, DP_mult_211_n528,
         DP_mult_211_n527, DP_mult_211_n526, DP_mult_211_n525,
         DP_mult_211_n524, DP_mult_211_n523, DP_mult_211_n522,
         DP_mult_211_n521, DP_mult_211_n520, DP_mult_211_n519,
         DP_mult_211_n518, DP_mult_211_n517, DP_mult_211_n516,
         DP_mult_211_n515, DP_mult_211_n514, DP_mult_211_n513,
         DP_mult_211_n329, DP_mult_211_n328, DP_mult_211_n327,
         DP_mult_211_n326, DP_mult_211_n325, DP_mult_211_n324,
         DP_mult_211_n323, DP_mult_211_n322, DP_mult_211_n321,
         DP_mult_211_n320, DP_mult_211_n319, DP_mult_211_n318,
         DP_mult_211_n317, DP_mult_211_n316, DP_mult_211_n315,
         DP_mult_211_n314, DP_mult_211_n313, DP_mult_211_n312,
         DP_mult_211_n311, DP_mult_211_n310, DP_mult_211_n309,
         DP_mult_211_n308, DP_mult_211_n307, DP_mult_211_n306,
         DP_mult_211_n305, DP_mult_211_n304, DP_mult_211_n303,
         DP_mult_211_n302, DP_mult_211_n301, DP_mult_211_n300,
         DP_mult_211_n299, DP_mult_211_n298, DP_mult_211_n296,
         DP_mult_211_n295, DP_mult_211_n294, DP_mult_211_n293,
         DP_mult_211_n292, DP_mult_211_n291, DP_mult_211_n290,
         DP_mult_211_n289, DP_mult_211_n288, DP_mult_211_n287,
         DP_mult_211_n286, DP_mult_211_n285, DP_mult_211_n284,
         DP_mult_211_n283, DP_mult_211_n282, DP_mult_211_n281,
         DP_mult_211_n280, DP_mult_211_n279, DP_mult_211_n278,
         DP_mult_211_n276, DP_mult_211_n275, DP_mult_211_n274,
         DP_mult_211_n273, DP_mult_211_n272, DP_mult_211_n271,
         DP_mult_211_n270, DP_mult_211_n269, DP_mult_211_n268,
         DP_mult_211_n267, DP_mult_211_n266, DP_mult_211_n265,
         DP_mult_211_n264, DP_mult_211_n263, DP_mult_211_n262,
         DP_mult_211_n261, DP_mult_211_n260, DP_mult_211_n259,
         DP_mult_211_n258, DP_mult_211_n257, DP_mult_211_n256,
         DP_mult_211_n255, DP_mult_211_n254, DP_mult_211_n253,
         DP_mult_211_n252, DP_mult_211_n251, DP_mult_211_n250,
         DP_mult_211_n249, DP_mult_211_n248, DP_mult_211_n247,
         DP_mult_211_n246, DP_mult_211_n245, DP_mult_211_n244,
         DP_mult_211_n243, DP_mult_211_n242, DP_mult_211_n241,
         DP_mult_211_n240, DP_mult_211_n239, DP_mult_211_n238,
         DP_mult_211_n237, DP_mult_211_n236, DP_mult_211_n235,
         DP_mult_211_n234, DP_mult_211_n233, DP_mult_211_n232,
         DP_mult_211_n231, DP_mult_211_n230, DP_mult_211_n229,
         DP_mult_211_n228, DP_mult_211_n227, DP_mult_211_n226,
         DP_mult_211_n225, DP_mult_211_n224, DP_mult_211_n223,
         DP_mult_211_n222, DP_mult_211_n221, DP_mult_211_n220,
         DP_mult_211_n219, DP_mult_211_n218, DP_mult_211_n217,
         DP_mult_211_n216, DP_mult_211_n215, DP_mult_211_n214,
         DP_mult_211_n213, DP_mult_211_n212, DP_mult_211_n211,
         DP_mult_211_n210, DP_mult_211_n209, DP_mult_211_n208,
         DP_mult_211_n207, DP_mult_211_n206, DP_mult_211_n205,
         DP_mult_211_n204, DP_mult_211_n203, DP_mult_211_n202,
         DP_mult_211_n201, DP_mult_211_n200, DP_mult_211_n199,
         DP_mult_211_n198, DP_mult_211_n197, DP_mult_211_n196,
         DP_mult_211_n195, DP_mult_211_n194, DP_mult_211_n193,
         DP_mult_211_n192, DP_mult_211_n191, DP_mult_211_n190,
         DP_mult_211_n189, DP_mult_211_n188, DP_mult_211_n187,
         DP_mult_211_n186, DP_mult_211_n185, DP_mult_211_n184,
         DP_mult_211_n183, DP_mult_211_n182, DP_mult_211_n181,
         DP_mult_211_n180, DP_mult_211_n179, DP_mult_211_n178,
         DP_mult_211_n177, DP_mult_211_n176, DP_mult_211_n175,
         DP_mult_211_n174, DP_mult_211_n173, DP_mult_211_n172,
         DP_mult_211_n171, DP_mult_211_n170, DP_mult_211_n169,
         DP_mult_211_n168, DP_mult_211_n167, DP_mult_211_n166,
         DP_mult_211_n165, DP_mult_211_n164, DP_mult_211_n163,
         DP_mult_211_n162, DP_mult_211_n161, DP_mult_211_n160,
         DP_mult_211_n159, DP_mult_211_n158, DP_mult_211_n157,
         DP_mult_211_n156, DP_mult_211_n155, DP_mult_211_n154,
         DP_mult_211_n153, DP_mult_211_n152, DP_mult_211_n151,
         DP_mult_211_n150, DP_mult_211_n149, DP_mult_211_n148,
         DP_mult_211_n147, DP_mult_211_n146, DP_mult_211_n145,
         DP_mult_211_n144, DP_mult_211_n143, DP_mult_211_n142,
         DP_mult_211_n141, DP_mult_211_n140, DP_mult_211_n139,
         DP_mult_211_n138, DP_mult_211_n137, DP_mult_211_n136,
         DP_mult_211_n135, DP_mult_211_n134, DP_mult_211_n133,
         DP_mult_211_n132, DP_mult_211_n131, DP_mult_211_n130,
         DP_mult_211_n129, DP_mult_211_n128, DP_mult_211_n127,
         DP_mult_211_n126, DP_mult_211_n125, DP_mult_211_n124,
         DP_mult_211_n123, DP_mult_211_n122, DP_mult_211_n121,
         DP_mult_211_n120, DP_sub_211_B_not_1_, DP_sub_211_B_not_2_,
         DP_sub_211_B_not_3_, DP_sub_211_B_not_4_, DP_sub_211_B_not_5_,
         DP_sub_211_B_not_6_, DP_sub_211_B_not_7_, DP_sub_211_B_not_8_,
         DP_sub_211_B_not_9_, DP_sub_211_B_not_10_, DP_sub_211_B_not_11_,
         DP_sub_211_B_not_12_, DP_sub_211_B_not_13_, DP_sub_211_B_not_14_,
         DP_sub_211_B_not_15_, DP_sub_211_B_not_16_, DP_sub_211_B_not_17_,
         DP_sub_211_B_not_18_, DP_sub_211_B_not_19_, DP_sub_211_B_not_20_,
         DP_sub_211_B_not_21_, DP_sub_211_B_not_22_, DP_sub_211_B_not_23_,
         DP_sub_211_carry_1_, DP_sub_211_carry_2_, DP_sub_211_carry_3_,
         DP_sub_211_carry_4_, DP_sub_211_carry_5_, DP_sub_211_carry_6_,
         DP_sub_211_carry_7_, DP_sub_211_carry_8_, DP_sub_211_carry_9_,
         DP_sub_211_carry_10_, DP_sub_211_carry_11_, DP_sub_211_carry_12_,
         DP_sub_211_carry_13_, DP_sub_211_carry_14_, DP_sub_211_carry_15_,
         DP_sub_211_carry_16_, DP_sub_211_carry_17_, DP_sub_211_carry_18_,
         DP_sub_211_carry_19_, DP_sub_211_carry_20_, DP_sub_211_carry_21_,
         DP_sub_211_carry_22_, DP_sub_211_carry_23_,
         DP_add_1_root_sub_0_root_sub_227_carry_1_,
         DP_add_1_root_sub_0_root_sub_227_carry_2_,
         DP_add_1_root_sub_0_root_sub_227_carry_3_,
         DP_add_1_root_sub_0_root_sub_227_carry_4_,
         DP_add_1_root_sub_0_root_sub_227_carry_5_,
         DP_add_1_root_sub_0_root_sub_227_carry_6_,
         DP_add_1_root_sub_0_root_sub_227_carry_7_,
         DP_add_1_root_sub_0_root_sub_227_carry_8_,
         DP_add_1_root_sub_0_root_sub_227_carry_9_,
         DP_add_1_root_sub_0_root_sub_227_carry_10_,
         DP_add_1_root_sub_0_root_sub_227_carry_11_,
         DP_add_1_root_sub_0_root_sub_227_carry_12_,
         DP_add_1_root_sub_0_root_sub_227_carry_13_,
         DP_add_1_root_sub_0_root_sub_227_carry_14_,
         DP_add_1_root_sub_0_root_sub_227_carry_15_,
         DP_add_1_root_sub_0_root_sub_227_carry_16_,
         DP_add_1_root_sub_0_root_sub_227_carry_17_,
         DP_add_1_root_sub_0_root_sub_227_carry_18_,
         DP_add_1_root_sub_0_root_sub_227_carry_19_,
         DP_add_1_root_sub_0_root_sub_227_carry_20_,
         DP_add_1_root_sub_0_root_sub_227_carry_21_,
         DP_add_1_root_sub_0_root_sub_227_carry_22_,
         DP_add_1_root_sub_0_root_sub_227_carry_23_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_1_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_2_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_3_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_4_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_5_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_6_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_7_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_8_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_9_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_10_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_11_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_12_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_13_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_14_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_15_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_16_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_17_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_18_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_19_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_20_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_21_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_22_,
         DP_sub_0_root_sub_0_root_sub_227_B_not_23_,
         DP_sub_0_root_sub_0_root_sub_227_carry_1_,
         DP_sub_0_root_sub_0_root_sub_227_carry_2_,
         DP_sub_0_root_sub_0_root_sub_227_carry_3_,
         DP_sub_0_root_sub_0_root_sub_227_carry_4_,
         DP_sub_0_root_sub_0_root_sub_227_carry_5_,
         DP_sub_0_root_sub_0_root_sub_227_carry_6_,
         DP_sub_0_root_sub_0_root_sub_227_carry_7_,
         DP_sub_0_root_sub_0_root_sub_227_carry_8_,
         DP_sub_0_root_sub_0_root_sub_227_carry_9_,
         DP_sub_0_root_sub_0_root_sub_227_carry_10_,
         DP_sub_0_root_sub_0_root_sub_227_carry_11_,
         DP_sub_0_root_sub_0_root_sub_227_carry_12_,
         DP_sub_0_root_sub_0_root_sub_227_carry_13_,
         DP_sub_0_root_sub_0_root_sub_227_carry_14_,
         DP_sub_0_root_sub_0_root_sub_227_carry_15_,
         DP_sub_0_root_sub_0_root_sub_227_carry_16_,
         DP_sub_0_root_sub_0_root_sub_227_carry_17_,
         DP_sub_0_root_sub_0_root_sub_227_carry_18_,
         DP_sub_0_root_sub_0_root_sub_227_carry_19_,
         DP_sub_0_root_sub_0_root_sub_227_carry_20_,
         DP_sub_0_root_sub_0_root_sub_227_carry_21_,
         DP_sub_0_root_sub_0_root_sub_227_carry_22_,
         DP_sub_0_root_sub_0_root_sub_227_carry_23_, CU_n2, CU_nextState_0_,
         CU_presentState_0_, reg_delay_0_n6, reg_delay_0_n5, reg_delay_0_n4,
         reg_delay_0_n3, reg_delay_0_n2, reg_delay_0_n1, reg_delay_1_n12,
         reg_delay_1_n11, reg_delay_1_n10, reg_delay_1_n9, reg_delay_1_n8,
         reg_delay_1_n7;
  wire   [0:23] DP_coeff_pipe03;
  wire   [0:23] DP_coeff_pipe02;
  wire   [0:23] DP_coeff_pipe01;
  wire   [0:23] DP_coeff_ret1;
  wire   [1:23] DP_coeff_ret0;
  wire   [0:11] DP_y_out;
  wire   [0:23] DP_pipe13;
  wire   [0:23] DP_pipe0_coeff_pipe03;
  wire   [0:23] DP_pipe12;
  wire   [0:23] DP_pipe0_coeff_pipe02;
  wire   [0:23] DP_pipe11;
  wire   [0:23] DP_pipe0_coeff_pipe01;
  wire   [0:23] DP_pipe10;
  wire   [0:23] DP_pipe0_b0;
  wire   [0:23] DP_pipe03;
  wire   [0:23] DP_pipe02;
  wire   [0:23] DP_pipe01;
  wire   [0:23] DP_pipe00;
  wire   [0:23] DP_ret1;
  wire   [0:23] DP_sw1_coeff_ret1;
  wire   [0:23] DP_ret0;
  wire   [0:23] DP_sw0_coeff_ret0;
  wire   [0:23] DP_sw2;

  OAI22_X1 DP_U42 ( .A1(DP_y_23), .A2(DP_n13), .B1(DP_y_23), .B2(DP_n11), .ZN(
        DP_N146) );
  AND2_X1 DP_U41 ( .A1(DP_n12), .A2(DP_n11), .ZN(DP_n13) );
  NOR2_X1 DP_U40 ( .A1(DP_n9), .A2(DP_n8), .ZN(DP_n10) );
  NAND3_X1 DP_U39 ( .A1(DP_y_23), .A2(DP_y_11_), .A3(DP_y_23), .ZN(DP_n9) );
  BUF_X1 DP_U38 ( .A(rst_n), .Z(DP_n7) );
  BUF_X1 DP_U37 ( .A(rst_n), .Z(DP_n1) );
  BUF_X1 DP_U36 ( .A(rst_n), .Z(DP_n6) );
  BUF_X1 DP_U35 ( .A(rst_n), .Z(DP_n5) );
  BUF_X1 DP_U34 ( .A(rst_n), .Z(DP_n4) );
  BUF_X1 DP_U33 ( .A(rst_n), .Z(DP_n3) );
  BUF_X1 DP_U32 ( .A(rst_n), .Z(DP_n2) );
  INV_X1 DP_U31 ( .A(DP_y_0_), .ZN(DP_n66) );
  OAI21_X1 DP_U30 ( .B1(DP_N148), .B2(DP_n66), .A(DP_n55), .ZN(DP_y_out[0]) );
  INV_X1 DP_U29 ( .A(DP_y_10_), .ZN(DP_n65) );
  OAI21_X1 DP_U28 ( .B1(DP_N148), .B2(DP_n65), .A(DP_n55), .ZN(DP_y_out[10])
         );
  INV_X1 DP_U27 ( .A(DP_y_9_), .ZN(DP_n54) );
  OAI21_X1 DP_U26 ( .B1(DP_N148), .B2(DP_n54), .A(DP_n55), .ZN(DP_y_out[9]) );
  INV_X1 DP_U25 ( .A(DP_y_8_), .ZN(DP_n56) );
  OAI21_X1 DP_U24 ( .B1(DP_N148), .B2(DP_n56), .A(DP_n55), .ZN(DP_y_out[8]) );
  INV_X1 DP_U23 ( .A(DP_y_7_), .ZN(DP_n57) );
  OAI21_X1 DP_U22 ( .B1(DP_N148), .B2(DP_n57), .A(DP_n55), .ZN(DP_y_out[7]) );
  INV_X1 DP_U21 ( .A(DP_y_6_), .ZN(DP_n58) );
  OAI21_X1 DP_U20 ( .B1(DP_N148), .B2(DP_n58), .A(DP_n55), .ZN(DP_y_out[6]) );
  INV_X1 DP_U19 ( .A(DP_y_5_), .ZN(DP_n59) );
  OAI21_X1 DP_U18 ( .B1(DP_N148), .B2(DP_n59), .A(DP_n55), .ZN(DP_y_out[5]) );
  INV_X1 DP_U17 ( .A(DP_y_4_), .ZN(DP_n60) );
  OAI21_X1 DP_U16 ( .B1(DP_N148), .B2(DP_n60), .A(DP_n55), .ZN(DP_y_out[4]) );
  INV_X1 DP_U15 ( .A(DP_y_3_), .ZN(DP_n61) );
  OAI21_X1 DP_U14 ( .B1(DP_N148), .B2(DP_n61), .A(DP_n55), .ZN(DP_y_out[3]) );
  INV_X1 DP_U13 ( .A(DP_y_2_), .ZN(DP_n62) );
  OAI21_X1 DP_U12 ( .B1(DP_N148), .B2(DP_n62), .A(DP_n55), .ZN(DP_y_out[2]) );
  INV_X1 DP_U11 ( .A(DP_y_1_), .ZN(DP_n63) );
  OAI21_X1 DP_U10 ( .B1(DP_N148), .B2(DP_n63), .A(DP_n55), .ZN(DP_y_out[1]) );
  INV_X1 DP_U9 ( .A(DP_y_23), .ZN(DP_n11) );
  NOR2_X1 DP_U8 ( .A1(DP_y_23), .A2(DP_N148), .ZN(DP_n64) );
  NOR2_X1 DP_U7 ( .A1(DP_N146), .A2(DP_n64), .ZN(DP_y_out[11]) );
  NOR2_X1 DP_U6 ( .A1(DP_y_23), .A2(DP_y_11_), .ZN(DP_n12) );
  NAND2_X1 DP_U5 ( .A1(DP_y_23), .A2(DP_y_23), .ZN(DP_n8) );
  OAI22_X2 DP_U4 ( .A1(DP_n10), .A2(DP_n11), .B1(DP_y_23), .B2(DP_n11), .ZN(
        DP_N148) );
  INV_X1 DP_U3 ( .A(DP_N146), .ZN(DP_n55) );
  NAND2_X1 DP_reg_in_U28 ( .A1(dIn[11]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n12) );
  OAI21_X1 DP_reg_in_U27 ( .B1(DP_reg_in_n37), .B2(DP_reg_in_n24), .A(
        DP_reg_in_n12), .ZN(DP_reg_in_n36) );
  NAND2_X1 DP_reg_in_U26 ( .A1(dIn[10]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n11) );
  OAI21_X1 DP_reg_in_U25 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n23), .A(
        DP_reg_in_n11), .ZN(DP_reg_in_n35) );
  NAND2_X1 DP_reg_in_U24 ( .A1(dIn[9]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n10)
         );
  OAI21_X1 DP_reg_in_U23 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n22), .A(
        DP_reg_in_n10), .ZN(DP_reg_in_n34) );
  NAND2_X1 DP_reg_in_U22 ( .A1(dIn[8]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n9)
         );
  OAI21_X1 DP_reg_in_U21 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n21), .A(
        DP_reg_in_n9), .ZN(DP_reg_in_n33) );
  NAND2_X1 DP_reg_in_U20 ( .A1(dIn[7]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n8)
         );
  OAI21_X1 DP_reg_in_U19 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n20), .A(
        DP_reg_in_n8), .ZN(DP_reg_in_n32) );
  NAND2_X1 DP_reg_in_U18 ( .A1(dIn[6]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n7)
         );
  OAI21_X1 DP_reg_in_U17 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n19), .A(
        DP_reg_in_n7), .ZN(DP_reg_in_n31) );
  NAND2_X1 DP_reg_in_U16 ( .A1(dIn[5]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n6)
         );
  OAI21_X1 DP_reg_in_U15 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n18), .A(
        DP_reg_in_n6), .ZN(DP_reg_in_n30) );
  NAND2_X1 DP_reg_in_U14 ( .A1(dIn[4]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n5)
         );
  OAI21_X1 DP_reg_in_U13 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n17), .A(
        DP_reg_in_n5), .ZN(DP_reg_in_n29) );
  NAND2_X1 DP_reg_in_U12 ( .A1(dIn[3]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n4)
         );
  OAI21_X1 DP_reg_in_U11 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n16), .A(
        DP_reg_in_n4), .ZN(DP_reg_in_n28) );
  NAND2_X1 DP_reg_in_U10 ( .A1(dIn[2]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n3)
         );
  OAI21_X1 DP_reg_in_U9 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n15), .A(
        DP_reg_in_n3), .ZN(DP_reg_in_n27) );
  NAND2_X1 DP_reg_in_U8 ( .A1(dIn[1]), .A2(DP_reg_in_n37), .ZN(DP_reg_in_n2)
         );
  OAI21_X1 DP_reg_in_U7 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n14), .A(
        DP_reg_in_n2), .ZN(DP_reg_in_n26) );
  NAND2_X1 DP_reg_in_U6 ( .A1(DP_reg_in_n38), .A2(dIn[0]), .ZN(DP_reg_in_n1)
         );
  OAI21_X1 DP_reg_in_U5 ( .B1(DP_reg_in_n38), .B2(DP_reg_in_n13), .A(
        DP_reg_in_n1), .ZN(DP_reg_in_n25) );
  BUF_X1 DP_reg_in_U4 ( .A(vIn), .Z(DP_reg_in_n38) );
  BUF_X1 DP_reg_in_U3 ( .A(vIn), .Z(DP_reg_in_n37) );
  BUF_X1 DP_reg_in_U2 ( .A(DP_n7), .Z(DP_reg_in_n39) );
  DFFR_X1 DP_reg_in_Q_reg_0_ ( .D(DP_reg_in_n25), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_0_), .QN(DP_reg_in_n13) );
  DFFR_X1 DP_reg_in_Q_reg_1_ ( .D(DP_reg_in_n26), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_1_), .QN(DP_reg_in_n14) );
  DFFR_X1 DP_reg_in_Q_reg_2_ ( .D(DP_reg_in_n27), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_2_), .QN(DP_reg_in_n15) );
  DFFR_X1 DP_reg_in_Q_reg_3_ ( .D(DP_reg_in_n28), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_3_), .QN(DP_reg_in_n16) );
  DFFR_X1 DP_reg_in_Q_reg_4_ ( .D(DP_reg_in_n29), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_4_), .QN(DP_reg_in_n17) );
  DFFR_X1 DP_reg_in_Q_reg_5_ ( .D(DP_reg_in_n30), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_5_), .QN(DP_reg_in_n18) );
  DFFR_X1 DP_reg_in_Q_reg_6_ ( .D(DP_reg_in_n31), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_6_), .QN(DP_reg_in_n19) );
  DFFR_X1 DP_reg_in_Q_reg_7_ ( .D(DP_reg_in_n32), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_7_), .QN(DP_reg_in_n20) );
  DFFR_X1 DP_reg_in_Q_reg_8_ ( .D(DP_reg_in_n33), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_8_), .QN(DP_reg_in_n21) );
  DFFR_X1 DP_reg_in_Q_reg_9_ ( .D(DP_reg_in_n34), .CK(clk), .RN(DP_reg_in_n39), 
        .Q(DP_x_9_), .QN(DP_reg_in_n22) );
  DFFR_X1 DP_reg_in_Q_reg_10_ ( .D(DP_reg_in_n35), .CK(clk), .RN(DP_reg_in_n39), .Q(DP_x_10_), .QN(DP_reg_in_n23) );
  DFFR_X1 DP_reg_in_Q_reg_11_ ( .D(DP_reg_in_n36), .CK(clk), .RN(DP_reg_in_n39), .Q(DP_x_11_), .QN(DP_reg_in_n24) );
  NAND2_X1 DP_reg_a_i_1_U28 ( .A1(a[23]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n64) );
  OAI21_X1 DP_reg_a_i_1_U27 ( .B1(DP_reg_a_i_1_n37), .B2(DP_reg_a_i_1_n52), 
        .A(DP_reg_a_i_1_n64), .ZN(DP_reg_a_i_1_n40) );
  NAND2_X1 DP_reg_a_i_1_U26 ( .A1(a[22]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n65) );
  OAI21_X1 DP_reg_a_i_1_U25 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n53), 
        .A(DP_reg_a_i_1_n65), .ZN(DP_reg_a_i_1_n41) );
  NAND2_X1 DP_reg_a_i_1_U24 ( .A1(a[21]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n66) );
  OAI21_X1 DP_reg_a_i_1_U23 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n54), 
        .A(DP_reg_a_i_1_n66), .ZN(DP_reg_a_i_1_n42) );
  NAND2_X1 DP_reg_a_i_1_U22 ( .A1(a[20]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n67) );
  OAI21_X1 DP_reg_a_i_1_U21 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n55), 
        .A(DP_reg_a_i_1_n67), .ZN(DP_reg_a_i_1_n43) );
  NAND2_X1 DP_reg_a_i_1_U20 ( .A1(a[19]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n68) );
  OAI21_X1 DP_reg_a_i_1_U19 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n56), 
        .A(DP_reg_a_i_1_n68), .ZN(DP_reg_a_i_1_n44) );
  NAND2_X1 DP_reg_a_i_1_U18 ( .A1(a[18]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n69) );
  OAI21_X1 DP_reg_a_i_1_U17 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n57), 
        .A(DP_reg_a_i_1_n69), .ZN(DP_reg_a_i_1_n45) );
  NAND2_X1 DP_reg_a_i_1_U16 ( .A1(a[17]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n70) );
  OAI21_X1 DP_reg_a_i_1_U15 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n58), 
        .A(DP_reg_a_i_1_n70), .ZN(DP_reg_a_i_1_n46) );
  NAND2_X1 DP_reg_a_i_1_U14 ( .A1(a[16]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n71) );
  OAI21_X1 DP_reg_a_i_1_U13 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n59), 
        .A(DP_reg_a_i_1_n71), .ZN(DP_reg_a_i_1_n47) );
  NAND2_X1 DP_reg_a_i_1_U12 ( .A1(a[15]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n72) );
  OAI21_X1 DP_reg_a_i_1_U11 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n60), 
        .A(DP_reg_a_i_1_n72), .ZN(DP_reg_a_i_1_n48) );
  NAND2_X1 DP_reg_a_i_1_U10 ( .A1(a[14]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n73) );
  OAI21_X1 DP_reg_a_i_1_U9 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n61), .A(
        DP_reg_a_i_1_n73), .ZN(DP_reg_a_i_1_n49) );
  NAND2_X1 DP_reg_a_i_1_U8 ( .A1(a[13]), .A2(DP_reg_a_i_1_n37), .ZN(
        DP_reg_a_i_1_n74) );
  OAI21_X1 DP_reg_a_i_1_U7 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n62), .A(
        DP_reg_a_i_1_n74), .ZN(DP_reg_a_i_1_n50) );
  NAND2_X1 DP_reg_a_i_1_U6 ( .A1(DP_reg_a_i_1_n38), .A2(a[12]), .ZN(
        DP_reg_a_i_1_n75) );
  OAI21_X1 DP_reg_a_i_1_U5 ( .B1(DP_reg_a_i_1_n38), .B2(DP_reg_a_i_1_n63), .A(
        DP_reg_a_i_1_n75), .ZN(DP_reg_a_i_1_n51) );
  BUF_X1 DP_reg_a_i_1_U4 ( .A(vIn), .Z(DP_reg_a_i_1_n38) );
  BUF_X1 DP_reg_a_i_1_U3 ( .A(vIn), .Z(DP_reg_a_i_1_n37) );
  BUF_X1 DP_reg_a_i_1_U2 ( .A(DP_n1), .Z(DP_reg_a_i_1_n39) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_0_ ( .D(DP_reg_a_i_1_n51), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_coeff_ret0[1]), .QN(DP_reg_a_i_1_n63) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_1_ ( .D(DP_reg_a_i_1_n50), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__1_), .QN(DP_reg_a_i_1_n62) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_2_ ( .D(DP_reg_a_i_1_n49), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__2_), .QN(DP_reg_a_i_1_n61) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_3_ ( .D(DP_reg_a_i_1_n48), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__3_), .QN(DP_reg_a_i_1_n60) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_4_ ( .D(DP_reg_a_i_1_n47), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__4_), .QN(DP_reg_a_i_1_n59) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_5_ ( .D(DP_reg_a_i_1_n46), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__5_), .QN(DP_reg_a_i_1_n58) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_6_ ( .D(DP_reg_a_i_1_n45), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__6_), .QN(DP_reg_a_i_1_n57) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_7_ ( .D(DP_reg_a_i_1_n44), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__7_), .QN(DP_reg_a_i_1_n56) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_8_ ( .D(DP_reg_a_i_1_n43), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__8_), .QN(DP_reg_a_i_1_n55) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_9_ ( .D(DP_reg_a_i_1_n42), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__9_), .QN(DP_reg_a_i_1_n54) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_10_ ( .D(DP_reg_a_i_1_n41), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__10_), .QN(DP_reg_a_i_1_n53) );
  DFFR_X1 DP_reg_a_i_1_Q_reg_11_ ( .D(DP_reg_a_i_1_n40), .CK(clk), .RN(
        DP_reg_a_i_1_n39), .Q(DP_a_int_1__11_), .QN(DP_reg_a_i_1_n52) );
  NAND2_X1 DP_reg_a_i_2_U28 ( .A1(a[11]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n64) );
  OAI21_X1 DP_reg_a_i_2_U27 ( .B1(DP_reg_a_i_2_n37), .B2(DP_reg_a_i_2_n52), 
        .A(DP_reg_a_i_2_n64), .ZN(DP_reg_a_i_2_n40) );
  NAND2_X1 DP_reg_a_i_2_U26 ( .A1(a[10]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n65) );
  OAI21_X1 DP_reg_a_i_2_U25 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n53), 
        .A(DP_reg_a_i_2_n65), .ZN(DP_reg_a_i_2_n41) );
  NAND2_X1 DP_reg_a_i_2_U24 ( .A1(a[9]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n66) );
  OAI21_X1 DP_reg_a_i_2_U23 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n54), 
        .A(DP_reg_a_i_2_n66), .ZN(DP_reg_a_i_2_n42) );
  NAND2_X1 DP_reg_a_i_2_U22 ( .A1(a[8]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n67) );
  OAI21_X1 DP_reg_a_i_2_U21 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n55), 
        .A(DP_reg_a_i_2_n67), .ZN(DP_reg_a_i_2_n43) );
  NAND2_X1 DP_reg_a_i_2_U20 ( .A1(a[7]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n68) );
  OAI21_X1 DP_reg_a_i_2_U19 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n56), 
        .A(DP_reg_a_i_2_n68), .ZN(DP_reg_a_i_2_n44) );
  NAND2_X1 DP_reg_a_i_2_U18 ( .A1(a[6]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n69) );
  OAI21_X1 DP_reg_a_i_2_U17 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n57), 
        .A(DP_reg_a_i_2_n69), .ZN(DP_reg_a_i_2_n45) );
  NAND2_X1 DP_reg_a_i_2_U16 ( .A1(a[5]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n70) );
  OAI21_X1 DP_reg_a_i_2_U15 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n58), 
        .A(DP_reg_a_i_2_n70), .ZN(DP_reg_a_i_2_n46) );
  NAND2_X1 DP_reg_a_i_2_U14 ( .A1(a[4]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n71) );
  OAI21_X1 DP_reg_a_i_2_U13 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n59), 
        .A(DP_reg_a_i_2_n71), .ZN(DP_reg_a_i_2_n47) );
  NAND2_X1 DP_reg_a_i_2_U12 ( .A1(a[3]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n72) );
  OAI21_X1 DP_reg_a_i_2_U11 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n60), 
        .A(DP_reg_a_i_2_n72), .ZN(DP_reg_a_i_2_n48) );
  NAND2_X1 DP_reg_a_i_2_U10 ( .A1(a[2]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n73) );
  OAI21_X1 DP_reg_a_i_2_U9 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n61), .A(
        DP_reg_a_i_2_n73), .ZN(DP_reg_a_i_2_n49) );
  NAND2_X1 DP_reg_a_i_2_U8 ( .A1(a[1]), .A2(DP_reg_a_i_2_n37), .ZN(
        DP_reg_a_i_2_n74) );
  OAI21_X1 DP_reg_a_i_2_U7 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n62), .A(
        DP_reg_a_i_2_n74), .ZN(DP_reg_a_i_2_n50) );
  NAND2_X1 DP_reg_a_i_2_U6 ( .A1(DP_reg_a_i_2_n38), .A2(a[0]), .ZN(
        DP_reg_a_i_2_n75) );
  OAI21_X1 DP_reg_a_i_2_U5 ( .B1(DP_reg_a_i_2_n38), .B2(DP_reg_a_i_2_n63), .A(
        DP_reg_a_i_2_n75), .ZN(DP_reg_a_i_2_n51) );
  BUF_X1 DP_reg_a_i_2_U4 ( .A(vIn), .Z(DP_reg_a_i_2_n38) );
  BUF_X1 DP_reg_a_i_2_U3 ( .A(vIn), .Z(DP_reg_a_i_2_n37) );
  BUF_X1 DP_reg_a_i_2_U2 ( .A(DP_n2), .Z(DP_reg_a_i_2_n39) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_0_ ( .D(DP_reg_a_i_2_n51), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N37), .QN(DP_reg_a_i_2_n63) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_1_ ( .D(DP_reg_a_i_2_n50), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N38), .QN(DP_reg_a_i_2_n62) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_2_ ( .D(DP_reg_a_i_2_n49), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N39), .QN(DP_reg_a_i_2_n61) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_3_ ( .D(DP_reg_a_i_2_n48), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N40), .QN(DP_reg_a_i_2_n60) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_4_ ( .D(DP_reg_a_i_2_n47), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N41), .QN(DP_reg_a_i_2_n59) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_5_ ( .D(DP_reg_a_i_2_n46), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N42), .QN(DP_reg_a_i_2_n58) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_6_ ( .D(DP_reg_a_i_2_n45), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N43), .QN(DP_reg_a_i_2_n57) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_7_ ( .D(DP_reg_a_i_2_n44), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N44), .QN(DP_reg_a_i_2_n56) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_8_ ( .D(DP_reg_a_i_2_n43), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N45), .QN(DP_reg_a_i_2_n55) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_9_ ( .D(DP_reg_a_i_2_n42), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N46), .QN(DP_reg_a_i_2_n54) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_10_ ( .D(DP_reg_a_i_2_n41), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N47), .QN(DP_reg_a_i_2_n53) );
  DFFR_X1 DP_reg_a_i_2_Q_reg_11_ ( .D(DP_reg_a_i_2_n40), .CK(clk), .RN(
        DP_reg_a_i_2_n39), .Q(DP_N49), .QN(DP_reg_a_i_2_n52) );
  NAND2_X1 DP_reg_b_i_0_U28 ( .A1(b[35]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n64) );
  OAI21_X1 DP_reg_b_i_0_U27 ( .B1(DP_reg_b_i_0_n37), .B2(DP_reg_b_i_0_n52), 
        .A(DP_reg_b_i_0_n64), .ZN(DP_reg_b_i_0_n40) );
  NAND2_X1 DP_reg_b_i_0_U26 ( .A1(b[34]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n65) );
  OAI21_X1 DP_reg_b_i_0_U25 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n53), 
        .A(DP_reg_b_i_0_n65), .ZN(DP_reg_b_i_0_n41) );
  NAND2_X1 DP_reg_b_i_0_U24 ( .A1(b[33]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n66) );
  OAI21_X1 DP_reg_b_i_0_U23 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n54), 
        .A(DP_reg_b_i_0_n66), .ZN(DP_reg_b_i_0_n42) );
  NAND2_X1 DP_reg_b_i_0_U22 ( .A1(b[32]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n67) );
  OAI21_X1 DP_reg_b_i_0_U21 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n55), 
        .A(DP_reg_b_i_0_n67), .ZN(DP_reg_b_i_0_n43) );
  NAND2_X1 DP_reg_b_i_0_U20 ( .A1(b[31]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n68) );
  OAI21_X1 DP_reg_b_i_0_U19 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n56), 
        .A(DP_reg_b_i_0_n68), .ZN(DP_reg_b_i_0_n44) );
  NAND2_X1 DP_reg_b_i_0_U18 ( .A1(b[30]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n69) );
  OAI21_X1 DP_reg_b_i_0_U17 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n57), 
        .A(DP_reg_b_i_0_n69), .ZN(DP_reg_b_i_0_n45) );
  NAND2_X1 DP_reg_b_i_0_U16 ( .A1(b[29]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n70) );
  OAI21_X1 DP_reg_b_i_0_U15 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n58), 
        .A(DP_reg_b_i_0_n70), .ZN(DP_reg_b_i_0_n46) );
  NAND2_X1 DP_reg_b_i_0_U14 ( .A1(b[28]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n71) );
  OAI21_X1 DP_reg_b_i_0_U13 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n59), 
        .A(DP_reg_b_i_0_n71), .ZN(DP_reg_b_i_0_n47) );
  NAND2_X1 DP_reg_b_i_0_U12 ( .A1(b[27]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n72) );
  OAI21_X1 DP_reg_b_i_0_U11 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n60), 
        .A(DP_reg_b_i_0_n72), .ZN(DP_reg_b_i_0_n48) );
  NAND2_X1 DP_reg_b_i_0_U10 ( .A1(b[26]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n73) );
  OAI21_X1 DP_reg_b_i_0_U9 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n61), .A(
        DP_reg_b_i_0_n73), .ZN(DP_reg_b_i_0_n49) );
  NAND2_X1 DP_reg_b_i_0_U8 ( .A1(b[25]), .A2(DP_reg_b_i_0_n37), .ZN(
        DP_reg_b_i_0_n74) );
  OAI21_X1 DP_reg_b_i_0_U7 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n62), .A(
        DP_reg_b_i_0_n74), .ZN(DP_reg_b_i_0_n50) );
  NAND2_X1 DP_reg_b_i_0_U6 ( .A1(DP_reg_b_i_0_n38), .A2(b[24]), .ZN(
        DP_reg_b_i_0_n75) );
  OAI21_X1 DP_reg_b_i_0_U5 ( .B1(DP_reg_b_i_0_n38), .B2(DP_reg_b_i_0_n63), .A(
        DP_reg_b_i_0_n75), .ZN(DP_reg_b_i_0_n51) );
  BUF_X1 DP_reg_b_i_0_U4 ( .A(vIn), .Z(DP_reg_b_i_0_n38) );
  BUF_X1 DP_reg_b_i_0_U3 ( .A(vIn), .Z(DP_reg_b_i_0_n37) );
  BUF_X1 DP_reg_b_i_0_U2 ( .A(DP_n3), .Z(DP_reg_b_i_0_n39) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_0_ ( .D(DP_reg_b_i_0_n51), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__0_), .QN(DP_reg_b_i_0_n63) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_1_ ( .D(DP_reg_b_i_0_n50), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__1_), .QN(DP_reg_b_i_0_n62) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_2_ ( .D(DP_reg_b_i_0_n49), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__2_), .QN(DP_reg_b_i_0_n61) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_3_ ( .D(DP_reg_b_i_0_n48), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__3_), .QN(DP_reg_b_i_0_n60) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_4_ ( .D(DP_reg_b_i_0_n47), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__4_), .QN(DP_reg_b_i_0_n59) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_5_ ( .D(DP_reg_b_i_0_n46), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__5_), .QN(DP_reg_b_i_0_n58) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_6_ ( .D(DP_reg_b_i_0_n45), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__6_), .QN(DP_reg_b_i_0_n57) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_7_ ( .D(DP_reg_b_i_0_n44), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__7_), .QN(DP_reg_b_i_0_n56) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_8_ ( .D(DP_reg_b_i_0_n43), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__8_), .QN(DP_reg_b_i_0_n55) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_9_ ( .D(DP_reg_b_i_0_n42), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__9_), .QN(DP_reg_b_i_0_n54) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_10_ ( .D(DP_reg_b_i_0_n41), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__10_), .QN(DP_reg_b_i_0_n53) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_11_ ( .D(DP_reg_b_i_0_n40), .CK(clk), .RN(
        DP_reg_b_i_0_n39), .Q(DP_b_int_0__11_), .QN(DP_reg_b_i_0_n52) );
  NAND2_X1 DP_reg_b_i_1_U28 ( .A1(b[23]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n64) );
  OAI21_X1 DP_reg_b_i_1_U27 ( .B1(DP_reg_b_i_1_n37), .B2(DP_reg_b_i_1_n52), 
        .A(DP_reg_b_i_1_n64), .ZN(DP_reg_b_i_1_n40) );
  NAND2_X1 DP_reg_b_i_1_U26 ( .A1(b[22]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n65) );
  OAI21_X1 DP_reg_b_i_1_U25 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n53), 
        .A(DP_reg_b_i_1_n65), .ZN(DP_reg_b_i_1_n41) );
  NAND2_X1 DP_reg_b_i_1_U24 ( .A1(b[21]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n66) );
  OAI21_X1 DP_reg_b_i_1_U23 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n54), 
        .A(DP_reg_b_i_1_n66), .ZN(DP_reg_b_i_1_n42) );
  NAND2_X1 DP_reg_b_i_1_U22 ( .A1(b[20]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n67) );
  OAI21_X1 DP_reg_b_i_1_U21 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n55), 
        .A(DP_reg_b_i_1_n67), .ZN(DP_reg_b_i_1_n43) );
  NAND2_X1 DP_reg_b_i_1_U20 ( .A1(b[19]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n68) );
  OAI21_X1 DP_reg_b_i_1_U19 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n56), 
        .A(DP_reg_b_i_1_n68), .ZN(DP_reg_b_i_1_n44) );
  NAND2_X1 DP_reg_b_i_1_U18 ( .A1(b[18]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n69) );
  OAI21_X1 DP_reg_b_i_1_U17 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n57), 
        .A(DP_reg_b_i_1_n69), .ZN(DP_reg_b_i_1_n45) );
  NAND2_X1 DP_reg_b_i_1_U16 ( .A1(b[17]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n70) );
  OAI21_X1 DP_reg_b_i_1_U15 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n58), 
        .A(DP_reg_b_i_1_n70), .ZN(DP_reg_b_i_1_n46) );
  NAND2_X1 DP_reg_b_i_1_U14 ( .A1(b[16]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n71) );
  OAI21_X1 DP_reg_b_i_1_U13 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n59), 
        .A(DP_reg_b_i_1_n71), .ZN(DP_reg_b_i_1_n47) );
  NAND2_X1 DP_reg_b_i_1_U12 ( .A1(b[15]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n72) );
  OAI21_X1 DP_reg_b_i_1_U11 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n60), 
        .A(DP_reg_b_i_1_n72), .ZN(DP_reg_b_i_1_n48) );
  NAND2_X1 DP_reg_b_i_1_U10 ( .A1(b[14]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n73) );
  OAI21_X1 DP_reg_b_i_1_U9 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n61), .A(
        DP_reg_b_i_1_n73), .ZN(DP_reg_b_i_1_n49) );
  NAND2_X1 DP_reg_b_i_1_U8 ( .A1(b[13]), .A2(DP_reg_b_i_1_n37), .ZN(
        DP_reg_b_i_1_n74) );
  OAI21_X1 DP_reg_b_i_1_U7 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n62), .A(
        DP_reg_b_i_1_n74), .ZN(DP_reg_b_i_1_n50) );
  NAND2_X1 DP_reg_b_i_1_U6 ( .A1(DP_reg_b_i_1_n38), .A2(b[12]), .ZN(
        DP_reg_b_i_1_n75) );
  OAI21_X1 DP_reg_b_i_1_U5 ( .B1(DP_reg_b_i_1_n38), .B2(DP_reg_b_i_1_n63), .A(
        DP_reg_b_i_1_n75), .ZN(DP_reg_b_i_1_n51) );
  BUF_X1 DP_reg_b_i_1_U4 ( .A(vIn), .Z(DP_reg_b_i_1_n38) );
  BUF_X1 DP_reg_b_i_1_U3 ( .A(vIn), .Z(DP_reg_b_i_1_n37) );
  BUF_X1 DP_reg_b_i_1_U2 ( .A(DP_n4), .Z(DP_reg_b_i_1_n39) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_0_ ( .D(DP_reg_b_i_1_n51), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__0_), .QN(DP_reg_b_i_1_n63) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_1_ ( .D(DP_reg_b_i_1_n50), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__1_), .QN(DP_reg_b_i_1_n62) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_2_ ( .D(DP_reg_b_i_1_n49), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__2_), .QN(DP_reg_b_i_1_n61) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_3_ ( .D(DP_reg_b_i_1_n48), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__3_), .QN(DP_reg_b_i_1_n60) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_4_ ( .D(DP_reg_b_i_1_n47), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__4_), .QN(DP_reg_b_i_1_n59) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_5_ ( .D(DP_reg_b_i_1_n46), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__5_), .QN(DP_reg_b_i_1_n58) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_6_ ( .D(DP_reg_b_i_1_n45), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__6_), .QN(DP_reg_b_i_1_n57) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_7_ ( .D(DP_reg_b_i_1_n44), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__7_), .QN(DP_reg_b_i_1_n56) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_8_ ( .D(DP_reg_b_i_1_n43), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__8_), .QN(DP_reg_b_i_1_n55) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_9_ ( .D(DP_reg_b_i_1_n42), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__9_), .QN(DP_reg_b_i_1_n54) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_10_ ( .D(DP_reg_b_i_1_n41), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__10_), .QN(DP_reg_b_i_1_n53) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_11_ ( .D(DP_reg_b_i_1_n40), .CK(clk), .RN(
        DP_reg_b_i_1_n39), .Q(DP_b_int_1__11_), .QN(DP_reg_b_i_1_n52) );
  NAND2_X1 DP_reg_b_i_2_U28 ( .A1(b[11]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n64) );
  OAI21_X1 DP_reg_b_i_2_U27 ( .B1(DP_reg_b_i_2_n37), .B2(DP_reg_b_i_2_n52), 
        .A(DP_reg_b_i_2_n64), .ZN(DP_reg_b_i_2_n40) );
  NAND2_X1 DP_reg_b_i_2_U26 ( .A1(b[10]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n65) );
  OAI21_X1 DP_reg_b_i_2_U25 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n53), 
        .A(DP_reg_b_i_2_n65), .ZN(DP_reg_b_i_2_n41) );
  NAND2_X1 DP_reg_b_i_2_U24 ( .A1(b[9]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n66) );
  OAI21_X1 DP_reg_b_i_2_U23 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n54), 
        .A(DP_reg_b_i_2_n66), .ZN(DP_reg_b_i_2_n42) );
  NAND2_X1 DP_reg_b_i_2_U22 ( .A1(b[8]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n67) );
  OAI21_X1 DP_reg_b_i_2_U21 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n55), 
        .A(DP_reg_b_i_2_n67), .ZN(DP_reg_b_i_2_n43) );
  NAND2_X1 DP_reg_b_i_2_U20 ( .A1(b[7]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n68) );
  OAI21_X1 DP_reg_b_i_2_U19 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n56), 
        .A(DP_reg_b_i_2_n68), .ZN(DP_reg_b_i_2_n44) );
  NAND2_X1 DP_reg_b_i_2_U18 ( .A1(b[6]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n69) );
  OAI21_X1 DP_reg_b_i_2_U17 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n57), 
        .A(DP_reg_b_i_2_n69), .ZN(DP_reg_b_i_2_n45) );
  NAND2_X1 DP_reg_b_i_2_U16 ( .A1(b[5]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n70) );
  OAI21_X1 DP_reg_b_i_2_U15 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n58), 
        .A(DP_reg_b_i_2_n70), .ZN(DP_reg_b_i_2_n46) );
  NAND2_X1 DP_reg_b_i_2_U14 ( .A1(b[4]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n71) );
  OAI21_X1 DP_reg_b_i_2_U13 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n59), 
        .A(DP_reg_b_i_2_n71), .ZN(DP_reg_b_i_2_n47) );
  NAND2_X1 DP_reg_b_i_2_U12 ( .A1(b[3]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n72) );
  OAI21_X1 DP_reg_b_i_2_U11 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n60), 
        .A(DP_reg_b_i_2_n72), .ZN(DP_reg_b_i_2_n48) );
  NAND2_X1 DP_reg_b_i_2_U10 ( .A1(b[2]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n73) );
  OAI21_X1 DP_reg_b_i_2_U9 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n61), .A(
        DP_reg_b_i_2_n73), .ZN(DP_reg_b_i_2_n49) );
  NAND2_X1 DP_reg_b_i_2_U8 ( .A1(b[1]), .A2(DP_reg_b_i_2_n37), .ZN(
        DP_reg_b_i_2_n74) );
  OAI21_X1 DP_reg_b_i_2_U7 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n62), .A(
        DP_reg_b_i_2_n74), .ZN(DP_reg_b_i_2_n50) );
  NAND2_X1 DP_reg_b_i_2_U6 ( .A1(DP_reg_b_i_2_n38), .A2(b[0]), .ZN(
        DP_reg_b_i_2_n75) );
  OAI21_X1 DP_reg_b_i_2_U5 ( .B1(DP_reg_b_i_2_n38), .B2(DP_reg_b_i_2_n63), .A(
        DP_reg_b_i_2_n75), .ZN(DP_reg_b_i_2_n51) );
  BUF_X1 DP_reg_b_i_2_U4 ( .A(vIn), .Z(DP_reg_b_i_2_n38) );
  BUF_X1 DP_reg_b_i_2_U3 ( .A(vIn), .Z(DP_reg_b_i_2_n37) );
  BUF_X1 DP_reg_b_i_2_U2 ( .A(DP_n5), .Z(DP_reg_b_i_2_n39) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_0_ ( .D(DP_reg_b_i_2_n51), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__0_), .QN(DP_reg_b_i_2_n63) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_1_ ( .D(DP_reg_b_i_2_n50), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__1_), .QN(DP_reg_b_i_2_n62) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_2_ ( .D(DP_reg_b_i_2_n49), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__2_), .QN(DP_reg_b_i_2_n61) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_3_ ( .D(DP_reg_b_i_2_n48), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__3_), .QN(DP_reg_b_i_2_n60) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_4_ ( .D(DP_reg_b_i_2_n47), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__4_), .QN(DP_reg_b_i_2_n59) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_5_ ( .D(DP_reg_b_i_2_n46), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__5_), .QN(DP_reg_b_i_2_n58) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_6_ ( .D(DP_reg_b_i_2_n45), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__6_), .QN(DP_reg_b_i_2_n57) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_7_ ( .D(DP_reg_b_i_2_n44), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__7_), .QN(DP_reg_b_i_2_n56) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_8_ ( .D(DP_reg_b_i_2_n43), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__8_), .QN(DP_reg_b_i_2_n55) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_9_ ( .D(DP_reg_b_i_2_n42), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__9_), .QN(DP_reg_b_i_2_n54) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_10_ ( .D(DP_reg_b_i_2_n41), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__10_), .QN(DP_reg_b_i_2_n53) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_11_ ( .D(DP_reg_b_i_2_n40), .CK(clk), .RN(
        DP_reg_b_i_2_n39), .Q(DP_b_int_2__11_), .QN(DP_reg_b_i_2_n52) );
  NAND2_X1 DP_reg_sw0_U57 ( .A1(DP_w_6_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n7) );
  OAI21_X1 DP_reg_sw0_U56 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n31), .A(
        DP_reg_sw0_n7), .ZN(DP_reg_sw0_n55) );
  NAND2_X1 DP_reg_sw0_U55 ( .A1(DP_w_3_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n4) );
  OAI21_X1 DP_reg_sw0_U54 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n28), .A(
        DP_reg_sw0_n4), .ZN(DP_reg_sw0_n52) );
  NAND2_X1 DP_reg_sw0_U53 ( .A1(DP_w_2_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n3) );
  OAI21_X1 DP_reg_sw0_U52 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n27), .A(
        DP_reg_sw0_n3), .ZN(DP_reg_sw0_n51) );
  NAND2_X1 DP_reg_sw0_U51 ( .A1(DP_w_1_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n2) );
  OAI21_X1 DP_reg_sw0_U50 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n26), .A(
        DP_reg_sw0_n2), .ZN(DP_reg_sw0_n50) );
  NAND2_X1 DP_reg_sw0_U49 ( .A1(DP_reg_sw0_n78), .A2(DP_w_0_), .ZN(
        DP_reg_sw0_n1) );
  OAI21_X1 DP_reg_sw0_U48 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n25), .A(
        DP_reg_sw0_n1), .ZN(DP_reg_sw0_n49) );
  NAND2_X1 DP_reg_sw0_U47 ( .A1(DP_w_5_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n6) );
  OAI21_X1 DP_reg_sw0_U46 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n30), .A(
        DP_reg_sw0_n6), .ZN(DP_reg_sw0_n54) );
  NAND2_X1 DP_reg_sw0_U45 ( .A1(DP_w_4_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n5) );
  OAI21_X1 DP_reg_sw0_U44 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n29), .A(
        DP_reg_sw0_n5), .ZN(DP_reg_sw0_n53) );
  NAND2_X1 DP_reg_sw0_U43 ( .A1(DP_w_13_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n14) );
  OAI21_X1 DP_reg_sw0_U42 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n38), .A(
        DP_reg_sw0_n14), .ZN(DP_reg_sw0_n62) );
  NAND2_X1 DP_reg_sw0_U41 ( .A1(DP_w_12_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n13) );
  OAI21_X1 DP_reg_sw0_U40 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n37), .A(
        DP_reg_sw0_n13), .ZN(DP_reg_sw0_n61) );
  NAND2_X1 DP_reg_sw0_U39 ( .A1(DP_w_11_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n12) );
  OAI21_X1 DP_reg_sw0_U38 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n36), .A(
        DP_reg_sw0_n12), .ZN(DP_reg_sw0_n60) );
  NAND2_X1 DP_reg_sw0_U37 ( .A1(DP_w_16_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n17) );
  OAI21_X1 DP_reg_sw0_U36 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n41), .A(
        DP_reg_sw0_n17), .ZN(DP_reg_sw0_n65) );
  NAND2_X1 DP_reg_sw0_U35 ( .A1(DP_w_15_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n16) );
  OAI21_X1 DP_reg_sw0_U34 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n40), .A(
        DP_reg_sw0_n16), .ZN(DP_reg_sw0_n64) );
  NAND2_X1 DP_reg_sw0_U33 ( .A1(DP_w_14_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n15) );
  OAI21_X1 DP_reg_sw0_U32 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n39), .A(
        DP_reg_sw0_n15), .ZN(DP_reg_sw0_n63) );
  NAND2_X1 DP_reg_sw0_U31 ( .A1(DP_w_10_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n11) );
  OAI21_X1 DP_reg_sw0_U30 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n35), .A(
        DP_reg_sw0_n11), .ZN(DP_reg_sw0_n59) );
  NAND2_X1 DP_reg_sw0_U29 ( .A1(DP_w_9_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n10) );
  OAI21_X1 DP_reg_sw0_U28 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n34), .A(
        DP_reg_sw0_n10), .ZN(DP_reg_sw0_n58) );
  NAND2_X1 DP_reg_sw0_U27 ( .A1(DP_w_8_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n9) );
  OAI21_X1 DP_reg_sw0_U26 ( .B1(DP_reg_sw0_n76), .B2(DP_reg_sw0_n33), .A(
        DP_reg_sw0_n9), .ZN(DP_reg_sw0_n57) );
  NAND2_X1 DP_reg_sw0_U25 ( .A1(DP_w_7_), .A2(DP_reg_sw0_n76), .ZN(
        DP_reg_sw0_n8) );
  OAI21_X1 DP_reg_sw0_U24 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n32), .A(
        DP_reg_sw0_n8), .ZN(DP_reg_sw0_n56) );
  NAND2_X1 DP_reg_sw0_U23 ( .A1(DP_w_23_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n24) );
  OAI21_X1 DP_reg_sw0_U22 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n48), .A(
        DP_reg_sw0_n24), .ZN(DP_reg_sw0_n72) );
  NAND2_X1 DP_reg_sw0_U21 ( .A1(DP_w_22_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n23) );
  OAI21_X1 DP_reg_sw0_U20 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n47), .A(
        DP_reg_sw0_n23), .ZN(DP_reg_sw0_n71) );
  NAND2_X1 DP_reg_sw0_U19 ( .A1(DP_w_20_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n21) );
  OAI21_X1 DP_reg_sw0_U18 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n45), .A(
        DP_reg_sw0_n21), .ZN(DP_reg_sw0_n69) );
  NAND2_X1 DP_reg_sw0_U17 ( .A1(DP_w_19_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n20) );
  OAI21_X1 DP_reg_sw0_U16 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n44), .A(
        DP_reg_sw0_n20), .ZN(DP_reg_sw0_n68) );
  NAND2_X1 DP_reg_sw0_U15 ( .A1(DP_w_18_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n19) );
  OAI21_X1 DP_reg_sw0_U14 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n43), .A(
        DP_reg_sw0_n19), .ZN(DP_reg_sw0_n67) );
  NAND2_X1 DP_reg_sw0_U13 ( .A1(DP_w_17_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n18) );
  OAI21_X1 DP_reg_sw0_U12 ( .B1(DP_reg_sw0_n77), .B2(DP_reg_sw0_n42), .A(
        DP_reg_sw0_n18), .ZN(DP_reg_sw0_n66) );
  NAND2_X1 DP_reg_sw0_U11 ( .A1(DP_w_21_), .A2(DP_reg_sw0_n75), .ZN(
        DP_reg_sw0_n22) );
  OAI21_X1 DP_reg_sw0_U10 ( .B1(DP_reg_sw0_n78), .B2(DP_reg_sw0_n46), .A(
        DP_reg_sw0_n22), .ZN(DP_reg_sw0_n70) );
  BUF_X1 DP_reg_sw0_U9 ( .A(DP_n1), .Z(DP_reg_sw0_n79) );
  BUF_X1 DP_reg_sw0_U8 ( .A(DP_n1), .Z(DP_reg_sw0_n80) );
  BUF_X1 DP_reg_sw0_U7 ( .A(sw_regs_en_int), .Z(DP_reg_sw0_n74) );
  BUF_X1 DP_reg_sw0_U6 ( .A(sw_regs_en_int), .Z(DP_reg_sw0_n73) );
  BUF_X1 DP_reg_sw0_U5 ( .A(DP_reg_sw0_n74), .Z(DP_reg_sw0_n78) );
  BUF_X1 DP_reg_sw0_U4 ( .A(DP_reg_sw0_n73), .Z(DP_reg_sw0_n76) );
  BUF_X1 DP_reg_sw0_U3 ( .A(DP_reg_sw0_n74), .Z(DP_reg_sw0_n77) );
  BUF_X1 DP_reg_sw0_U2 ( .A(DP_reg_sw0_n73), .Z(DP_reg_sw0_n75) );
  DFFR_X1 DP_reg_sw0_Q_reg_0_ ( .D(DP_reg_sw0_n49), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_0_), .QN(DP_reg_sw0_n25) );
  DFFR_X1 DP_reg_sw0_Q_reg_1_ ( .D(DP_reg_sw0_n50), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_1_), .QN(DP_reg_sw0_n26) );
  DFFR_X1 DP_reg_sw0_Q_reg_2_ ( .D(DP_reg_sw0_n51), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_2_), .QN(DP_reg_sw0_n27) );
  DFFR_X1 DP_reg_sw0_Q_reg_3_ ( .D(DP_reg_sw0_n52), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_3_), .QN(DP_reg_sw0_n28) );
  DFFR_X1 DP_reg_sw0_Q_reg_4_ ( .D(DP_reg_sw0_n53), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_4_), .QN(DP_reg_sw0_n29) );
  DFFR_X1 DP_reg_sw0_Q_reg_5_ ( .D(DP_reg_sw0_n54), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_5_), .QN(DP_reg_sw0_n30) );
  DFFR_X1 DP_reg_sw0_Q_reg_6_ ( .D(DP_reg_sw0_n55), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_6_), .QN(DP_reg_sw0_n31) );
  DFFR_X1 DP_reg_sw0_Q_reg_7_ ( .D(DP_reg_sw0_n56), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_7_), .QN(DP_reg_sw0_n32) );
  DFFR_X1 DP_reg_sw0_Q_reg_8_ ( .D(DP_reg_sw0_n57), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_8_), .QN(DP_reg_sw0_n33) );
  DFFR_X1 DP_reg_sw0_Q_reg_9_ ( .D(DP_reg_sw0_n58), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_9_), .QN(DP_reg_sw0_n34) );
  DFFR_X1 DP_reg_sw0_Q_reg_10_ ( .D(DP_reg_sw0_n59), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_10_), .QN(DP_reg_sw0_n35) );
  DFFR_X1 DP_reg_sw0_Q_reg_11_ ( .D(DP_reg_sw0_n60), .CK(clk), .RN(
        DP_reg_sw0_n80), .Q(DP_sw0_11_), .QN(DP_reg_sw0_n36) );
  DFFR_X1 DP_reg_sw0_Q_reg_12_ ( .D(DP_reg_sw0_n61), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_12_), .QN(DP_reg_sw0_n37) );
  DFFR_X1 DP_reg_sw0_Q_reg_13_ ( .D(DP_reg_sw0_n62), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_13_), .QN(DP_reg_sw0_n38) );
  DFFR_X1 DP_reg_sw0_Q_reg_14_ ( .D(DP_reg_sw0_n63), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_14_), .QN(DP_reg_sw0_n39) );
  DFFR_X1 DP_reg_sw0_Q_reg_15_ ( .D(DP_reg_sw0_n64), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_15_), .QN(DP_reg_sw0_n40) );
  DFFR_X1 DP_reg_sw0_Q_reg_16_ ( .D(DP_reg_sw0_n65), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_16_), .QN(DP_reg_sw0_n41) );
  DFFR_X1 DP_reg_sw0_Q_reg_17_ ( .D(DP_reg_sw0_n66), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_17_), .QN(DP_reg_sw0_n42) );
  DFFR_X1 DP_reg_sw0_Q_reg_18_ ( .D(DP_reg_sw0_n67), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_18_), .QN(DP_reg_sw0_n43) );
  DFFR_X1 DP_reg_sw0_Q_reg_19_ ( .D(DP_reg_sw0_n68), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_19_), .QN(DP_reg_sw0_n44) );
  DFFR_X1 DP_reg_sw0_Q_reg_20_ ( .D(DP_reg_sw0_n69), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_20_), .QN(DP_reg_sw0_n45) );
  DFFR_X1 DP_reg_sw0_Q_reg_21_ ( .D(DP_reg_sw0_n70), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_21_), .QN(DP_reg_sw0_n46) );
  DFFR_X1 DP_reg_sw0_Q_reg_22_ ( .D(DP_reg_sw0_n71), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_22_), .QN(DP_reg_sw0_n47) );
  DFFR_X1 DP_reg_sw0_Q_reg_23_ ( .D(DP_reg_sw0_n72), .CK(clk), .RN(
        DP_reg_sw0_n79), .Q(DP_sw0_23_), .QN(DP_reg_sw0_n48) );
  NAND2_X1 DP_reg_sw1_U57 ( .A1(DP_sw0_23_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n129) );
  OAI21_X1 DP_reg_sw1_U56 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n105), .A(
        DP_reg_sw1_n129), .ZN(DP_reg_sw1_n81) );
  NAND2_X1 DP_reg_sw1_U55 ( .A1(DP_sw0_22_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n130) );
  OAI21_X1 DP_reg_sw1_U54 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n106), .A(
        DP_reg_sw1_n130), .ZN(DP_reg_sw1_n82) );
  NAND2_X1 DP_reg_sw1_U53 ( .A1(DP_sw0_20_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n132) );
  OAI21_X1 DP_reg_sw1_U52 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n108), .A(
        DP_reg_sw1_n132), .ZN(DP_reg_sw1_n84) );
  NAND2_X1 DP_reg_sw1_U51 ( .A1(DP_sw0_19_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n133) );
  OAI21_X1 DP_reg_sw1_U50 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n109), .A(
        DP_reg_sw1_n133), .ZN(DP_reg_sw1_n85) );
  NAND2_X1 DP_reg_sw1_U49 ( .A1(DP_sw0_6_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n146) );
  OAI21_X1 DP_reg_sw1_U48 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n122), .A(
        DP_reg_sw1_n146), .ZN(DP_reg_sw1_n98) );
  NAND2_X1 DP_reg_sw1_U47 ( .A1(DP_sw0_3_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n149) );
  OAI21_X1 DP_reg_sw1_U46 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n125), .A(
        DP_reg_sw1_n149), .ZN(DP_reg_sw1_n101) );
  NAND2_X1 DP_reg_sw1_U45 ( .A1(DP_sw0_2_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n150) );
  OAI21_X1 DP_reg_sw1_U44 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n126), .A(
        DP_reg_sw1_n150), .ZN(DP_reg_sw1_n102) );
  NAND2_X1 DP_reg_sw1_U43 ( .A1(DP_sw0_1_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n151) );
  OAI21_X1 DP_reg_sw1_U42 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n127), .A(
        DP_reg_sw1_n151), .ZN(DP_reg_sw1_n103) );
  NAND2_X1 DP_reg_sw1_U41 ( .A1(DP_reg_sw1_n78), .A2(DP_sw0_0_), .ZN(
        DP_reg_sw1_n152) );
  OAI21_X1 DP_reg_sw1_U40 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n128), .A(
        DP_reg_sw1_n152), .ZN(DP_reg_sw1_n104) );
  NAND2_X1 DP_reg_sw1_U39 ( .A1(DP_sw0_8_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n144) );
  OAI21_X1 DP_reg_sw1_U38 ( .B1(DP_reg_sw1_n76), .B2(DP_reg_sw1_n120), .A(
        DP_reg_sw1_n144), .ZN(DP_reg_sw1_n96) );
  NAND2_X1 DP_reg_sw1_U37 ( .A1(DP_sw0_18_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n134) );
  OAI21_X1 DP_reg_sw1_U36 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n110), .A(
        DP_reg_sw1_n134), .ZN(DP_reg_sw1_n86) );
  NAND2_X1 DP_reg_sw1_U35 ( .A1(DP_sw0_17_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n135) );
  OAI21_X1 DP_reg_sw1_U34 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n111), .A(
        DP_reg_sw1_n135), .ZN(DP_reg_sw1_n87) );
  NAND2_X1 DP_reg_sw1_U33 ( .A1(DP_sw0_16_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n136) );
  OAI21_X1 DP_reg_sw1_U32 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n112), .A(
        DP_reg_sw1_n136), .ZN(DP_reg_sw1_n88) );
  NAND2_X1 DP_reg_sw1_U31 ( .A1(DP_sw0_15_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n137) );
  OAI21_X1 DP_reg_sw1_U30 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n113), .A(
        DP_reg_sw1_n137), .ZN(DP_reg_sw1_n89) );
  NAND2_X1 DP_reg_sw1_U29 ( .A1(DP_sw0_14_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n138) );
  OAI21_X1 DP_reg_sw1_U28 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n114), .A(
        DP_reg_sw1_n138), .ZN(DP_reg_sw1_n90) );
  NAND2_X1 DP_reg_sw1_U27 ( .A1(DP_sw0_13_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n139) );
  OAI21_X1 DP_reg_sw1_U26 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n115), .A(
        DP_reg_sw1_n139), .ZN(DP_reg_sw1_n91) );
  NAND2_X1 DP_reg_sw1_U25 ( .A1(DP_sw0_12_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n140) );
  OAI21_X1 DP_reg_sw1_U24 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n116), .A(
        DP_reg_sw1_n140), .ZN(DP_reg_sw1_n92) );
  NAND2_X1 DP_reg_sw1_U23 ( .A1(DP_sw0_11_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n141) );
  OAI21_X1 DP_reg_sw1_U22 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n117), .A(
        DP_reg_sw1_n141), .ZN(DP_reg_sw1_n93) );
  NAND2_X1 DP_reg_sw1_U21 ( .A1(DP_sw0_10_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n142) );
  OAI21_X1 DP_reg_sw1_U20 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n118), .A(
        DP_reg_sw1_n142), .ZN(DP_reg_sw1_n94) );
  NAND2_X1 DP_reg_sw1_U19 ( .A1(DP_sw0_9_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n143) );
  OAI21_X1 DP_reg_sw1_U18 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n119), .A(
        DP_reg_sw1_n143), .ZN(DP_reg_sw1_n95) );
  NAND2_X1 DP_reg_sw1_U17 ( .A1(DP_sw0_7_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n145) );
  OAI21_X1 DP_reg_sw1_U16 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n121), .A(
        DP_reg_sw1_n145), .ZN(DP_reg_sw1_n97) );
  NAND2_X1 DP_reg_sw1_U15 ( .A1(DP_sw0_5_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n147) );
  OAI21_X1 DP_reg_sw1_U14 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n123), .A(
        DP_reg_sw1_n147), .ZN(DP_reg_sw1_n99) );
  NAND2_X1 DP_reg_sw1_U13 ( .A1(DP_sw0_4_), .A2(DP_reg_sw1_n76), .ZN(
        DP_reg_sw1_n148) );
  OAI21_X1 DP_reg_sw1_U12 ( .B1(DP_reg_sw1_n77), .B2(DP_reg_sw1_n124), .A(
        DP_reg_sw1_n148), .ZN(DP_reg_sw1_n100) );
  NAND2_X1 DP_reg_sw1_U11 ( .A1(DP_sw0_21_), .A2(DP_reg_sw1_n75), .ZN(
        DP_reg_sw1_n131) );
  OAI21_X1 DP_reg_sw1_U10 ( .B1(DP_reg_sw1_n78), .B2(DP_reg_sw1_n107), .A(
        DP_reg_sw1_n131), .ZN(DP_reg_sw1_n83) );
  BUF_X1 DP_reg_sw1_U9 ( .A(DP_n4), .Z(DP_reg_sw1_n79) );
  BUF_X1 DP_reg_sw1_U8 ( .A(DP_n4), .Z(DP_reg_sw1_n80) );
  BUF_X1 DP_reg_sw1_U7 ( .A(sw_regs_en_int), .Z(DP_reg_sw1_n74) );
  BUF_X1 DP_reg_sw1_U6 ( .A(sw_regs_en_int), .Z(DP_reg_sw1_n73) );
  BUF_X1 DP_reg_sw1_U5 ( .A(DP_reg_sw1_n74), .Z(DP_reg_sw1_n78) );
  BUF_X1 DP_reg_sw1_U4 ( .A(DP_reg_sw1_n73), .Z(DP_reg_sw1_n76) );
  BUF_X1 DP_reg_sw1_U3 ( .A(DP_reg_sw1_n74), .Z(DP_reg_sw1_n77) );
  BUF_X1 DP_reg_sw1_U2 ( .A(DP_reg_sw1_n73), .Z(DP_reg_sw1_n75) );
  DFFR_X1 DP_reg_sw1_Q_reg_0_ ( .D(DP_reg_sw1_n104), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_0_), .QN(DP_reg_sw1_n128) );
  DFFR_X1 DP_reg_sw1_Q_reg_1_ ( .D(DP_reg_sw1_n103), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_1_), .QN(DP_reg_sw1_n127) );
  DFFR_X1 DP_reg_sw1_Q_reg_2_ ( .D(DP_reg_sw1_n102), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_2_), .QN(DP_reg_sw1_n126) );
  DFFR_X1 DP_reg_sw1_Q_reg_3_ ( .D(DP_reg_sw1_n101), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_3_), .QN(DP_reg_sw1_n125) );
  DFFR_X1 DP_reg_sw1_Q_reg_4_ ( .D(DP_reg_sw1_n100), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_4_), .QN(DP_reg_sw1_n124) );
  DFFR_X1 DP_reg_sw1_Q_reg_5_ ( .D(DP_reg_sw1_n99), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_5_), .QN(DP_reg_sw1_n123) );
  DFFR_X1 DP_reg_sw1_Q_reg_6_ ( .D(DP_reg_sw1_n98), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_6_), .QN(DP_reg_sw1_n122) );
  DFFR_X1 DP_reg_sw1_Q_reg_7_ ( .D(DP_reg_sw1_n97), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_7_), .QN(DP_reg_sw1_n121) );
  DFFR_X1 DP_reg_sw1_Q_reg_8_ ( .D(DP_reg_sw1_n96), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_8_), .QN(DP_reg_sw1_n120) );
  DFFR_X1 DP_reg_sw1_Q_reg_9_ ( .D(DP_reg_sw1_n95), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_9_), .QN(DP_reg_sw1_n119) );
  DFFR_X1 DP_reg_sw1_Q_reg_10_ ( .D(DP_reg_sw1_n94), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_10_), .QN(DP_reg_sw1_n118) );
  DFFR_X1 DP_reg_sw1_Q_reg_11_ ( .D(DP_reg_sw1_n93), .CK(clk), .RN(
        DP_reg_sw1_n80), .Q(DP_sw1_11_), .QN(DP_reg_sw1_n117) );
  DFFR_X1 DP_reg_sw1_Q_reg_12_ ( .D(DP_reg_sw1_n92), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_12_), .QN(DP_reg_sw1_n116) );
  DFFR_X1 DP_reg_sw1_Q_reg_13_ ( .D(DP_reg_sw1_n91), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_13_), .QN(DP_reg_sw1_n115) );
  DFFR_X1 DP_reg_sw1_Q_reg_14_ ( .D(DP_reg_sw1_n90), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_14_), .QN(DP_reg_sw1_n114) );
  DFFR_X1 DP_reg_sw1_Q_reg_15_ ( .D(DP_reg_sw1_n89), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_15_), .QN(DP_reg_sw1_n113) );
  DFFR_X1 DP_reg_sw1_Q_reg_16_ ( .D(DP_reg_sw1_n88), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_16_), .QN(DP_reg_sw1_n112) );
  DFFR_X1 DP_reg_sw1_Q_reg_17_ ( .D(DP_reg_sw1_n87), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_17_), .QN(DP_reg_sw1_n111) );
  DFFR_X1 DP_reg_sw1_Q_reg_18_ ( .D(DP_reg_sw1_n86), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_18_), .QN(DP_reg_sw1_n110) );
  DFFR_X1 DP_reg_sw1_Q_reg_19_ ( .D(DP_reg_sw1_n85), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_19_), .QN(DP_reg_sw1_n109) );
  DFFR_X1 DP_reg_sw1_Q_reg_20_ ( .D(DP_reg_sw1_n84), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_20_), .QN(DP_reg_sw1_n108) );
  DFFR_X1 DP_reg_sw1_Q_reg_21_ ( .D(DP_reg_sw1_n83), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_21_), .QN(DP_reg_sw1_n107) );
  DFFR_X1 DP_reg_sw1_Q_reg_22_ ( .D(DP_reg_sw1_n82), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_22_), .QN(DP_reg_sw1_n106) );
  DFFR_X1 DP_reg_sw1_Q_reg_23_ ( .D(DP_reg_sw1_n81), .CK(clk), .RN(
        DP_reg_sw1_n79), .Q(DP_sw1_23_), .QN(DP_reg_sw1_n105) );
  NAND2_X1 DP_reg_sw2_U57 ( .A1(DP_sw1_23_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n129) );
  OAI21_X1 DP_reg_sw2_U56 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n105), .A(
        DP_reg_sw2_n129), .ZN(DP_reg_sw2_n81) );
  NAND2_X1 DP_reg_sw2_U55 ( .A1(DP_sw1_22_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n130) );
  OAI21_X1 DP_reg_sw2_U54 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n106), .A(
        DP_reg_sw2_n130), .ZN(DP_reg_sw2_n82) );
  NAND2_X1 DP_reg_sw2_U53 ( .A1(DP_sw1_20_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n132) );
  OAI21_X1 DP_reg_sw2_U52 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n108), .A(
        DP_reg_sw2_n132), .ZN(DP_reg_sw2_n84) );
  NAND2_X1 DP_reg_sw2_U51 ( .A1(DP_sw1_19_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n133) );
  OAI21_X1 DP_reg_sw2_U50 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n109), .A(
        DP_reg_sw2_n133), .ZN(DP_reg_sw2_n85) );
  NAND2_X1 DP_reg_sw2_U49 ( .A1(DP_sw1_6_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n146) );
  OAI21_X1 DP_reg_sw2_U48 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n122), .A(
        DP_reg_sw2_n146), .ZN(DP_reg_sw2_n98) );
  NAND2_X1 DP_reg_sw2_U47 ( .A1(DP_sw1_3_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n149) );
  OAI21_X1 DP_reg_sw2_U46 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n125), .A(
        DP_reg_sw2_n149), .ZN(DP_reg_sw2_n101) );
  NAND2_X1 DP_reg_sw2_U45 ( .A1(DP_sw1_2_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n150) );
  OAI21_X1 DP_reg_sw2_U44 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n126), .A(
        DP_reg_sw2_n150), .ZN(DP_reg_sw2_n102) );
  NAND2_X1 DP_reg_sw2_U43 ( .A1(DP_sw1_1_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n151) );
  OAI21_X1 DP_reg_sw2_U42 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n127), .A(
        DP_reg_sw2_n151), .ZN(DP_reg_sw2_n103) );
  NAND2_X1 DP_reg_sw2_U41 ( .A1(DP_reg_sw2_n78), .A2(DP_sw1_0_), .ZN(
        DP_reg_sw2_n152) );
  OAI21_X1 DP_reg_sw2_U40 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n128), .A(
        DP_reg_sw2_n152), .ZN(DP_reg_sw2_n104) );
  NAND2_X1 DP_reg_sw2_U39 ( .A1(DP_sw1_8_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n144) );
  OAI21_X1 DP_reg_sw2_U38 ( .B1(DP_reg_sw2_n76), .B2(DP_reg_sw2_n120), .A(
        DP_reg_sw2_n144), .ZN(DP_reg_sw2_n96) );
  NAND2_X1 DP_reg_sw2_U37 ( .A1(DP_sw1_18_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n134) );
  OAI21_X1 DP_reg_sw2_U36 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n110), .A(
        DP_reg_sw2_n134), .ZN(DP_reg_sw2_n86) );
  NAND2_X1 DP_reg_sw2_U35 ( .A1(DP_sw1_17_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n135) );
  OAI21_X1 DP_reg_sw2_U34 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n111), .A(
        DP_reg_sw2_n135), .ZN(DP_reg_sw2_n87) );
  NAND2_X1 DP_reg_sw2_U33 ( .A1(DP_sw1_16_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n136) );
  OAI21_X1 DP_reg_sw2_U32 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n112), .A(
        DP_reg_sw2_n136), .ZN(DP_reg_sw2_n88) );
  NAND2_X1 DP_reg_sw2_U31 ( .A1(DP_sw1_15_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n137) );
  OAI21_X1 DP_reg_sw2_U30 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n113), .A(
        DP_reg_sw2_n137), .ZN(DP_reg_sw2_n89) );
  NAND2_X1 DP_reg_sw2_U29 ( .A1(DP_sw1_14_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n138) );
  OAI21_X1 DP_reg_sw2_U28 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n114), .A(
        DP_reg_sw2_n138), .ZN(DP_reg_sw2_n90) );
  NAND2_X1 DP_reg_sw2_U27 ( .A1(DP_sw1_13_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n139) );
  OAI21_X1 DP_reg_sw2_U26 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n115), .A(
        DP_reg_sw2_n139), .ZN(DP_reg_sw2_n91) );
  NAND2_X1 DP_reg_sw2_U25 ( .A1(DP_sw1_12_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n140) );
  OAI21_X1 DP_reg_sw2_U24 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n116), .A(
        DP_reg_sw2_n140), .ZN(DP_reg_sw2_n92) );
  NAND2_X1 DP_reg_sw2_U23 ( .A1(DP_sw1_11_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n141) );
  OAI21_X1 DP_reg_sw2_U22 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n117), .A(
        DP_reg_sw2_n141), .ZN(DP_reg_sw2_n93) );
  NAND2_X1 DP_reg_sw2_U21 ( .A1(DP_sw1_10_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n142) );
  OAI21_X1 DP_reg_sw2_U20 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n118), .A(
        DP_reg_sw2_n142), .ZN(DP_reg_sw2_n94) );
  NAND2_X1 DP_reg_sw2_U19 ( .A1(DP_sw1_9_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n143) );
  OAI21_X1 DP_reg_sw2_U18 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n119), .A(
        DP_reg_sw2_n143), .ZN(DP_reg_sw2_n95) );
  NAND2_X1 DP_reg_sw2_U17 ( .A1(DP_sw1_7_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n145) );
  OAI21_X1 DP_reg_sw2_U16 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n121), .A(
        DP_reg_sw2_n145), .ZN(DP_reg_sw2_n97) );
  NAND2_X1 DP_reg_sw2_U15 ( .A1(DP_sw1_5_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n147) );
  OAI21_X1 DP_reg_sw2_U14 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n123), .A(
        DP_reg_sw2_n147), .ZN(DP_reg_sw2_n99) );
  NAND2_X1 DP_reg_sw2_U13 ( .A1(DP_sw1_4_), .A2(DP_reg_sw2_n76), .ZN(
        DP_reg_sw2_n148) );
  OAI21_X1 DP_reg_sw2_U12 ( .B1(DP_reg_sw2_n77), .B2(DP_reg_sw2_n124), .A(
        DP_reg_sw2_n148), .ZN(DP_reg_sw2_n100) );
  NAND2_X1 DP_reg_sw2_U11 ( .A1(DP_sw1_21_), .A2(DP_reg_sw2_n75), .ZN(
        DP_reg_sw2_n131) );
  OAI21_X1 DP_reg_sw2_U10 ( .B1(DP_reg_sw2_n78), .B2(DP_reg_sw2_n107), .A(
        DP_reg_sw2_n131), .ZN(DP_reg_sw2_n83) );
  BUF_X1 DP_reg_sw2_U9 ( .A(DP_n7), .Z(DP_reg_sw2_n79) );
  BUF_X1 DP_reg_sw2_U8 ( .A(DP_n7), .Z(DP_reg_sw2_n80) );
  BUF_X1 DP_reg_sw2_U7 ( .A(sw_regs_en_int), .Z(DP_reg_sw2_n74) );
  BUF_X1 DP_reg_sw2_U6 ( .A(sw_regs_en_int), .Z(DP_reg_sw2_n73) );
  BUF_X1 DP_reg_sw2_U5 ( .A(DP_reg_sw2_n74), .Z(DP_reg_sw2_n78) );
  BUF_X1 DP_reg_sw2_U4 ( .A(DP_reg_sw2_n73), .Z(DP_reg_sw2_n76) );
  BUF_X1 DP_reg_sw2_U3 ( .A(DP_reg_sw2_n74), .Z(DP_reg_sw2_n77) );
  BUF_X1 DP_reg_sw2_U2 ( .A(DP_reg_sw2_n73), .Z(DP_reg_sw2_n75) );
  DFFR_X1 DP_reg_sw2_Q_reg_0_ ( .D(DP_reg_sw2_n104), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[0]), .QN(DP_reg_sw2_n128) );
  DFFR_X1 DP_reg_sw2_Q_reg_1_ ( .D(DP_reg_sw2_n103), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[1]), .QN(DP_reg_sw2_n127) );
  DFFR_X1 DP_reg_sw2_Q_reg_2_ ( .D(DP_reg_sw2_n102), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[2]), .QN(DP_reg_sw2_n126) );
  DFFR_X1 DP_reg_sw2_Q_reg_3_ ( .D(DP_reg_sw2_n101), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[3]), .QN(DP_reg_sw2_n125) );
  DFFR_X1 DP_reg_sw2_Q_reg_4_ ( .D(DP_reg_sw2_n100), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[4]), .QN(DP_reg_sw2_n124) );
  DFFR_X1 DP_reg_sw2_Q_reg_5_ ( .D(DP_reg_sw2_n99), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[5]), .QN(DP_reg_sw2_n123) );
  DFFR_X1 DP_reg_sw2_Q_reg_6_ ( .D(DP_reg_sw2_n98), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[6]), .QN(DP_reg_sw2_n122) );
  DFFR_X1 DP_reg_sw2_Q_reg_7_ ( .D(DP_reg_sw2_n97), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[7]), .QN(DP_reg_sw2_n121) );
  DFFR_X1 DP_reg_sw2_Q_reg_8_ ( .D(DP_reg_sw2_n96), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[8]), .QN(DP_reg_sw2_n120) );
  DFFR_X1 DP_reg_sw2_Q_reg_9_ ( .D(DP_reg_sw2_n95), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[9]), .QN(DP_reg_sw2_n119) );
  DFFR_X1 DP_reg_sw2_Q_reg_10_ ( .D(DP_reg_sw2_n94), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[10]), .QN(DP_reg_sw2_n118) );
  DFFR_X1 DP_reg_sw2_Q_reg_11_ ( .D(DP_reg_sw2_n93), .CK(clk), .RN(
        DP_reg_sw2_n80), .Q(DP_sw2[11]), .QN(DP_reg_sw2_n117) );
  DFFR_X1 DP_reg_sw2_Q_reg_12_ ( .D(DP_reg_sw2_n92), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[12]), .QN(DP_reg_sw2_n116) );
  DFFR_X1 DP_reg_sw2_Q_reg_13_ ( .D(DP_reg_sw2_n91), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[13]), .QN(DP_reg_sw2_n115) );
  DFFR_X1 DP_reg_sw2_Q_reg_14_ ( .D(DP_reg_sw2_n90), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[14]), .QN(DP_reg_sw2_n114) );
  DFFR_X1 DP_reg_sw2_Q_reg_15_ ( .D(DP_reg_sw2_n89), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[15]), .QN(DP_reg_sw2_n113) );
  DFFR_X1 DP_reg_sw2_Q_reg_16_ ( .D(DP_reg_sw2_n88), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[16]), .QN(DP_reg_sw2_n112) );
  DFFR_X1 DP_reg_sw2_Q_reg_17_ ( .D(DP_reg_sw2_n87), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[17]), .QN(DP_reg_sw2_n111) );
  DFFR_X1 DP_reg_sw2_Q_reg_18_ ( .D(DP_reg_sw2_n86), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[18]), .QN(DP_reg_sw2_n110) );
  DFFR_X1 DP_reg_sw2_Q_reg_19_ ( .D(DP_reg_sw2_n85), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[19]), .QN(DP_reg_sw2_n109) );
  DFFR_X1 DP_reg_sw2_Q_reg_20_ ( .D(DP_reg_sw2_n84), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[20]), .QN(DP_reg_sw2_n108) );
  DFFR_X1 DP_reg_sw2_Q_reg_21_ ( .D(DP_reg_sw2_n83), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[21]), .QN(DP_reg_sw2_n107) );
  DFFR_X1 DP_reg_sw2_Q_reg_22_ ( .D(DP_reg_sw2_n82), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[22]), .QN(DP_reg_sw2_n106) );
  DFFR_X1 DP_reg_sw2_Q_reg_23_ ( .D(DP_reg_sw2_n81), .CK(clk), .RN(
        DP_reg_sw2_n79), .Q(DP_sw2[23]), .QN(DP_reg_sw2_n105) );
  NAND2_X1 DP_reg_ret0_U51 ( .A1(DP_sw0_coeff_ret0[9]), .A2(1'b1), .ZN(
        DP_reg_ret0_n137) );
  OAI21_X1 DP_reg_ret0_U50 ( .B1(1'b1), .B2(DP_reg_ret0_n113), .A(
        DP_reg_ret0_n137), .ZN(DP_reg_ret0_n89) );
  NAND2_X1 DP_reg_ret0_U49 ( .A1(DP_sw0_coeff_ret0[8]), .A2(1'b1), .ZN(
        DP_reg_ret0_n138) );
  OAI21_X1 DP_reg_ret0_U48 ( .B1(1'b1), .B2(DP_reg_ret0_n114), .A(
        DP_reg_ret0_n138), .ZN(DP_reg_ret0_n90) );
  NAND2_X1 DP_reg_ret0_U47 ( .A1(DP_sw0_coeff_ret0[7]), .A2(1'b1), .ZN(
        DP_reg_ret0_n139) );
  OAI21_X1 DP_reg_ret0_U46 ( .B1(1'b1), .B2(DP_reg_ret0_n115), .A(
        DP_reg_ret0_n139), .ZN(DP_reg_ret0_n91) );
  NAND2_X1 DP_reg_ret0_U45 ( .A1(DP_sw0_coeff_ret0[6]), .A2(1'b1), .ZN(
        DP_reg_ret0_n140) );
  OAI21_X1 DP_reg_ret0_U44 ( .B1(1'b1), .B2(DP_reg_ret0_n116), .A(
        DP_reg_ret0_n140), .ZN(DP_reg_ret0_n92) );
  NAND2_X1 DP_reg_ret0_U43 ( .A1(DP_sw0_coeff_ret0[5]), .A2(1'b1), .ZN(
        DP_reg_ret0_n141) );
  OAI21_X1 DP_reg_ret0_U42 ( .B1(1'b1), .B2(DP_reg_ret0_n117), .A(
        DP_reg_ret0_n141), .ZN(DP_reg_ret0_n93) );
  NAND2_X1 DP_reg_ret0_U41 ( .A1(DP_sw0_coeff_ret0[4]), .A2(1'b1), .ZN(
        DP_reg_ret0_n142) );
  OAI21_X1 DP_reg_ret0_U40 ( .B1(1'b1), .B2(DP_reg_ret0_n118), .A(
        DP_reg_ret0_n142), .ZN(DP_reg_ret0_n94) );
  NAND2_X1 DP_reg_ret0_U39 ( .A1(DP_sw0_coeff_ret0[3]), .A2(1'b1), .ZN(
        DP_reg_ret0_n143) );
  OAI21_X1 DP_reg_ret0_U38 ( .B1(1'b1), .B2(DP_reg_ret0_n119), .A(
        DP_reg_ret0_n143), .ZN(DP_reg_ret0_n95) );
  NAND2_X1 DP_reg_ret0_U37 ( .A1(DP_sw0_coeff_ret0[2]), .A2(1'b1), .ZN(
        DP_reg_ret0_n144) );
  OAI21_X1 DP_reg_ret0_U36 ( .B1(1'b1), .B2(DP_reg_ret0_n120), .A(
        DP_reg_ret0_n144), .ZN(DP_reg_ret0_n96) );
  NAND2_X1 DP_reg_ret0_U35 ( .A1(DP_sw0_coeff_ret0[1]), .A2(1'b1), .ZN(
        DP_reg_ret0_n145) );
  OAI21_X1 DP_reg_ret0_U34 ( .B1(1'b1), .B2(DP_reg_ret0_n121), .A(
        DP_reg_ret0_n145), .ZN(DP_reg_ret0_n97) );
  NAND2_X1 DP_reg_ret0_U33 ( .A1(1'b1), .A2(DP_sw0_coeff_ret0[0]), .ZN(
        DP_reg_ret0_n146) );
  OAI21_X1 DP_reg_ret0_U32 ( .B1(1'b1), .B2(DP_reg_ret0_n122), .A(
        DP_reg_ret0_n146), .ZN(DP_reg_ret0_n98) );
  NAND2_X1 DP_reg_ret0_U31 ( .A1(DP_sw0_coeff_ret0[20]), .A2(1'b1), .ZN(
        DP_reg_ret0_n126) );
  OAI21_X1 DP_reg_ret0_U30 ( .B1(1'b1), .B2(DP_reg_ret0_n102), .A(
        DP_reg_ret0_n126), .ZN(DP_reg_ret0_n78) );
  NAND2_X1 DP_reg_ret0_U29 ( .A1(DP_sw0_coeff_ret0[19]), .A2(1'b1), .ZN(
        DP_reg_ret0_n127) );
  OAI21_X1 DP_reg_ret0_U28 ( .B1(1'b1), .B2(DP_reg_ret0_n103), .A(
        DP_reg_ret0_n127), .ZN(DP_reg_ret0_n79) );
  NAND2_X1 DP_reg_ret0_U27 ( .A1(DP_sw0_coeff_ret0[18]), .A2(1'b1), .ZN(
        DP_reg_ret0_n128) );
  OAI21_X1 DP_reg_ret0_U26 ( .B1(1'b1), .B2(DP_reg_ret0_n104), .A(
        DP_reg_ret0_n128), .ZN(DP_reg_ret0_n80) );
  NAND2_X1 DP_reg_ret0_U25 ( .A1(DP_sw0_coeff_ret0[17]), .A2(1'b1), .ZN(
        DP_reg_ret0_n129) );
  OAI21_X1 DP_reg_ret0_U24 ( .B1(1'b1), .B2(DP_reg_ret0_n105), .A(
        DP_reg_ret0_n129), .ZN(DP_reg_ret0_n81) );
  NAND2_X1 DP_reg_ret0_U23 ( .A1(DP_sw0_coeff_ret0[16]), .A2(1'b1), .ZN(
        DP_reg_ret0_n130) );
  OAI21_X1 DP_reg_ret0_U22 ( .B1(1'b1), .B2(DP_reg_ret0_n106), .A(
        DP_reg_ret0_n130), .ZN(DP_reg_ret0_n82) );
  NAND2_X1 DP_reg_ret0_U21 ( .A1(DP_sw0_coeff_ret0[15]), .A2(1'b1), .ZN(
        DP_reg_ret0_n131) );
  OAI21_X1 DP_reg_ret0_U20 ( .B1(1'b1), .B2(DP_reg_ret0_n107), .A(
        DP_reg_ret0_n131), .ZN(DP_reg_ret0_n83) );
  NAND2_X1 DP_reg_ret0_U19 ( .A1(DP_sw0_coeff_ret0[14]), .A2(1'b1), .ZN(
        DP_reg_ret0_n132) );
  OAI21_X1 DP_reg_ret0_U18 ( .B1(1'b1), .B2(DP_reg_ret0_n108), .A(
        DP_reg_ret0_n132), .ZN(DP_reg_ret0_n84) );
  NAND2_X1 DP_reg_ret0_U17 ( .A1(DP_sw0_coeff_ret0[13]), .A2(1'b1), .ZN(
        DP_reg_ret0_n133) );
  OAI21_X1 DP_reg_ret0_U16 ( .B1(1'b1), .B2(DP_reg_ret0_n109), .A(
        DP_reg_ret0_n133), .ZN(DP_reg_ret0_n85) );
  NAND2_X1 DP_reg_ret0_U15 ( .A1(DP_sw0_coeff_ret0[12]), .A2(1'b1), .ZN(
        DP_reg_ret0_n134) );
  OAI21_X1 DP_reg_ret0_U14 ( .B1(1'b1), .B2(DP_reg_ret0_n110), .A(
        DP_reg_ret0_n134), .ZN(DP_reg_ret0_n86) );
  NAND2_X1 DP_reg_ret0_U13 ( .A1(DP_sw0_coeff_ret0[11]), .A2(1'b1), .ZN(
        DP_reg_ret0_n135) );
  OAI21_X1 DP_reg_ret0_U12 ( .B1(1'b1), .B2(DP_reg_ret0_n111), .A(
        DP_reg_ret0_n135), .ZN(DP_reg_ret0_n87) );
  NAND2_X1 DP_reg_ret0_U11 ( .A1(DP_sw0_coeff_ret0[10]), .A2(1'b1), .ZN(
        DP_reg_ret0_n136) );
  OAI21_X1 DP_reg_ret0_U10 ( .B1(1'b1), .B2(DP_reg_ret0_n112), .A(
        DP_reg_ret0_n136), .ZN(DP_reg_ret0_n88) );
  NAND2_X1 DP_reg_ret0_U9 ( .A1(DP_sw0_coeff_ret0[22]), .A2(1'b1), .ZN(
        DP_reg_ret0_n124) );
  OAI21_X1 DP_reg_ret0_U8 ( .B1(1'b1), .B2(DP_reg_ret0_n100), .A(
        DP_reg_ret0_n124), .ZN(DP_reg_ret0_n76) );
  NAND2_X1 DP_reg_ret0_U7 ( .A1(DP_sw0_coeff_ret0[21]), .A2(1'b1), .ZN(
        DP_reg_ret0_n125) );
  OAI21_X1 DP_reg_ret0_U6 ( .B1(1'b1), .B2(DP_reg_ret0_n101), .A(
        DP_reg_ret0_n125), .ZN(DP_reg_ret0_n77) );
  NAND2_X1 DP_reg_ret0_U5 ( .A1(DP_sw0_coeff_ret0[23]), .A2(1'b1), .ZN(
        DP_reg_ret0_n123) );
  OAI21_X1 DP_reg_ret0_U4 ( .B1(1'b1), .B2(DP_reg_ret0_n99), .A(
        DP_reg_ret0_n123), .ZN(DP_reg_ret0_n75) );
  BUF_X1 DP_reg_ret0_U3 ( .A(DP_n6), .Z(DP_reg_ret0_n73) );
  BUF_X1 DP_reg_ret0_U2 ( .A(DP_n6), .Z(DP_reg_ret0_n74) );
  DFFR_X1 DP_reg_ret0_Q_reg_0_ ( .D(DP_reg_ret0_n98), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[0]), .QN(DP_reg_ret0_n122) );
  DFFR_X1 DP_reg_ret0_Q_reg_1_ ( .D(DP_reg_ret0_n97), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[1]), .QN(DP_reg_ret0_n121) );
  DFFR_X1 DP_reg_ret0_Q_reg_2_ ( .D(DP_reg_ret0_n96), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[2]), .QN(DP_reg_ret0_n120) );
  DFFR_X1 DP_reg_ret0_Q_reg_3_ ( .D(DP_reg_ret0_n95), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[3]), .QN(DP_reg_ret0_n119) );
  DFFR_X1 DP_reg_ret0_Q_reg_4_ ( .D(DP_reg_ret0_n94), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[4]), .QN(DP_reg_ret0_n118) );
  DFFR_X1 DP_reg_ret0_Q_reg_5_ ( .D(DP_reg_ret0_n93), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[5]), .QN(DP_reg_ret0_n117) );
  DFFR_X1 DP_reg_ret0_Q_reg_6_ ( .D(DP_reg_ret0_n92), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[6]), .QN(DP_reg_ret0_n116) );
  DFFR_X1 DP_reg_ret0_Q_reg_7_ ( .D(DP_reg_ret0_n91), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[7]), .QN(DP_reg_ret0_n115) );
  DFFR_X1 DP_reg_ret0_Q_reg_8_ ( .D(DP_reg_ret0_n90), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[8]), .QN(DP_reg_ret0_n114) );
  DFFR_X1 DP_reg_ret0_Q_reg_9_ ( .D(DP_reg_ret0_n89), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[9]), .QN(DP_reg_ret0_n113) );
  DFFR_X1 DP_reg_ret0_Q_reg_10_ ( .D(DP_reg_ret0_n88), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[10]), .QN(DP_reg_ret0_n112) );
  DFFR_X1 DP_reg_ret0_Q_reg_11_ ( .D(DP_reg_ret0_n87), .CK(clk), .RN(
        DP_reg_ret0_n74), .Q(DP_ret0[11]), .QN(DP_reg_ret0_n111) );
  DFFR_X1 DP_reg_ret0_Q_reg_12_ ( .D(DP_reg_ret0_n86), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[12]), .QN(DP_reg_ret0_n110) );
  DFFR_X1 DP_reg_ret0_Q_reg_13_ ( .D(DP_reg_ret0_n85), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[13]), .QN(DP_reg_ret0_n109) );
  DFFR_X1 DP_reg_ret0_Q_reg_14_ ( .D(DP_reg_ret0_n84), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[14]), .QN(DP_reg_ret0_n108) );
  DFFR_X1 DP_reg_ret0_Q_reg_15_ ( .D(DP_reg_ret0_n83), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[15]), .QN(DP_reg_ret0_n107) );
  DFFR_X1 DP_reg_ret0_Q_reg_16_ ( .D(DP_reg_ret0_n82), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[16]), .QN(DP_reg_ret0_n106) );
  DFFR_X1 DP_reg_ret0_Q_reg_17_ ( .D(DP_reg_ret0_n81), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[17]), .QN(DP_reg_ret0_n105) );
  DFFR_X1 DP_reg_ret0_Q_reg_18_ ( .D(DP_reg_ret0_n80), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[18]), .QN(DP_reg_ret0_n104) );
  DFFR_X1 DP_reg_ret0_Q_reg_19_ ( .D(DP_reg_ret0_n79), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[19]), .QN(DP_reg_ret0_n103) );
  DFFR_X1 DP_reg_ret0_Q_reg_20_ ( .D(DP_reg_ret0_n78), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[20]), .QN(DP_reg_ret0_n102) );
  DFFR_X1 DP_reg_ret0_Q_reg_21_ ( .D(DP_reg_ret0_n77), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[21]), .QN(DP_reg_ret0_n101) );
  DFFR_X1 DP_reg_ret0_Q_reg_22_ ( .D(DP_reg_ret0_n76), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[22]), .QN(DP_reg_ret0_n100) );
  DFFR_X1 DP_reg_ret0_Q_reg_23_ ( .D(DP_reg_ret0_n75), .CK(clk), .RN(
        DP_reg_ret0_n73), .Q(DP_ret0[23]), .QN(DP_reg_ret0_n99) );
  NAND2_X1 DP_reg_ret1_U51 ( .A1(DP_sw1_coeff_ret1[7]), .A2(1'b1), .ZN(
        DP_reg_ret1_n139) );
  OAI21_X1 DP_reg_ret1_U50 ( .B1(1'b1), .B2(DP_reg_ret1_n115), .A(
        DP_reg_ret1_n139), .ZN(DP_reg_ret1_n91) );
  NAND2_X1 DP_reg_ret1_U49 ( .A1(DP_sw1_coeff_ret1[6]), .A2(1'b1), .ZN(
        DP_reg_ret1_n140) );
  OAI21_X1 DP_reg_ret1_U48 ( .B1(1'b1), .B2(DP_reg_ret1_n116), .A(
        DP_reg_ret1_n140), .ZN(DP_reg_ret1_n92) );
  NAND2_X1 DP_reg_ret1_U47 ( .A1(DP_sw1_coeff_ret1[5]), .A2(1'b1), .ZN(
        DP_reg_ret1_n141) );
  OAI21_X1 DP_reg_ret1_U46 ( .B1(1'b1), .B2(DP_reg_ret1_n117), .A(
        DP_reg_ret1_n141), .ZN(DP_reg_ret1_n93) );
  NAND2_X1 DP_reg_ret1_U45 ( .A1(DP_sw1_coeff_ret1[4]), .A2(1'b1), .ZN(
        DP_reg_ret1_n142) );
  OAI21_X1 DP_reg_ret1_U44 ( .B1(1'b1), .B2(DP_reg_ret1_n118), .A(
        DP_reg_ret1_n142), .ZN(DP_reg_ret1_n94) );
  NAND2_X1 DP_reg_ret1_U43 ( .A1(DP_sw1_coeff_ret1[3]), .A2(1'b1), .ZN(
        DP_reg_ret1_n143) );
  OAI21_X1 DP_reg_ret1_U42 ( .B1(1'b1), .B2(DP_reg_ret1_n119), .A(
        DP_reg_ret1_n143), .ZN(DP_reg_ret1_n95) );
  NAND2_X1 DP_reg_ret1_U41 ( .A1(DP_sw1_coeff_ret1[2]), .A2(1'b1), .ZN(
        DP_reg_ret1_n144) );
  OAI21_X1 DP_reg_ret1_U40 ( .B1(1'b1), .B2(DP_reg_ret1_n120), .A(
        DP_reg_ret1_n144), .ZN(DP_reg_ret1_n96) );
  NAND2_X1 DP_reg_ret1_U39 ( .A1(DP_sw1_coeff_ret1[1]), .A2(1'b1), .ZN(
        DP_reg_ret1_n145) );
  OAI21_X1 DP_reg_ret1_U38 ( .B1(1'b1), .B2(DP_reg_ret1_n121), .A(
        DP_reg_ret1_n145), .ZN(DP_reg_ret1_n97) );
  NAND2_X1 DP_reg_ret1_U37 ( .A1(1'b1), .A2(DP_sw1_coeff_ret1[0]), .ZN(
        DP_reg_ret1_n146) );
  OAI21_X1 DP_reg_ret1_U36 ( .B1(1'b1), .B2(DP_reg_ret1_n122), .A(
        DP_reg_ret1_n146), .ZN(DP_reg_ret1_n98) );
  NAND2_X1 DP_reg_ret1_U35 ( .A1(DP_sw1_coeff_ret1[18]), .A2(1'b1), .ZN(
        DP_reg_ret1_n128) );
  OAI21_X1 DP_reg_ret1_U34 ( .B1(1'b1), .B2(DP_reg_ret1_n104), .A(
        DP_reg_ret1_n128), .ZN(DP_reg_ret1_n80) );
  NAND2_X1 DP_reg_ret1_U33 ( .A1(DP_sw1_coeff_ret1[17]), .A2(1'b1), .ZN(
        DP_reg_ret1_n129) );
  OAI21_X1 DP_reg_ret1_U32 ( .B1(1'b1), .B2(DP_reg_ret1_n105), .A(
        DP_reg_ret1_n129), .ZN(DP_reg_ret1_n81) );
  NAND2_X1 DP_reg_ret1_U31 ( .A1(DP_sw1_coeff_ret1[16]), .A2(1'b1), .ZN(
        DP_reg_ret1_n130) );
  OAI21_X1 DP_reg_ret1_U30 ( .B1(1'b1), .B2(DP_reg_ret1_n106), .A(
        DP_reg_ret1_n130), .ZN(DP_reg_ret1_n82) );
  NAND2_X1 DP_reg_ret1_U29 ( .A1(DP_sw1_coeff_ret1[15]), .A2(1'b1), .ZN(
        DP_reg_ret1_n131) );
  OAI21_X1 DP_reg_ret1_U28 ( .B1(1'b1), .B2(DP_reg_ret1_n107), .A(
        DP_reg_ret1_n131), .ZN(DP_reg_ret1_n83) );
  NAND2_X1 DP_reg_ret1_U27 ( .A1(DP_sw1_coeff_ret1[14]), .A2(1'b1), .ZN(
        DP_reg_ret1_n132) );
  OAI21_X1 DP_reg_ret1_U26 ( .B1(1'b1), .B2(DP_reg_ret1_n108), .A(
        DP_reg_ret1_n132), .ZN(DP_reg_ret1_n84) );
  NAND2_X1 DP_reg_ret1_U25 ( .A1(DP_sw1_coeff_ret1[13]), .A2(1'b1), .ZN(
        DP_reg_ret1_n133) );
  OAI21_X1 DP_reg_ret1_U24 ( .B1(1'b1), .B2(DP_reg_ret1_n109), .A(
        DP_reg_ret1_n133), .ZN(DP_reg_ret1_n85) );
  NAND2_X1 DP_reg_ret1_U23 ( .A1(DP_sw1_coeff_ret1[12]), .A2(1'b1), .ZN(
        DP_reg_ret1_n134) );
  OAI21_X1 DP_reg_ret1_U22 ( .B1(1'b1), .B2(DP_reg_ret1_n110), .A(
        DP_reg_ret1_n134), .ZN(DP_reg_ret1_n86) );
  NAND2_X1 DP_reg_ret1_U21 ( .A1(DP_sw1_coeff_ret1[11]), .A2(1'b1), .ZN(
        DP_reg_ret1_n135) );
  OAI21_X1 DP_reg_ret1_U20 ( .B1(1'b1), .B2(DP_reg_ret1_n111), .A(
        DP_reg_ret1_n135), .ZN(DP_reg_ret1_n87) );
  NAND2_X1 DP_reg_ret1_U19 ( .A1(DP_sw1_coeff_ret1[10]), .A2(1'b1), .ZN(
        DP_reg_ret1_n136) );
  OAI21_X1 DP_reg_ret1_U18 ( .B1(1'b1), .B2(DP_reg_ret1_n112), .A(
        DP_reg_ret1_n136), .ZN(DP_reg_ret1_n88) );
  NAND2_X1 DP_reg_ret1_U17 ( .A1(DP_sw1_coeff_ret1[9]), .A2(1'b1), .ZN(
        DP_reg_ret1_n137) );
  OAI21_X1 DP_reg_ret1_U16 ( .B1(1'b1), .B2(DP_reg_ret1_n113), .A(
        DP_reg_ret1_n137), .ZN(DP_reg_ret1_n89) );
  NAND2_X1 DP_reg_ret1_U15 ( .A1(DP_sw1_coeff_ret1[8]), .A2(1'b1), .ZN(
        DP_reg_ret1_n138) );
  OAI21_X1 DP_reg_ret1_U14 ( .B1(1'b1), .B2(DP_reg_ret1_n114), .A(
        DP_reg_ret1_n138), .ZN(DP_reg_ret1_n90) );
  NAND2_X1 DP_reg_ret1_U13 ( .A1(DP_sw1_coeff_ret1[22]), .A2(1'b1), .ZN(
        DP_reg_ret1_n124) );
  OAI21_X1 DP_reg_ret1_U12 ( .B1(1'b1), .B2(DP_reg_ret1_n100), .A(
        DP_reg_ret1_n124), .ZN(DP_reg_ret1_n76) );
  NAND2_X1 DP_reg_ret1_U11 ( .A1(DP_sw1_coeff_ret1[21]), .A2(1'b1), .ZN(
        DP_reg_ret1_n125) );
  OAI21_X1 DP_reg_ret1_U10 ( .B1(1'b1), .B2(DP_reg_ret1_n101), .A(
        DP_reg_ret1_n125), .ZN(DP_reg_ret1_n77) );
  NAND2_X1 DP_reg_ret1_U9 ( .A1(DP_sw1_coeff_ret1[20]), .A2(1'b1), .ZN(
        DP_reg_ret1_n126) );
  OAI21_X1 DP_reg_ret1_U8 ( .B1(1'b1), .B2(DP_reg_ret1_n102), .A(
        DP_reg_ret1_n126), .ZN(DP_reg_ret1_n78) );
  NAND2_X1 DP_reg_ret1_U7 ( .A1(DP_sw1_coeff_ret1[19]), .A2(1'b1), .ZN(
        DP_reg_ret1_n127) );
  OAI21_X1 DP_reg_ret1_U6 ( .B1(1'b1), .B2(DP_reg_ret1_n103), .A(
        DP_reg_ret1_n127), .ZN(DP_reg_ret1_n79) );
  NAND2_X1 DP_reg_ret1_U5 ( .A1(DP_sw1_coeff_ret1[23]), .A2(1'b1), .ZN(
        DP_reg_ret1_n123) );
  OAI21_X1 DP_reg_ret1_U4 ( .B1(1'b1), .B2(DP_reg_ret1_n99), .A(
        DP_reg_ret1_n123), .ZN(DP_reg_ret1_n75) );
  BUF_X1 DP_reg_ret1_U3 ( .A(DP_n6), .Z(DP_reg_ret1_n73) );
  BUF_X1 DP_reg_ret1_U2 ( .A(DP_n6), .Z(DP_reg_ret1_n74) );
  DFFR_X1 DP_reg_ret1_Q_reg_0_ ( .D(DP_reg_ret1_n98), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[0]), .QN(DP_reg_ret1_n122) );
  DFFR_X1 DP_reg_ret1_Q_reg_1_ ( .D(DP_reg_ret1_n97), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[1]), .QN(DP_reg_ret1_n121) );
  DFFR_X1 DP_reg_ret1_Q_reg_2_ ( .D(DP_reg_ret1_n96), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[2]), .QN(DP_reg_ret1_n120) );
  DFFR_X1 DP_reg_ret1_Q_reg_3_ ( .D(DP_reg_ret1_n95), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[3]), .QN(DP_reg_ret1_n119) );
  DFFR_X1 DP_reg_ret1_Q_reg_4_ ( .D(DP_reg_ret1_n94), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[4]), .QN(DP_reg_ret1_n118) );
  DFFR_X1 DP_reg_ret1_Q_reg_5_ ( .D(DP_reg_ret1_n93), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[5]), .QN(DP_reg_ret1_n117) );
  DFFR_X1 DP_reg_ret1_Q_reg_6_ ( .D(DP_reg_ret1_n92), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[6]), .QN(DP_reg_ret1_n116) );
  DFFR_X1 DP_reg_ret1_Q_reg_7_ ( .D(DP_reg_ret1_n91), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[7]), .QN(DP_reg_ret1_n115) );
  DFFR_X1 DP_reg_ret1_Q_reg_8_ ( .D(DP_reg_ret1_n90), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[8]), .QN(DP_reg_ret1_n114) );
  DFFR_X1 DP_reg_ret1_Q_reg_9_ ( .D(DP_reg_ret1_n89), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[9]), .QN(DP_reg_ret1_n113) );
  DFFR_X1 DP_reg_ret1_Q_reg_10_ ( .D(DP_reg_ret1_n88), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[10]), .QN(DP_reg_ret1_n112) );
  DFFR_X1 DP_reg_ret1_Q_reg_11_ ( .D(DP_reg_ret1_n87), .CK(clk), .RN(
        DP_reg_ret1_n74), .Q(DP_ret1[11]), .QN(DP_reg_ret1_n111) );
  DFFR_X1 DP_reg_ret1_Q_reg_12_ ( .D(DP_reg_ret1_n86), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[12]), .QN(DP_reg_ret1_n110) );
  DFFR_X1 DP_reg_ret1_Q_reg_13_ ( .D(DP_reg_ret1_n85), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[13]), .QN(DP_reg_ret1_n109) );
  DFFR_X1 DP_reg_ret1_Q_reg_14_ ( .D(DP_reg_ret1_n84), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[14]), .QN(DP_reg_ret1_n108) );
  DFFR_X1 DP_reg_ret1_Q_reg_15_ ( .D(DP_reg_ret1_n83), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[15]), .QN(DP_reg_ret1_n107) );
  DFFR_X1 DP_reg_ret1_Q_reg_16_ ( .D(DP_reg_ret1_n82), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[16]), .QN(DP_reg_ret1_n106) );
  DFFR_X1 DP_reg_ret1_Q_reg_17_ ( .D(DP_reg_ret1_n81), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[17]), .QN(DP_reg_ret1_n105) );
  DFFR_X1 DP_reg_ret1_Q_reg_18_ ( .D(DP_reg_ret1_n80), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[18]), .QN(DP_reg_ret1_n104) );
  DFFR_X1 DP_reg_ret1_Q_reg_19_ ( .D(DP_reg_ret1_n79), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[19]), .QN(DP_reg_ret1_n103) );
  DFFR_X1 DP_reg_ret1_Q_reg_20_ ( .D(DP_reg_ret1_n78), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[20]), .QN(DP_reg_ret1_n102) );
  DFFR_X1 DP_reg_ret1_Q_reg_21_ ( .D(DP_reg_ret1_n77), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[21]), .QN(DP_reg_ret1_n101) );
  DFFR_X1 DP_reg_ret1_Q_reg_22_ ( .D(DP_reg_ret1_n76), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[22]), .QN(DP_reg_ret1_n100) );
  DFFR_X1 DP_reg_ret1_Q_reg_23_ ( .D(DP_reg_ret1_n75), .CK(clk), .RN(
        DP_reg_ret1_n73), .Q(DP_ret1[23]), .QN(DP_reg_ret1_n99) );
  NAND2_X1 DP_reg_pipe00_U51 ( .A1(DP_w_6_), .A2(1'b1), .ZN(DP_reg_pipe00_n140) );
  OAI21_X1 DP_reg_pipe00_U50 ( .B1(1'b1), .B2(DP_reg_pipe00_n116), .A(
        DP_reg_pipe00_n140), .ZN(DP_reg_pipe00_n92) );
  NAND2_X1 DP_reg_pipe00_U49 ( .A1(DP_w_5_), .A2(1'b1), .ZN(DP_reg_pipe00_n141) );
  OAI21_X1 DP_reg_pipe00_U48 ( .B1(1'b1), .B2(DP_reg_pipe00_n117), .A(
        DP_reg_pipe00_n141), .ZN(DP_reg_pipe00_n93) );
  NAND2_X1 DP_reg_pipe00_U47 ( .A1(DP_w_4_), .A2(1'b1), .ZN(DP_reg_pipe00_n142) );
  OAI21_X1 DP_reg_pipe00_U46 ( .B1(1'b1), .B2(DP_reg_pipe00_n118), .A(
        DP_reg_pipe00_n142), .ZN(DP_reg_pipe00_n94) );
  NAND2_X1 DP_reg_pipe00_U45 ( .A1(DP_w_3_), .A2(1'b1), .ZN(DP_reg_pipe00_n143) );
  OAI21_X1 DP_reg_pipe00_U44 ( .B1(1'b1), .B2(DP_reg_pipe00_n119), .A(
        DP_reg_pipe00_n143), .ZN(DP_reg_pipe00_n95) );
  NAND2_X1 DP_reg_pipe00_U43 ( .A1(DP_w_2_), .A2(1'b1), .ZN(DP_reg_pipe00_n144) );
  OAI21_X1 DP_reg_pipe00_U42 ( .B1(1'b1), .B2(DP_reg_pipe00_n120), .A(
        DP_reg_pipe00_n144), .ZN(DP_reg_pipe00_n96) );
  NAND2_X1 DP_reg_pipe00_U41 ( .A1(DP_w_1_), .A2(1'b1), .ZN(DP_reg_pipe00_n145) );
  OAI21_X1 DP_reg_pipe00_U40 ( .B1(1'b1), .B2(DP_reg_pipe00_n121), .A(
        DP_reg_pipe00_n145), .ZN(DP_reg_pipe00_n97) );
  NAND2_X1 DP_reg_pipe00_U39 ( .A1(1'b1), .A2(DP_w_0_), .ZN(DP_reg_pipe00_n146) );
  OAI21_X1 DP_reg_pipe00_U38 ( .B1(1'b1), .B2(DP_reg_pipe00_n122), .A(
        DP_reg_pipe00_n146), .ZN(DP_reg_pipe00_n98) );
  NAND2_X1 DP_reg_pipe00_U37 ( .A1(DP_w_14_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n132) );
  OAI21_X1 DP_reg_pipe00_U36 ( .B1(1'b1), .B2(DP_reg_pipe00_n108), .A(
        DP_reg_pipe00_n132), .ZN(DP_reg_pipe00_n84) );
  NAND2_X1 DP_reg_pipe00_U35 ( .A1(DP_w_13_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n133) );
  OAI21_X1 DP_reg_pipe00_U34 ( .B1(1'b1), .B2(DP_reg_pipe00_n109), .A(
        DP_reg_pipe00_n133), .ZN(DP_reg_pipe00_n85) );
  NAND2_X1 DP_reg_pipe00_U33 ( .A1(DP_w_12_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n134) );
  OAI21_X1 DP_reg_pipe00_U32 ( .B1(1'b1), .B2(DP_reg_pipe00_n110), .A(
        DP_reg_pipe00_n134), .ZN(DP_reg_pipe00_n86) );
  NAND2_X1 DP_reg_pipe00_U31 ( .A1(DP_w_11_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n135) );
  OAI21_X1 DP_reg_pipe00_U30 ( .B1(1'b1), .B2(DP_reg_pipe00_n111), .A(
        DP_reg_pipe00_n135), .ZN(DP_reg_pipe00_n87) );
  NAND2_X1 DP_reg_pipe00_U29 ( .A1(DP_w_16_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n130) );
  OAI21_X1 DP_reg_pipe00_U28 ( .B1(1'b1), .B2(DP_reg_pipe00_n106), .A(
        DP_reg_pipe00_n130), .ZN(DP_reg_pipe00_n82) );
  NAND2_X1 DP_reg_pipe00_U27 ( .A1(DP_w_15_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n131) );
  OAI21_X1 DP_reg_pipe00_U26 ( .B1(1'b1), .B2(DP_reg_pipe00_n107), .A(
        DP_reg_pipe00_n131), .ZN(DP_reg_pipe00_n83) );
  NAND2_X1 DP_reg_pipe00_U25 ( .A1(DP_w_10_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n136) );
  OAI21_X1 DP_reg_pipe00_U24 ( .B1(1'b1), .B2(DP_reg_pipe00_n112), .A(
        DP_reg_pipe00_n136), .ZN(DP_reg_pipe00_n88) );
  NAND2_X1 DP_reg_pipe00_U23 ( .A1(DP_w_9_), .A2(1'b1), .ZN(DP_reg_pipe00_n137) );
  OAI21_X1 DP_reg_pipe00_U22 ( .B1(1'b1), .B2(DP_reg_pipe00_n113), .A(
        DP_reg_pipe00_n137), .ZN(DP_reg_pipe00_n89) );
  NAND2_X1 DP_reg_pipe00_U21 ( .A1(DP_w_8_), .A2(1'b1), .ZN(DP_reg_pipe00_n138) );
  OAI21_X1 DP_reg_pipe00_U20 ( .B1(1'b1), .B2(DP_reg_pipe00_n114), .A(
        DP_reg_pipe00_n138), .ZN(DP_reg_pipe00_n90) );
  NAND2_X1 DP_reg_pipe00_U19 ( .A1(DP_w_7_), .A2(1'b1), .ZN(DP_reg_pipe00_n139) );
  OAI21_X1 DP_reg_pipe00_U18 ( .B1(1'b1), .B2(DP_reg_pipe00_n115), .A(
        DP_reg_pipe00_n139), .ZN(DP_reg_pipe00_n91) );
  NAND2_X1 DP_reg_pipe00_U17 ( .A1(DP_w_23_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n123) );
  OAI21_X1 DP_reg_pipe00_U16 ( .B1(1'b1), .B2(DP_reg_pipe00_n99), .A(
        DP_reg_pipe00_n123), .ZN(DP_reg_pipe00_n75) );
  NAND2_X1 DP_reg_pipe00_U15 ( .A1(DP_w_22_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n124) );
  OAI21_X1 DP_reg_pipe00_U14 ( .B1(1'b1), .B2(DP_reg_pipe00_n100), .A(
        DP_reg_pipe00_n124), .ZN(DP_reg_pipe00_n76) );
  NAND2_X1 DP_reg_pipe00_U13 ( .A1(DP_w_20_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n126) );
  OAI21_X1 DP_reg_pipe00_U12 ( .B1(1'b1), .B2(DP_reg_pipe00_n102), .A(
        DP_reg_pipe00_n126), .ZN(DP_reg_pipe00_n78) );
  NAND2_X1 DP_reg_pipe00_U11 ( .A1(DP_w_19_), .A2(1'b1), .ZN(
        DP_reg_pipe00_n127) );
  OAI21_X1 DP_reg_pipe00_U10 ( .B1(1'b1), .B2(DP_reg_pipe00_n103), .A(
        DP_reg_pipe00_n127), .ZN(DP_reg_pipe00_n79) );
  NAND2_X1 DP_reg_pipe00_U9 ( .A1(DP_w_18_), .A2(1'b1), .ZN(DP_reg_pipe00_n128) );
  OAI21_X1 DP_reg_pipe00_U8 ( .B1(1'b1), .B2(DP_reg_pipe00_n104), .A(
        DP_reg_pipe00_n128), .ZN(DP_reg_pipe00_n80) );
  NAND2_X1 DP_reg_pipe00_U7 ( .A1(DP_w_17_), .A2(1'b1), .ZN(DP_reg_pipe00_n129) );
  OAI21_X1 DP_reg_pipe00_U6 ( .B1(1'b1), .B2(DP_reg_pipe00_n105), .A(
        DP_reg_pipe00_n129), .ZN(DP_reg_pipe00_n81) );
  NAND2_X1 DP_reg_pipe00_U5 ( .A1(DP_w_21_), .A2(1'b1), .ZN(DP_reg_pipe00_n125) );
  OAI21_X1 DP_reg_pipe00_U4 ( .B1(1'b1), .B2(DP_reg_pipe00_n101), .A(
        DP_reg_pipe00_n125), .ZN(DP_reg_pipe00_n77) );
  BUF_X1 DP_reg_pipe00_U3 ( .A(DP_n5), .Z(DP_reg_pipe00_n73) );
  BUF_X1 DP_reg_pipe00_U2 ( .A(DP_n5), .Z(DP_reg_pipe00_n74) );
  DFFR_X1 DP_reg_pipe00_Q_reg_0_ ( .D(DP_reg_pipe00_n98), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[0]), .QN(DP_reg_pipe00_n122) );
  DFFR_X1 DP_reg_pipe00_Q_reg_1_ ( .D(DP_reg_pipe00_n97), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[1]), .QN(DP_reg_pipe00_n121) );
  DFFR_X1 DP_reg_pipe00_Q_reg_2_ ( .D(DP_reg_pipe00_n96), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[2]), .QN(DP_reg_pipe00_n120) );
  DFFR_X1 DP_reg_pipe00_Q_reg_3_ ( .D(DP_reg_pipe00_n95), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[3]), .QN(DP_reg_pipe00_n119) );
  DFFR_X1 DP_reg_pipe00_Q_reg_4_ ( .D(DP_reg_pipe00_n94), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[4]), .QN(DP_reg_pipe00_n118) );
  DFFR_X1 DP_reg_pipe00_Q_reg_5_ ( .D(DP_reg_pipe00_n93), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[5]), .QN(DP_reg_pipe00_n117) );
  DFFR_X1 DP_reg_pipe00_Q_reg_6_ ( .D(DP_reg_pipe00_n92), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[6]), .QN(DP_reg_pipe00_n116) );
  DFFR_X1 DP_reg_pipe00_Q_reg_7_ ( .D(DP_reg_pipe00_n91), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[7]), .QN(DP_reg_pipe00_n115) );
  DFFR_X1 DP_reg_pipe00_Q_reg_8_ ( .D(DP_reg_pipe00_n90), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[8]), .QN(DP_reg_pipe00_n114) );
  DFFR_X1 DP_reg_pipe00_Q_reg_9_ ( .D(DP_reg_pipe00_n89), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[9]), .QN(DP_reg_pipe00_n113) );
  DFFR_X1 DP_reg_pipe00_Q_reg_10_ ( .D(DP_reg_pipe00_n88), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[10]), .QN(DP_reg_pipe00_n112) );
  DFFR_X1 DP_reg_pipe00_Q_reg_11_ ( .D(DP_reg_pipe00_n87), .CK(clk), .RN(
        DP_reg_pipe00_n74), .Q(DP_pipe00[11]), .QN(DP_reg_pipe00_n111) );
  DFFR_X1 DP_reg_pipe00_Q_reg_12_ ( .D(DP_reg_pipe00_n86), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[12]), .QN(DP_reg_pipe00_n110) );
  DFFR_X1 DP_reg_pipe00_Q_reg_13_ ( .D(DP_reg_pipe00_n85), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[13]), .QN(DP_reg_pipe00_n109) );
  DFFR_X1 DP_reg_pipe00_Q_reg_14_ ( .D(DP_reg_pipe00_n84), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[14]), .QN(DP_reg_pipe00_n108) );
  DFFR_X1 DP_reg_pipe00_Q_reg_15_ ( .D(DP_reg_pipe00_n83), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[15]), .QN(DP_reg_pipe00_n107) );
  DFFR_X1 DP_reg_pipe00_Q_reg_16_ ( .D(DP_reg_pipe00_n82), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[16]), .QN(DP_reg_pipe00_n106) );
  DFFR_X1 DP_reg_pipe00_Q_reg_17_ ( .D(DP_reg_pipe00_n81), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[17]), .QN(DP_reg_pipe00_n105) );
  DFFR_X1 DP_reg_pipe00_Q_reg_18_ ( .D(DP_reg_pipe00_n80), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[18]), .QN(DP_reg_pipe00_n104) );
  DFFR_X1 DP_reg_pipe00_Q_reg_19_ ( .D(DP_reg_pipe00_n79), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[19]), .QN(DP_reg_pipe00_n103) );
  DFFR_X1 DP_reg_pipe00_Q_reg_20_ ( .D(DP_reg_pipe00_n78), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[20]), .QN(DP_reg_pipe00_n102) );
  DFFR_X1 DP_reg_pipe00_Q_reg_21_ ( .D(DP_reg_pipe00_n77), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[21]), .QN(DP_reg_pipe00_n101) );
  DFFR_X1 DP_reg_pipe00_Q_reg_22_ ( .D(DP_reg_pipe00_n76), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[22]), .QN(DP_reg_pipe00_n100) );
  DFFR_X1 DP_reg_pipe00_Q_reg_23_ ( .D(DP_reg_pipe00_n75), .CK(clk), .RN(
        DP_reg_pipe00_n73), .Q(DP_pipe00[23]), .QN(DP_reg_pipe00_n99) );
  NAND2_X1 DP_reg_pipe01_U51 ( .A1(DP_sw0_23_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n123) );
  OAI21_X1 DP_reg_pipe01_U50 ( .B1(1'b1), .B2(DP_reg_pipe01_n99), .A(
        DP_reg_pipe01_n123), .ZN(DP_reg_pipe01_n75) );
  NAND2_X1 DP_reg_pipe01_U49 ( .A1(DP_sw0_22_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n124) );
  OAI21_X1 DP_reg_pipe01_U48 ( .B1(1'b1), .B2(DP_reg_pipe01_n100), .A(
        DP_reg_pipe01_n124), .ZN(DP_reg_pipe01_n76) );
  NAND2_X1 DP_reg_pipe01_U47 ( .A1(DP_sw0_21_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n125) );
  OAI21_X1 DP_reg_pipe01_U46 ( .B1(1'b1), .B2(DP_reg_pipe01_n101), .A(
        DP_reg_pipe01_n125), .ZN(DP_reg_pipe01_n77) );
  NAND2_X1 DP_reg_pipe01_U45 ( .A1(DP_sw0_20_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n126) );
  OAI21_X1 DP_reg_pipe01_U44 ( .B1(1'b1), .B2(DP_reg_pipe01_n102), .A(
        DP_reg_pipe01_n126), .ZN(DP_reg_pipe01_n78) );
  NAND2_X1 DP_reg_pipe01_U43 ( .A1(DP_sw0_19_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n127) );
  OAI21_X1 DP_reg_pipe01_U42 ( .B1(1'b1), .B2(DP_reg_pipe01_n103), .A(
        DP_reg_pipe01_n127), .ZN(DP_reg_pipe01_n79) );
  NAND2_X1 DP_reg_pipe01_U41 ( .A1(DP_sw0_18_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n128) );
  OAI21_X1 DP_reg_pipe01_U40 ( .B1(1'b1), .B2(DP_reg_pipe01_n104), .A(
        DP_reg_pipe01_n128), .ZN(DP_reg_pipe01_n80) );
  NAND2_X1 DP_reg_pipe01_U39 ( .A1(DP_sw0_17_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n129) );
  OAI21_X1 DP_reg_pipe01_U38 ( .B1(1'b1), .B2(DP_reg_pipe01_n105), .A(
        DP_reg_pipe01_n129), .ZN(DP_reg_pipe01_n81) );
  NAND2_X1 DP_reg_pipe01_U37 ( .A1(DP_sw0_16_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n130) );
  OAI21_X1 DP_reg_pipe01_U36 ( .B1(1'b1), .B2(DP_reg_pipe01_n106), .A(
        DP_reg_pipe01_n130), .ZN(DP_reg_pipe01_n82) );
  NAND2_X1 DP_reg_pipe01_U35 ( .A1(DP_sw0_15_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n131) );
  OAI21_X1 DP_reg_pipe01_U34 ( .B1(1'b1), .B2(DP_reg_pipe01_n107), .A(
        DP_reg_pipe01_n131), .ZN(DP_reg_pipe01_n83) );
  NAND2_X1 DP_reg_pipe01_U33 ( .A1(DP_sw0_14_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n132) );
  OAI21_X1 DP_reg_pipe01_U32 ( .B1(1'b1), .B2(DP_reg_pipe01_n108), .A(
        DP_reg_pipe01_n132), .ZN(DP_reg_pipe01_n84) );
  NAND2_X1 DP_reg_pipe01_U31 ( .A1(DP_sw0_13_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n133) );
  OAI21_X1 DP_reg_pipe01_U30 ( .B1(1'b1), .B2(DP_reg_pipe01_n109), .A(
        DP_reg_pipe01_n133), .ZN(DP_reg_pipe01_n85) );
  NAND2_X1 DP_reg_pipe01_U29 ( .A1(DP_sw0_12_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n134) );
  OAI21_X1 DP_reg_pipe01_U28 ( .B1(1'b1), .B2(DP_reg_pipe01_n110), .A(
        DP_reg_pipe01_n134), .ZN(DP_reg_pipe01_n86) );
  NAND2_X1 DP_reg_pipe01_U27 ( .A1(DP_sw0_11_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n135) );
  OAI21_X1 DP_reg_pipe01_U26 ( .B1(1'b1), .B2(DP_reg_pipe01_n111), .A(
        DP_reg_pipe01_n135), .ZN(DP_reg_pipe01_n87) );
  NAND2_X1 DP_reg_pipe01_U25 ( .A1(DP_sw0_10_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n136) );
  OAI21_X1 DP_reg_pipe01_U24 ( .B1(1'b1), .B2(DP_reg_pipe01_n112), .A(
        DP_reg_pipe01_n136), .ZN(DP_reg_pipe01_n88) );
  NAND2_X1 DP_reg_pipe01_U23 ( .A1(DP_sw0_9_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n137) );
  OAI21_X1 DP_reg_pipe01_U22 ( .B1(1'b1), .B2(DP_reg_pipe01_n113), .A(
        DP_reg_pipe01_n137), .ZN(DP_reg_pipe01_n89) );
  NAND2_X1 DP_reg_pipe01_U21 ( .A1(DP_sw0_8_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n138) );
  OAI21_X1 DP_reg_pipe01_U20 ( .B1(1'b1), .B2(DP_reg_pipe01_n114), .A(
        DP_reg_pipe01_n138), .ZN(DP_reg_pipe01_n90) );
  NAND2_X1 DP_reg_pipe01_U19 ( .A1(DP_sw0_7_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n139) );
  OAI21_X1 DP_reg_pipe01_U18 ( .B1(1'b1), .B2(DP_reg_pipe01_n115), .A(
        DP_reg_pipe01_n139), .ZN(DP_reg_pipe01_n91) );
  NAND2_X1 DP_reg_pipe01_U17 ( .A1(DP_sw0_6_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n140) );
  OAI21_X1 DP_reg_pipe01_U16 ( .B1(1'b1), .B2(DP_reg_pipe01_n116), .A(
        DP_reg_pipe01_n140), .ZN(DP_reg_pipe01_n92) );
  NAND2_X1 DP_reg_pipe01_U15 ( .A1(DP_sw0_5_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n141) );
  OAI21_X1 DP_reg_pipe01_U14 ( .B1(1'b1), .B2(DP_reg_pipe01_n117), .A(
        DP_reg_pipe01_n141), .ZN(DP_reg_pipe01_n93) );
  NAND2_X1 DP_reg_pipe01_U13 ( .A1(DP_sw0_4_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n142) );
  OAI21_X1 DP_reg_pipe01_U12 ( .B1(1'b1), .B2(DP_reg_pipe01_n118), .A(
        DP_reg_pipe01_n142), .ZN(DP_reg_pipe01_n94) );
  NAND2_X1 DP_reg_pipe01_U11 ( .A1(DP_sw0_3_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n143) );
  OAI21_X1 DP_reg_pipe01_U10 ( .B1(1'b1), .B2(DP_reg_pipe01_n119), .A(
        DP_reg_pipe01_n143), .ZN(DP_reg_pipe01_n95) );
  NAND2_X1 DP_reg_pipe01_U9 ( .A1(DP_sw0_2_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n144) );
  OAI21_X1 DP_reg_pipe01_U8 ( .B1(1'b1), .B2(DP_reg_pipe01_n120), .A(
        DP_reg_pipe01_n144), .ZN(DP_reg_pipe01_n96) );
  NAND2_X1 DP_reg_pipe01_U7 ( .A1(DP_sw0_1_), .A2(1'b1), .ZN(
        DP_reg_pipe01_n145) );
  OAI21_X1 DP_reg_pipe01_U6 ( .B1(1'b1), .B2(DP_reg_pipe01_n121), .A(
        DP_reg_pipe01_n145), .ZN(DP_reg_pipe01_n97) );
  NAND2_X1 DP_reg_pipe01_U5 ( .A1(1'b1), .A2(DP_sw0_0_), .ZN(
        DP_reg_pipe01_n146) );
  OAI21_X1 DP_reg_pipe01_U4 ( .B1(1'b1), .B2(DP_reg_pipe01_n122), .A(
        DP_reg_pipe01_n146), .ZN(DP_reg_pipe01_n98) );
  BUF_X1 DP_reg_pipe01_U3 ( .A(DP_n5), .Z(DP_reg_pipe01_n73) );
  BUF_X1 DP_reg_pipe01_U2 ( .A(DP_n5), .Z(DP_reg_pipe01_n74) );
  DFFR_X1 DP_reg_pipe01_Q_reg_0_ ( .D(DP_reg_pipe01_n98), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[0]), .QN(DP_reg_pipe01_n122) );
  DFFR_X1 DP_reg_pipe01_Q_reg_1_ ( .D(DP_reg_pipe01_n97), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[1]), .QN(DP_reg_pipe01_n121) );
  DFFR_X1 DP_reg_pipe01_Q_reg_2_ ( .D(DP_reg_pipe01_n96), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[2]), .QN(DP_reg_pipe01_n120) );
  DFFR_X1 DP_reg_pipe01_Q_reg_3_ ( .D(DP_reg_pipe01_n95), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[3]), .QN(DP_reg_pipe01_n119) );
  DFFR_X1 DP_reg_pipe01_Q_reg_4_ ( .D(DP_reg_pipe01_n94), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[4]), .QN(DP_reg_pipe01_n118) );
  DFFR_X1 DP_reg_pipe01_Q_reg_5_ ( .D(DP_reg_pipe01_n93), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[5]), .QN(DP_reg_pipe01_n117) );
  DFFR_X1 DP_reg_pipe01_Q_reg_6_ ( .D(DP_reg_pipe01_n92), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[6]), .QN(DP_reg_pipe01_n116) );
  DFFR_X1 DP_reg_pipe01_Q_reg_7_ ( .D(DP_reg_pipe01_n91), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[7]), .QN(DP_reg_pipe01_n115) );
  DFFR_X1 DP_reg_pipe01_Q_reg_8_ ( .D(DP_reg_pipe01_n90), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[8]), .QN(DP_reg_pipe01_n114) );
  DFFR_X1 DP_reg_pipe01_Q_reg_9_ ( .D(DP_reg_pipe01_n89), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[9]), .QN(DP_reg_pipe01_n113) );
  DFFR_X1 DP_reg_pipe01_Q_reg_10_ ( .D(DP_reg_pipe01_n88), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[10]), .QN(DP_reg_pipe01_n112) );
  DFFR_X1 DP_reg_pipe01_Q_reg_11_ ( .D(DP_reg_pipe01_n87), .CK(clk), .RN(
        DP_reg_pipe01_n74), .Q(DP_pipe01[11]), .QN(DP_reg_pipe01_n111) );
  DFFR_X1 DP_reg_pipe01_Q_reg_12_ ( .D(DP_reg_pipe01_n86), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[12]), .QN(DP_reg_pipe01_n110) );
  DFFR_X1 DP_reg_pipe01_Q_reg_13_ ( .D(DP_reg_pipe01_n85), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[13]), .QN(DP_reg_pipe01_n109) );
  DFFR_X1 DP_reg_pipe01_Q_reg_14_ ( .D(DP_reg_pipe01_n84), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[14]), .QN(DP_reg_pipe01_n108) );
  DFFR_X1 DP_reg_pipe01_Q_reg_15_ ( .D(DP_reg_pipe01_n83), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[15]), .QN(DP_reg_pipe01_n107) );
  DFFR_X1 DP_reg_pipe01_Q_reg_16_ ( .D(DP_reg_pipe01_n82), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[16]), .QN(DP_reg_pipe01_n106) );
  DFFR_X1 DP_reg_pipe01_Q_reg_17_ ( .D(DP_reg_pipe01_n81), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[17]), .QN(DP_reg_pipe01_n105) );
  DFFR_X1 DP_reg_pipe01_Q_reg_18_ ( .D(DP_reg_pipe01_n80), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[18]), .QN(DP_reg_pipe01_n104) );
  DFFR_X1 DP_reg_pipe01_Q_reg_19_ ( .D(DP_reg_pipe01_n79), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[19]), .QN(DP_reg_pipe01_n103) );
  DFFR_X1 DP_reg_pipe01_Q_reg_20_ ( .D(DP_reg_pipe01_n78), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[20]), .QN(DP_reg_pipe01_n102) );
  DFFR_X1 DP_reg_pipe01_Q_reg_21_ ( .D(DP_reg_pipe01_n77), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[21]), .QN(DP_reg_pipe01_n101) );
  DFFR_X1 DP_reg_pipe01_Q_reg_22_ ( .D(DP_reg_pipe01_n76), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[22]), .QN(DP_reg_pipe01_n100) );
  DFFR_X1 DP_reg_pipe01_Q_reg_23_ ( .D(DP_reg_pipe01_n75), .CK(clk), .RN(
        DP_reg_pipe01_n73), .Q(DP_pipe01[23]), .QN(DP_reg_pipe01_n99) );
  NAND2_X1 DP_reg_pipe02_U51 ( .A1(DP_sw1_23_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n123) );
  OAI21_X1 DP_reg_pipe02_U50 ( .B1(1'b1), .B2(DP_reg_pipe02_n99), .A(
        DP_reg_pipe02_n123), .ZN(DP_reg_pipe02_n75) );
  NAND2_X1 DP_reg_pipe02_U49 ( .A1(DP_sw1_22_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n124) );
  OAI21_X1 DP_reg_pipe02_U48 ( .B1(1'b1), .B2(DP_reg_pipe02_n100), .A(
        DP_reg_pipe02_n124), .ZN(DP_reg_pipe02_n76) );
  NAND2_X1 DP_reg_pipe02_U47 ( .A1(DP_sw1_21_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n125) );
  OAI21_X1 DP_reg_pipe02_U46 ( .B1(1'b1), .B2(DP_reg_pipe02_n101), .A(
        DP_reg_pipe02_n125), .ZN(DP_reg_pipe02_n77) );
  NAND2_X1 DP_reg_pipe02_U45 ( .A1(DP_sw1_20_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n126) );
  OAI21_X1 DP_reg_pipe02_U44 ( .B1(1'b1), .B2(DP_reg_pipe02_n102), .A(
        DP_reg_pipe02_n126), .ZN(DP_reg_pipe02_n78) );
  NAND2_X1 DP_reg_pipe02_U43 ( .A1(DP_sw1_19_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n127) );
  OAI21_X1 DP_reg_pipe02_U42 ( .B1(1'b1), .B2(DP_reg_pipe02_n103), .A(
        DP_reg_pipe02_n127), .ZN(DP_reg_pipe02_n79) );
  NAND2_X1 DP_reg_pipe02_U41 ( .A1(DP_sw1_18_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n128) );
  OAI21_X1 DP_reg_pipe02_U40 ( .B1(1'b1), .B2(DP_reg_pipe02_n104), .A(
        DP_reg_pipe02_n128), .ZN(DP_reg_pipe02_n80) );
  NAND2_X1 DP_reg_pipe02_U39 ( .A1(DP_sw1_17_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n129) );
  OAI21_X1 DP_reg_pipe02_U38 ( .B1(1'b1), .B2(DP_reg_pipe02_n105), .A(
        DP_reg_pipe02_n129), .ZN(DP_reg_pipe02_n81) );
  NAND2_X1 DP_reg_pipe02_U37 ( .A1(DP_sw1_16_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n130) );
  OAI21_X1 DP_reg_pipe02_U36 ( .B1(1'b1), .B2(DP_reg_pipe02_n106), .A(
        DP_reg_pipe02_n130), .ZN(DP_reg_pipe02_n82) );
  NAND2_X1 DP_reg_pipe02_U35 ( .A1(DP_sw1_15_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n131) );
  OAI21_X1 DP_reg_pipe02_U34 ( .B1(1'b1), .B2(DP_reg_pipe02_n107), .A(
        DP_reg_pipe02_n131), .ZN(DP_reg_pipe02_n83) );
  NAND2_X1 DP_reg_pipe02_U33 ( .A1(DP_sw1_14_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n132) );
  OAI21_X1 DP_reg_pipe02_U32 ( .B1(1'b1), .B2(DP_reg_pipe02_n108), .A(
        DP_reg_pipe02_n132), .ZN(DP_reg_pipe02_n84) );
  NAND2_X1 DP_reg_pipe02_U31 ( .A1(DP_sw1_13_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n133) );
  OAI21_X1 DP_reg_pipe02_U30 ( .B1(1'b1), .B2(DP_reg_pipe02_n109), .A(
        DP_reg_pipe02_n133), .ZN(DP_reg_pipe02_n85) );
  NAND2_X1 DP_reg_pipe02_U29 ( .A1(DP_sw1_12_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n134) );
  OAI21_X1 DP_reg_pipe02_U28 ( .B1(1'b1), .B2(DP_reg_pipe02_n110), .A(
        DP_reg_pipe02_n134), .ZN(DP_reg_pipe02_n86) );
  NAND2_X1 DP_reg_pipe02_U27 ( .A1(DP_sw1_11_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n135) );
  OAI21_X1 DP_reg_pipe02_U26 ( .B1(1'b1), .B2(DP_reg_pipe02_n111), .A(
        DP_reg_pipe02_n135), .ZN(DP_reg_pipe02_n87) );
  NAND2_X1 DP_reg_pipe02_U25 ( .A1(DP_sw1_10_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n136) );
  OAI21_X1 DP_reg_pipe02_U24 ( .B1(1'b1), .B2(DP_reg_pipe02_n112), .A(
        DP_reg_pipe02_n136), .ZN(DP_reg_pipe02_n88) );
  NAND2_X1 DP_reg_pipe02_U23 ( .A1(DP_sw1_9_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n137) );
  OAI21_X1 DP_reg_pipe02_U22 ( .B1(1'b1), .B2(DP_reg_pipe02_n113), .A(
        DP_reg_pipe02_n137), .ZN(DP_reg_pipe02_n89) );
  NAND2_X1 DP_reg_pipe02_U21 ( .A1(DP_sw1_8_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n138) );
  OAI21_X1 DP_reg_pipe02_U20 ( .B1(1'b1), .B2(DP_reg_pipe02_n114), .A(
        DP_reg_pipe02_n138), .ZN(DP_reg_pipe02_n90) );
  NAND2_X1 DP_reg_pipe02_U19 ( .A1(DP_sw1_7_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n139) );
  OAI21_X1 DP_reg_pipe02_U18 ( .B1(1'b1), .B2(DP_reg_pipe02_n115), .A(
        DP_reg_pipe02_n139), .ZN(DP_reg_pipe02_n91) );
  NAND2_X1 DP_reg_pipe02_U17 ( .A1(DP_sw1_6_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n140) );
  OAI21_X1 DP_reg_pipe02_U16 ( .B1(1'b1), .B2(DP_reg_pipe02_n116), .A(
        DP_reg_pipe02_n140), .ZN(DP_reg_pipe02_n92) );
  NAND2_X1 DP_reg_pipe02_U15 ( .A1(DP_sw1_5_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n141) );
  OAI21_X1 DP_reg_pipe02_U14 ( .B1(1'b1), .B2(DP_reg_pipe02_n117), .A(
        DP_reg_pipe02_n141), .ZN(DP_reg_pipe02_n93) );
  NAND2_X1 DP_reg_pipe02_U13 ( .A1(DP_sw1_4_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n142) );
  OAI21_X1 DP_reg_pipe02_U12 ( .B1(1'b1), .B2(DP_reg_pipe02_n118), .A(
        DP_reg_pipe02_n142), .ZN(DP_reg_pipe02_n94) );
  NAND2_X1 DP_reg_pipe02_U11 ( .A1(DP_sw1_3_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n143) );
  OAI21_X1 DP_reg_pipe02_U10 ( .B1(1'b1), .B2(DP_reg_pipe02_n119), .A(
        DP_reg_pipe02_n143), .ZN(DP_reg_pipe02_n95) );
  NAND2_X1 DP_reg_pipe02_U9 ( .A1(DP_sw1_2_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n144) );
  OAI21_X1 DP_reg_pipe02_U8 ( .B1(1'b1), .B2(DP_reg_pipe02_n120), .A(
        DP_reg_pipe02_n144), .ZN(DP_reg_pipe02_n96) );
  NAND2_X1 DP_reg_pipe02_U7 ( .A1(DP_sw1_1_), .A2(1'b1), .ZN(
        DP_reg_pipe02_n145) );
  OAI21_X1 DP_reg_pipe02_U6 ( .B1(1'b1), .B2(DP_reg_pipe02_n121), .A(
        DP_reg_pipe02_n145), .ZN(DP_reg_pipe02_n97) );
  NAND2_X1 DP_reg_pipe02_U5 ( .A1(1'b1), .A2(DP_sw1_0_), .ZN(
        DP_reg_pipe02_n146) );
  OAI21_X1 DP_reg_pipe02_U4 ( .B1(1'b1), .B2(DP_reg_pipe02_n122), .A(
        DP_reg_pipe02_n146), .ZN(DP_reg_pipe02_n98) );
  BUF_X1 DP_reg_pipe02_U3 ( .A(DP_n4), .Z(DP_reg_pipe02_n73) );
  BUF_X1 DP_reg_pipe02_U2 ( .A(DP_n4), .Z(DP_reg_pipe02_n74) );
  DFFR_X1 DP_reg_pipe02_Q_reg_0_ ( .D(DP_reg_pipe02_n98), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[0]), .QN(DP_reg_pipe02_n122) );
  DFFR_X1 DP_reg_pipe02_Q_reg_1_ ( .D(DP_reg_pipe02_n97), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[1]), .QN(DP_reg_pipe02_n121) );
  DFFR_X1 DP_reg_pipe02_Q_reg_2_ ( .D(DP_reg_pipe02_n96), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[2]), .QN(DP_reg_pipe02_n120) );
  DFFR_X1 DP_reg_pipe02_Q_reg_3_ ( .D(DP_reg_pipe02_n95), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[3]), .QN(DP_reg_pipe02_n119) );
  DFFR_X1 DP_reg_pipe02_Q_reg_4_ ( .D(DP_reg_pipe02_n94), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[4]), .QN(DP_reg_pipe02_n118) );
  DFFR_X1 DP_reg_pipe02_Q_reg_5_ ( .D(DP_reg_pipe02_n93), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[5]), .QN(DP_reg_pipe02_n117) );
  DFFR_X1 DP_reg_pipe02_Q_reg_6_ ( .D(DP_reg_pipe02_n92), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[6]), .QN(DP_reg_pipe02_n116) );
  DFFR_X1 DP_reg_pipe02_Q_reg_7_ ( .D(DP_reg_pipe02_n91), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[7]), .QN(DP_reg_pipe02_n115) );
  DFFR_X1 DP_reg_pipe02_Q_reg_8_ ( .D(DP_reg_pipe02_n90), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[8]), .QN(DP_reg_pipe02_n114) );
  DFFR_X1 DP_reg_pipe02_Q_reg_9_ ( .D(DP_reg_pipe02_n89), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[9]), .QN(DP_reg_pipe02_n113) );
  DFFR_X1 DP_reg_pipe02_Q_reg_10_ ( .D(DP_reg_pipe02_n88), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[10]), .QN(DP_reg_pipe02_n112) );
  DFFR_X1 DP_reg_pipe02_Q_reg_11_ ( .D(DP_reg_pipe02_n87), .CK(clk), .RN(
        DP_reg_pipe02_n74), .Q(DP_pipe02[11]), .QN(DP_reg_pipe02_n111) );
  DFFR_X1 DP_reg_pipe02_Q_reg_12_ ( .D(DP_reg_pipe02_n86), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[12]), .QN(DP_reg_pipe02_n110) );
  DFFR_X1 DP_reg_pipe02_Q_reg_13_ ( .D(DP_reg_pipe02_n85), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[13]), .QN(DP_reg_pipe02_n109) );
  DFFR_X1 DP_reg_pipe02_Q_reg_14_ ( .D(DP_reg_pipe02_n84), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[14]), .QN(DP_reg_pipe02_n108) );
  DFFR_X1 DP_reg_pipe02_Q_reg_15_ ( .D(DP_reg_pipe02_n83), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[15]), .QN(DP_reg_pipe02_n107) );
  DFFR_X1 DP_reg_pipe02_Q_reg_16_ ( .D(DP_reg_pipe02_n82), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[16]), .QN(DP_reg_pipe02_n106) );
  DFFR_X1 DP_reg_pipe02_Q_reg_17_ ( .D(DP_reg_pipe02_n81), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[17]), .QN(DP_reg_pipe02_n105) );
  DFFR_X1 DP_reg_pipe02_Q_reg_18_ ( .D(DP_reg_pipe02_n80), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[18]), .QN(DP_reg_pipe02_n104) );
  DFFR_X1 DP_reg_pipe02_Q_reg_19_ ( .D(DP_reg_pipe02_n79), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[19]), .QN(DP_reg_pipe02_n103) );
  DFFR_X1 DP_reg_pipe02_Q_reg_20_ ( .D(DP_reg_pipe02_n78), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[20]), .QN(DP_reg_pipe02_n102) );
  DFFR_X1 DP_reg_pipe02_Q_reg_21_ ( .D(DP_reg_pipe02_n77), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[21]), .QN(DP_reg_pipe02_n101) );
  DFFR_X1 DP_reg_pipe02_Q_reg_22_ ( .D(DP_reg_pipe02_n76), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[22]), .QN(DP_reg_pipe02_n100) );
  DFFR_X1 DP_reg_pipe02_Q_reg_23_ ( .D(DP_reg_pipe02_n75), .CK(clk), .RN(
        DP_reg_pipe02_n73), .Q(DP_pipe02[23]), .QN(DP_reg_pipe02_n99) );
  NAND2_X1 DP_reg_pipe03_U51 ( .A1(DP_sw2[23]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n123) );
  OAI21_X1 DP_reg_pipe03_U50 ( .B1(1'b1), .B2(DP_reg_pipe03_n99), .A(
        DP_reg_pipe03_n123), .ZN(DP_reg_pipe03_n75) );
  NAND2_X1 DP_reg_pipe03_U49 ( .A1(DP_sw2[22]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n124) );
  OAI21_X1 DP_reg_pipe03_U48 ( .B1(1'b1), .B2(DP_reg_pipe03_n100), .A(
        DP_reg_pipe03_n124), .ZN(DP_reg_pipe03_n76) );
  NAND2_X1 DP_reg_pipe03_U47 ( .A1(DP_sw2[21]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n125) );
  OAI21_X1 DP_reg_pipe03_U46 ( .B1(1'b1), .B2(DP_reg_pipe03_n101), .A(
        DP_reg_pipe03_n125), .ZN(DP_reg_pipe03_n77) );
  NAND2_X1 DP_reg_pipe03_U45 ( .A1(DP_sw2[20]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n126) );
  OAI21_X1 DP_reg_pipe03_U44 ( .B1(1'b1), .B2(DP_reg_pipe03_n102), .A(
        DP_reg_pipe03_n126), .ZN(DP_reg_pipe03_n78) );
  NAND2_X1 DP_reg_pipe03_U43 ( .A1(DP_sw2[19]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n127) );
  OAI21_X1 DP_reg_pipe03_U42 ( .B1(1'b1), .B2(DP_reg_pipe03_n103), .A(
        DP_reg_pipe03_n127), .ZN(DP_reg_pipe03_n79) );
  NAND2_X1 DP_reg_pipe03_U41 ( .A1(DP_sw2[18]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n128) );
  OAI21_X1 DP_reg_pipe03_U40 ( .B1(1'b1), .B2(DP_reg_pipe03_n104), .A(
        DP_reg_pipe03_n128), .ZN(DP_reg_pipe03_n80) );
  NAND2_X1 DP_reg_pipe03_U39 ( .A1(DP_sw2[17]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n129) );
  OAI21_X1 DP_reg_pipe03_U38 ( .B1(1'b1), .B2(DP_reg_pipe03_n105), .A(
        DP_reg_pipe03_n129), .ZN(DP_reg_pipe03_n81) );
  NAND2_X1 DP_reg_pipe03_U37 ( .A1(DP_sw2[16]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n130) );
  OAI21_X1 DP_reg_pipe03_U36 ( .B1(1'b1), .B2(DP_reg_pipe03_n106), .A(
        DP_reg_pipe03_n130), .ZN(DP_reg_pipe03_n82) );
  NAND2_X1 DP_reg_pipe03_U35 ( .A1(DP_sw2[15]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n131) );
  OAI21_X1 DP_reg_pipe03_U34 ( .B1(1'b1), .B2(DP_reg_pipe03_n107), .A(
        DP_reg_pipe03_n131), .ZN(DP_reg_pipe03_n83) );
  NAND2_X1 DP_reg_pipe03_U33 ( .A1(DP_sw2[14]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n132) );
  OAI21_X1 DP_reg_pipe03_U32 ( .B1(1'b1), .B2(DP_reg_pipe03_n108), .A(
        DP_reg_pipe03_n132), .ZN(DP_reg_pipe03_n84) );
  NAND2_X1 DP_reg_pipe03_U31 ( .A1(DP_sw2[13]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n133) );
  OAI21_X1 DP_reg_pipe03_U30 ( .B1(1'b1), .B2(DP_reg_pipe03_n109), .A(
        DP_reg_pipe03_n133), .ZN(DP_reg_pipe03_n85) );
  NAND2_X1 DP_reg_pipe03_U29 ( .A1(DP_sw2[12]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n134) );
  OAI21_X1 DP_reg_pipe03_U28 ( .B1(1'b1), .B2(DP_reg_pipe03_n110), .A(
        DP_reg_pipe03_n134), .ZN(DP_reg_pipe03_n86) );
  NAND2_X1 DP_reg_pipe03_U27 ( .A1(DP_sw2[11]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n135) );
  OAI21_X1 DP_reg_pipe03_U26 ( .B1(1'b1), .B2(DP_reg_pipe03_n111), .A(
        DP_reg_pipe03_n135), .ZN(DP_reg_pipe03_n87) );
  NAND2_X1 DP_reg_pipe03_U25 ( .A1(DP_sw2[10]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n136) );
  OAI21_X1 DP_reg_pipe03_U24 ( .B1(1'b1), .B2(DP_reg_pipe03_n112), .A(
        DP_reg_pipe03_n136), .ZN(DP_reg_pipe03_n88) );
  NAND2_X1 DP_reg_pipe03_U23 ( .A1(DP_sw2[9]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n137) );
  OAI21_X1 DP_reg_pipe03_U22 ( .B1(1'b1), .B2(DP_reg_pipe03_n113), .A(
        DP_reg_pipe03_n137), .ZN(DP_reg_pipe03_n89) );
  NAND2_X1 DP_reg_pipe03_U21 ( .A1(DP_sw2[8]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n138) );
  OAI21_X1 DP_reg_pipe03_U20 ( .B1(1'b1), .B2(DP_reg_pipe03_n114), .A(
        DP_reg_pipe03_n138), .ZN(DP_reg_pipe03_n90) );
  NAND2_X1 DP_reg_pipe03_U19 ( .A1(DP_sw2[7]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n139) );
  OAI21_X1 DP_reg_pipe03_U18 ( .B1(1'b1), .B2(DP_reg_pipe03_n115), .A(
        DP_reg_pipe03_n139), .ZN(DP_reg_pipe03_n91) );
  NAND2_X1 DP_reg_pipe03_U17 ( .A1(DP_sw2[6]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n140) );
  OAI21_X1 DP_reg_pipe03_U16 ( .B1(1'b1), .B2(DP_reg_pipe03_n116), .A(
        DP_reg_pipe03_n140), .ZN(DP_reg_pipe03_n92) );
  NAND2_X1 DP_reg_pipe03_U15 ( .A1(DP_sw2[5]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n141) );
  OAI21_X1 DP_reg_pipe03_U14 ( .B1(1'b1), .B2(DP_reg_pipe03_n117), .A(
        DP_reg_pipe03_n141), .ZN(DP_reg_pipe03_n93) );
  NAND2_X1 DP_reg_pipe03_U13 ( .A1(DP_sw2[4]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n142) );
  OAI21_X1 DP_reg_pipe03_U12 ( .B1(1'b1), .B2(DP_reg_pipe03_n118), .A(
        DP_reg_pipe03_n142), .ZN(DP_reg_pipe03_n94) );
  NAND2_X1 DP_reg_pipe03_U11 ( .A1(DP_sw2[3]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n143) );
  OAI21_X1 DP_reg_pipe03_U10 ( .B1(1'b1), .B2(DP_reg_pipe03_n119), .A(
        DP_reg_pipe03_n143), .ZN(DP_reg_pipe03_n95) );
  NAND2_X1 DP_reg_pipe03_U9 ( .A1(DP_sw2[2]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n144) );
  OAI21_X1 DP_reg_pipe03_U8 ( .B1(1'b1), .B2(DP_reg_pipe03_n120), .A(
        DP_reg_pipe03_n144), .ZN(DP_reg_pipe03_n96) );
  NAND2_X1 DP_reg_pipe03_U7 ( .A1(DP_sw2[1]), .A2(1'b1), .ZN(
        DP_reg_pipe03_n145) );
  OAI21_X1 DP_reg_pipe03_U6 ( .B1(1'b1), .B2(DP_reg_pipe03_n121), .A(
        DP_reg_pipe03_n145), .ZN(DP_reg_pipe03_n97) );
  NAND2_X1 DP_reg_pipe03_U5 ( .A1(1'b1), .A2(DP_sw2[0]), .ZN(
        DP_reg_pipe03_n146) );
  OAI21_X1 DP_reg_pipe03_U4 ( .B1(1'b1), .B2(DP_reg_pipe03_n122), .A(
        DP_reg_pipe03_n146), .ZN(DP_reg_pipe03_n98) );
  BUF_X1 DP_reg_pipe03_U3 ( .A(DP_n3), .Z(DP_reg_pipe03_n73) );
  BUF_X1 DP_reg_pipe03_U2 ( .A(DP_n3), .Z(DP_reg_pipe03_n74) );
  DFFR_X1 DP_reg_pipe03_Q_reg_0_ ( .D(DP_reg_pipe03_n98), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[0]), .QN(DP_reg_pipe03_n122) );
  DFFR_X1 DP_reg_pipe03_Q_reg_1_ ( .D(DP_reg_pipe03_n97), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[1]), .QN(DP_reg_pipe03_n121) );
  DFFR_X1 DP_reg_pipe03_Q_reg_2_ ( .D(DP_reg_pipe03_n96), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[2]), .QN(DP_reg_pipe03_n120) );
  DFFR_X1 DP_reg_pipe03_Q_reg_3_ ( .D(DP_reg_pipe03_n95), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[3]), .QN(DP_reg_pipe03_n119) );
  DFFR_X1 DP_reg_pipe03_Q_reg_4_ ( .D(DP_reg_pipe03_n94), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[4]), .QN(DP_reg_pipe03_n118) );
  DFFR_X1 DP_reg_pipe03_Q_reg_5_ ( .D(DP_reg_pipe03_n93), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[5]), .QN(DP_reg_pipe03_n117) );
  DFFR_X1 DP_reg_pipe03_Q_reg_6_ ( .D(DP_reg_pipe03_n92), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[6]), .QN(DP_reg_pipe03_n116) );
  DFFR_X1 DP_reg_pipe03_Q_reg_7_ ( .D(DP_reg_pipe03_n91), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[7]), .QN(DP_reg_pipe03_n115) );
  DFFR_X1 DP_reg_pipe03_Q_reg_8_ ( .D(DP_reg_pipe03_n90), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[8]), .QN(DP_reg_pipe03_n114) );
  DFFR_X1 DP_reg_pipe03_Q_reg_9_ ( .D(DP_reg_pipe03_n89), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[9]), .QN(DP_reg_pipe03_n113) );
  DFFR_X1 DP_reg_pipe03_Q_reg_10_ ( .D(DP_reg_pipe03_n88), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[10]), .QN(DP_reg_pipe03_n112) );
  DFFR_X1 DP_reg_pipe03_Q_reg_11_ ( .D(DP_reg_pipe03_n87), .CK(clk), .RN(
        DP_reg_pipe03_n74), .Q(DP_pipe03[11]), .QN(DP_reg_pipe03_n111) );
  DFFR_X1 DP_reg_pipe03_Q_reg_12_ ( .D(DP_reg_pipe03_n86), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[12]), .QN(DP_reg_pipe03_n110) );
  DFFR_X1 DP_reg_pipe03_Q_reg_13_ ( .D(DP_reg_pipe03_n85), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[13]), .QN(DP_reg_pipe03_n109) );
  DFFR_X1 DP_reg_pipe03_Q_reg_14_ ( .D(DP_reg_pipe03_n84), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[14]), .QN(DP_reg_pipe03_n108) );
  DFFR_X1 DP_reg_pipe03_Q_reg_15_ ( .D(DP_reg_pipe03_n83), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[15]), .QN(DP_reg_pipe03_n107) );
  DFFR_X1 DP_reg_pipe03_Q_reg_16_ ( .D(DP_reg_pipe03_n82), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[16]), .QN(DP_reg_pipe03_n106) );
  DFFR_X1 DP_reg_pipe03_Q_reg_17_ ( .D(DP_reg_pipe03_n81), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[17]), .QN(DP_reg_pipe03_n105) );
  DFFR_X1 DP_reg_pipe03_Q_reg_18_ ( .D(DP_reg_pipe03_n80), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[18]), .QN(DP_reg_pipe03_n104) );
  DFFR_X1 DP_reg_pipe03_Q_reg_19_ ( .D(DP_reg_pipe03_n79), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[19]), .QN(DP_reg_pipe03_n103) );
  DFFR_X1 DP_reg_pipe03_Q_reg_20_ ( .D(DP_reg_pipe03_n78), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[20]), .QN(DP_reg_pipe03_n102) );
  DFFR_X1 DP_reg_pipe03_Q_reg_21_ ( .D(DP_reg_pipe03_n77), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[21]), .QN(DP_reg_pipe03_n101) );
  DFFR_X1 DP_reg_pipe03_Q_reg_22_ ( .D(DP_reg_pipe03_n76), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[22]), .QN(DP_reg_pipe03_n100) );
  DFFR_X1 DP_reg_pipe03_Q_reg_23_ ( .D(DP_reg_pipe03_n75), .CK(clk), .RN(
        DP_reg_pipe03_n73), .Q(DP_pipe03[23]), .QN(DP_reg_pipe03_n99) );
  NAND2_X1 DP_reg_pipe10_U51 ( .A1(DP_pipe0_b0[1]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n145) );
  OAI21_X1 DP_reg_pipe10_U50 ( .B1(1'b1), .B2(DP_reg_pipe10_n121), .A(
        DP_reg_pipe10_n145), .ZN(DP_reg_pipe10_n97) );
  NAND2_X1 DP_reg_pipe10_U49 ( .A1(1'b1), .A2(DP_pipe0_b0[0]), .ZN(
        DP_reg_pipe10_n146) );
  OAI21_X1 DP_reg_pipe10_U48 ( .B1(1'b1), .B2(DP_reg_pipe10_n122), .A(
        DP_reg_pipe10_n146), .ZN(DP_reg_pipe10_n98) );
  NAND2_X1 DP_reg_pipe10_U47 ( .A1(DP_pipe0_b0[12]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n134) );
  OAI21_X1 DP_reg_pipe10_U46 ( .B1(1'b1), .B2(DP_reg_pipe10_n110), .A(
        DP_reg_pipe10_n134), .ZN(DP_reg_pipe10_n86) );
  NAND2_X1 DP_reg_pipe10_U45 ( .A1(DP_pipe0_b0[11]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n135) );
  OAI21_X1 DP_reg_pipe10_U44 ( .B1(1'b1), .B2(DP_reg_pipe10_n111), .A(
        DP_reg_pipe10_n135), .ZN(DP_reg_pipe10_n87) );
  NAND2_X1 DP_reg_pipe10_U43 ( .A1(DP_pipe0_b0[10]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n136) );
  OAI21_X1 DP_reg_pipe10_U42 ( .B1(1'b1), .B2(DP_reg_pipe10_n112), .A(
        DP_reg_pipe10_n136), .ZN(DP_reg_pipe10_n88) );
  NAND2_X1 DP_reg_pipe10_U41 ( .A1(DP_pipe0_b0[9]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n137) );
  OAI21_X1 DP_reg_pipe10_U40 ( .B1(1'b1), .B2(DP_reg_pipe10_n113), .A(
        DP_reg_pipe10_n137), .ZN(DP_reg_pipe10_n89) );
  NAND2_X1 DP_reg_pipe10_U39 ( .A1(DP_pipe0_b0[8]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n138) );
  OAI21_X1 DP_reg_pipe10_U38 ( .B1(1'b1), .B2(DP_reg_pipe10_n114), .A(
        DP_reg_pipe10_n138), .ZN(DP_reg_pipe10_n90) );
  NAND2_X1 DP_reg_pipe10_U37 ( .A1(DP_pipe0_b0[7]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n139) );
  OAI21_X1 DP_reg_pipe10_U36 ( .B1(1'b1), .B2(DP_reg_pipe10_n115), .A(
        DP_reg_pipe10_n139), .ZN(DP_reg_pipe10_n91) );
  NAND2_X1 DP_reg_pipe10_U35 ( .A1(DP_pipe0_b0[6]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n140) );
  OAI21_X1 DP_reg_pipe10_U34 ( .B1(1'b1), .B2(DP_reg_pipe10_n116), .A(
        DP_reg_pipe10_n140), .ZN(DP_reg_pipe10_n92) );
  NAND2_X1 DP_reg_pipe10_U33 ( .A1(DP_pipe0_b0[5]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n141) );
  OAI21_X1 DP_reg_pipe10_U32 ( .B1(1'b1), .B2(DP_reg_pipe10_n117), .A(
        DP_reg_pipe10_n141), .ZN(DP_reg_pipe10_n93) );
  NAND2_X1 DP_reg_pipe10_U31 ( .A1(DP_pipe0_b0[4]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n142) );
  OAI21_X1 DP_reg_pipe10_U30 ( .B1(1'b1), .B2(DP_reg_pipe10_n118), .A(
        DP_reg_pipe10_n142), .ZN(DP_reg_pipe10_n94) );
  NAND2_X1 DP_reg_pipe10_U29 ( .A1(DP_pipe0_b0[3]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n143) );
  OAI21_X1 DP_reg_pipe10_U28 ( .B1(1'b1), .B2(DP_reg_pipe10_n119), .A(
        DP_reg_pipe10_n143), .ZN(DP_reg_pipe10_n95) );
  NAND2_X1 DP_reg_pipe10_U27 ( .A1(DP_pipe0_b0[2]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n144) );
  OAI21_X1 DP_reg_pipe10_U26 ( .B1(1'b1), .B2(DP_reg_pipe10_n120), .A(
        DP_reg_pipe10_n144), .ZN(DP_reg_pipe10_n96) );
  NAND2_X1 DP_reg_pipe10_U25 ( .A1(DP_pipe0_b0[22]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n124) );
  OAI21_X1 DP_reg_pipe10_U24 ( .B1(1'b1), .B2(DP_reg_pipe10_n100), .A(
        DP_reg_pipe10_n124), .ZN(DP_reg_pipe10_n76) );
  NAND2_X1 DP_reg_pipe10_U23 ( .A1(DP_pipe0_b0[19]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n127) );
  OAI21_X1 DP_reg_pipe10_U22 ( .B1(1'b1), .B2(DP_reg_pipe10_n103), .A(
        DP_reg_pipe10_n127), .ZN(DP_reg_pipe10_n79) );
  NAND2_X1 DP_reg_pipe10_U21 ( .A1(DP_pipe0_b0[18]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n128) );
  OAI21_X1 DP_reg_pipe10_U20 ( .B1(1'b1), .B2(DP_reg_pipe10_n104), .A(
        DP_reg_pipe10_n128), .ZN(DP_reg_pipe10_n80) );
  NAND2_X1 DP_reg_pipe10_U19 ( .A1(DP_pipe0_b0[15]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n131) );
  OAI21_X1 DP_reg_pipe10_U18 ( .B1(1'b1), .B2(DP_reg_pipe10_n107), .A(
        DP_reg_pipe10_n131), .ZN(DP_reg_pipe10_n83) );
  NAND2_X1 DP_reg_pipe10_U17 ( .A1(DP_pipe0_b0[14]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n132) );
  OAI21_X1 DP_reg_pipe10_U16 ( .B1(1'b1), .B2(DP_reg_pipe10_n108), .A(
        DP_reg_pipe10_n132), .ZN(DP_reg_pipe10_n84) );
  NAND2_X1 DP_reg_pipe10_U15 ( .A1(DP_pipe0_b0[13]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n133) );
  OAI21_X1 DP_reg_pipe10_U14 ( .B1(1'b1), .B2(DP_reg_pipe10_n109), .A(
        DP_reg_pipe10_n133), .ZN(DP_reg_pipe10_n85) );
  NAND2_X1 DP_reg_pipe10_U13 ( .A1(DP_pipe0_b0[21]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n125) );
  OAI21_X1 DP_reg_pipe10_U12 ( .B1(1'b1), .B2(DP_reg_pipe10_n101), .A(
        DP_reg_pipe10_n125), .ZN(DP_reg_pipe10_n77) );
  NAND2_X1 DP_reg_pipe10_U11 ( .A1(DP_pipe0_b0[20]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n126) );
  OAI21_X1 DP_reg_pipe10_U10 ( .B1(1'b1), .B2(DP_reg_pipe10_n102), .A(
        DP_reg_pipe10_n126), .ZN(DP_reg_pipe10_n78) );
  NAND2_X1 DP_reg_pipe10_U9 ( .A1(DP_pipe0_b0[17]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n129) );
  OAI21_X1 DP_reg_pipe10_U8 ( .B1(1'b1), .B2(DP_reg_pipe10_n105), .A(
        DP_reg_pipe10_n129), .ZN(DP_reg_pipe10_n81) );
  NAND2_X1 DP_reg_pipe10_U7 ( .A1(DP_pipe0_b0[16]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n130) );
  OAI21_X1 DP_reg_pipe10_U6 ( .B1(1'b1), .B2(DP_reg_pipe10_n106), .A(
        DP_reg_pipe10_n130), .ZN(DP_reg_pipe10_n82) );
  NAND2_X1 DP_reg_pipe10_U5 ( .A1(DP_pipe0_b0[23]), .A2(1'b1), .ZN(
        DP_reg_pipe10_n123) );
  OAI21_X1 DP_reg_pipe10_U4 ( .B1(1'b1), .B2(DP_reg_pipe10_n99), .A(
        DP_reg_pipe10_n123), .ZN(DP_reg_pipe10_n75) );
  BUF_X1 DP_reg_pipe10_U3 ( .A(DP_n3), .Z(DP_reg_pipe10_n73) );
  BUF_X1 DP_reg_pipe10_U2 ( .A(DP_n3), .Z(DP_reg_pipe10_n74) );
  DFFR_X1 DP_reg_pipe10_Q_reg_0_ ( .D(DP_reg_pipe10_n98), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[0]), .QN(DP_reg_pipe10_n122) );
  DFFR_X1 DP_reg_pipe10_Q_reg_1_ ( .D(DP_reg_pipe10_n97), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[1]), .QN(DP_reg_pipe10_n121) );
  DFFR_X1 DP_reg_pipe10_Q_reg_2_ ( .D(DP_reg_pipe10_n96), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[2]), .QN(DP_reg_pipe10_n120) );
  DFFR_X1 DP_reg_pipe10_Q_reg_3_ ( .D(DP_reg_pipe10_n95), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[3]), .QN(DP_reg_pipe10_n119) );
  DFFR_X1 DP_reg_pipe10_Q_reg_4_ ( .D(DP_reg_pipe10_n94), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[4]), .QN(DP_reg_pipe10_n118) );
  DFFR_X1 DP_reg_pipe10_Q_reg_5_ ( .D(DP_reg_pipe10_n93), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[5]), .QN(DP_reg_pipe10_n117) );
  DFFR_X1 DP_reg_pipe10_Q_reg_6_ ( .D(DP_reg_pipe10_n92), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[6]), .QN(DP_reg_pipe10_n116) );
  DFFR_X1 DP_reg_pipe10_Q_reg_7_ ( .D(DP_reg_pipe10_n91), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[7]), .QN(DP_reg_pipe10_n115) );
  DFFR_X1 DP_reg_pipe10_Q_reg_8_ ( .D(DP_reg_pipe10_n90), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[8]), .QN(DP_reg_pipe10_n114) );
  DFFR_X1 DP_reg_pipe10_Q_reg_9_ ( .D(DP_reg_pipe10_n89), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[9]), .QN(DP_reg_pipe10_n113) );
  DFFR_X1 DP_reg_pipe10_Q_reg_10_ ( .D(DP_reg_pipe10_n88), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[10]), .QN(DP_reg_pipe10_n112) );
  DFFR_X1 DP_reg_pipe10_Q_reg_11_ ( .D(DP_reg_pipe10_n87), .CK(clk), .RN(
        DP_reg_pipe10_n74), .Q(DP_pipe10[11]), .QN(DP_reg_pipe10_n111) );
  DFFR_X1 DP_reg_pipe10_Q_reg_12_ ( .D(DP_reg_pipe10_n86), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[12]), .QN(DP_reg_pipe10_n110) );
  DFFR_X1 DP_reg_pipe10_Q_reg_13_ ( .D(DP_reg_pipe10_n85), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[13]), .QN(DP_reg_pipe10_n109) );
  DFFR_X1 DP_reg_pipe10_Q_reg_14_ ( .D(DP_reg_pipe10_n84), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[14]), .QN(DP_reg_pipe10_n108) );
  DFFR_X1 DP_reg_pipe10_Q_reg_15_ ( .D(DP_reg_pipe10_n83), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[15]), .QN(DP_reg_pipe10_n107) );
  DFFR_X1 DP_reg_pipe10_Q_reg_16_ ( .D(DP_reg_pipe10_n82), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[16]), .QN(DP_reg_pipe10_n106) );
  DFFR_X1 DP_reg_pipe10_Q_reg_17_ ( .D(DP_reg_pipe10_n81), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[17]), .QN(DP_reg_pipe10_n105) );
  DFFR_X1 DP_reg_pipe10_Q_reg_18_ ( .D(DP_reg_pipe10_n80), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[18]), .QN(DP_reg_pipe10_n104) );
  DFFR_X1 DP_reg_pipe10_Q_reg_19_ ( .D(DP_reg_pipe10_n79), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[19]), .QN(DP_reg_pipe10_n103) );
  DFFR_X1 DP_reg_pipe10_Q_reg_20_ ( .D(DP_reg_pipe10_n78), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[20]), .QN(DP_reg_pipe10_n102) );
  DFFR_X1 DP_reg_pipe10_Q_reg_21_ ( .D(DP_reg_pipe10_n77), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[21]), .QN(DP_reg_pipe10_n101) );
  DFFR_X1 DP_reg_pipe10_Q_reg_22_ ( .D(DP_reg_pipe10_n76), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[22]), .QN(DP_reg_pipe10_n100) );
  DFFR_X1 DP_reg_pipe10_Q_reg_23_ ( .D(DP_reg_pipe10_n75), .CK(clk), .RN(
        DP_reg_pipe10_n73), .Q(DP_pipe10[23]), .QN(DP_reg_pipe10_n99) );
  NAND2_X1 DP_reg_pipe11_U51 ( .A1(DP_pipe0_coeff_pipe01[6]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n140) );
  OAI21_X1 DP_reg_pipe11_U50 ( .B1(1'b1), .B2(DP_reg_pipe11_n116), .A(
        DP_reg_pipe11_n140), .ZN(DP_reg_pipe11_n92) );
  NAND2_X1 DP_reg_pipe11_U49 ( .A1(DP_pipe0_coeff_pipe01[5]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n141) );
  OAI21_X1 DP_reg_pipe11_U48 ( .B1(1'b1), .B2(DP_reg_pipe11_n117), .A(
        DP_reg_pipe11_n141), .ZN(DP_reg_pipe11_n93) );
  NAND2_X1 DP_reg_pipe11_U47 ( .A1(DP_pipe0_coeff_pipe01[4]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n142) );
  OAI21_X1 DP_reg_pipe11_U46 ( .B1(1'b1), .B2(DP_reg_pipe11_n118), .A(
        DP_reg_pipe11_n142), .ZN(DP_reg_pipe11_n94) );
  NAND2_X1 DP_reg_pipe11_U45 ( .A1(DP_pipe0_coeff_pipe01[3]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n143) );
  OAI21_X1 DP_reg_pipe11_U44 ( .B1(1'b1), .B2(DP_reg_pipe11_n119), .A(
        DP_reg_pipe11_n143), .ZN(DP_reg_pipe11_n95) );
  NAND2_X1 DP_reg_pipe11_U43 ( .A1(DP_pipe0_coeff_pipe01[2]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n144) );
  OAI21_X1 DP_reg_pipe11_U42 ( .B1(1'b1), .B2(DP_reg_pipe11_n120), .A(
        DP_reg_pipe11_n144), .ZN(DP_reg_pipe11_n96) );
  NAND2_X1 DP_reg_pipe11_U41 ( .A1(DP_pipe0_coeff_pipe01[1]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n145) );
  OAI21_X1 DP_reg_pipe11_U40 ( .B1(1'b1), .B2(DP_reg_pipe11_n121), .A(
        DP_reg_pipe11_n145), .ZN(DP_reg_pipe11_n97) );
  NAND2_X1 DP_reg_pipe11_U39 ( .A1(1'b1), .A2(DP_pipe0_coeff_pipe01[0]), .ZN(
        DP_reg_pipe11_n146) );
  OAI21_X1 DP_reg_pipe11_U38 ( .B1(1'b1), .B2(DP_reg_pipe11_n122), .A(
        DP_reg_pipe11_n146), .ZN(DP_reg_pipe11_n98) );
  NAND2_X1 DP_reg_pipe11_U37 ( .A1(DP_pipe0_coeff_pipe01[17]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n129) );
  OAI21_X1 DP_reg_pipe11_U36 ( .B1(1'b1), .B2(DP_reg_pipe11_n105), .A(
        DP_reg_pipe11_n129), .ZN(DP_reg_pipe11_n81) );
  NAND2_X1 DP_reg_pipe11_U35 ( .A1(DP_pipe0_coeff_pipe01[16]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n130) );
  OAI21_X1 DP_reg_pipe11_U34 ( .B1(1'b1), .B2(DP_reg_pipe11_n106), .A(
        DP_reg_pipe11_n130), .ZN(DP_reg_pipe11_n82) );
  NAND2_X1 DP_reg_pipe11_U33 ( .A1(DP_pipe0_coeff_pipe01[15]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n131) );
  OAI21_X1 DP_reg_pipe11_U32 ( .B1(1'b1), .B2(DP_reg_pipe11_n107), .A(
        DP_reg_pipe11_n131), .ZN(DP_reg_pipe11_n83) );
  NAND2_X1 DP_reg_pipe11_U31 ( .A1(DP_pipe0_coeff_pipe01[14]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n132) );
  OAI21_X1 DP_reg_pipe11_U30 ( .B1(1'b1), .B2(DP_reg_pipe11_n108), .A(
        DP_reg_pipe11_n132), .ZN(DP_reg_pipe11_n84) );
  NAND2_X1 DP_reg_pipe11_U29 ( .A1(DP_pipe0_coeff_pipe01[13]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n133) );
  OAI21_X1 DP_reg_pipe11_U28 ( .B1(1'b1), .B2(DP_reg_pipe11_n109), .A(
        DP_reg_pipe11_n133), .ZN(DP_reg_pipe11_n85) );
  NAND2_X1 DP_reg_pipe11_U27 ( .A1(DP_pipe0_coeff_pipe01[12]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n134) );
  OAI21_X1 DP_reg_pipe11_U26 ( .B1(1'b1), .B2(DP_reg_pipe11_n110), .A(
        DP_reg_pipe11_n134), .ZN(DP_reg_pipe11_n86) );
  NAND2_X1 DP_reg_pipe11_U25 ( .A1(DP_pipe0_coeff_pipe01[11]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n135) );
  OAI21_X1 DP_reg_pipe11_U24 ( .B1(1'b1), .B2(DP_reg_pipe11_n111), .A(
        DP_reg_pipe11_n135), .ZN(DP_reg_pipe11_n87) );
  NAND2_X1 DP_reg_pipe11_U23 ( .A1(DP_pipe0_coeff_pipe01[10]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n136) );
  OAI21_X1 DP_reg_pipe11_U22 ( .B1(1'b1), .B2(DP_reg_pipe11_n112), .A(
        DP_reg_pipe11_n136), .ZN(DP_reg_pipe11_n88) );
  NAND2_X1 DP_reg_pipe11_U21 ( .A1(DP_pipe0_coeff_pipe01[9]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n137) );
  OAI21_X1 DP_reg_pipe11_U20 ( .B1(1'b1), .B2(DP_reg_pipe11_n113), .A(
        DP_reg_pipe11_n137), .ZN(DP_reg_pipe11_n89) );
  NAND2_X1 DP_reg_pipe11_U19 ( .A1(DP_pipe0_coeff_pipe01[8]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n138) );
  OAI21_X1 DP_reg_pipe11_U18 ( .B1(1'b1), .B2(DP_reg_pipe11_n114), .A(
        DP_reg_pipe11_n138), .ZN(DP_reg_pipe11_n90) );
  NAND2_X1 DP_reg_pipe11_U17 ( .A1(DP_pipe0_coeff_pipe01[7]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n139) );
  OAI21_X1 DP_reg_pipe11_U16 ( .B1(1'b1), .B2(DP_reg_pipe11_n115), .A(
        DP_reg_pipe11_n139), .ZN(DP_reg_pipe11_n91) );
  NAND2_X1 DP_reg_pipe11_U15 ( .A1(DP_pipe0_coeff_pipe01[22]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n124) );
  OAI21_X1 DP_reg_pipe11_U14 ( .B1(1'b1), .B2(DP_reg_pipe11_n100), .A(
        DP_reg_pipe11_n124), .ZN(DP_reg_pipe11_n76) );
  NAND2_X1 DP_reg_pipe11_U13 ( .A1(DP_pipe0_coeff_pipe01[21]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n125) );
  OAI21_X1 DP_reg_pipe11_U12 ( .B1(1'b1), .B2(DP_reg_pipe11_n101), .A(
        DP_reg_pipe11_n125), .ZN(DP_reg_pipe11_n77) );
  NAND2_X1 DP_reg_pipe11_U11 ( .A1(DP_pipe0_coeff_pipe01[20]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n126) );
  OAI21_X1 DP_reg_pipe11_U10 ( .B1(1'b1), .B2(DP_reg_pipe11_n102), .A(
        DP_reg_pipe11_n126), .ZN(DP_reg_pipe11_n78) );
  NAND2_X1 DP_reg_pipe11_U9 ( .A1(DP_pipe0_coeff_pipe01[19]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n127) );
  OAI21_X1 DP_reg_pipe11_U8 ( .B1(1'b1), .B2(DP_reg_pipe11_n103), .A(
        DP_reg_pipe11_n127), .ZN(DP_reg_pipe11_n79) );
  NAND2_X1 DP_reg_pipe11_U7 ( .A1(DP_pipe0_coeff_pipe01[18]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n128) );
  OAI21_X1 DP_reg_pipe11_U6 ( .B1(1'b1), .B2(DP_reg_pipe11_n104), .A(
        DP_reg_pipe11_n128), .ZN(DP_reg_pipe11_n80) );
  NAND2_X1 DP_reg_pipe11_U5 ( .A1(DP_pipe0_coeff_pipe01[23]), .A2(1'b1), .ZN(
        DP_reg_pipe11_n123) );
  OAI21_X1 DP_reg_pipe11_U4 ( .B1(1'b1), .B2(DP_reg_pipe11_n99), .A(
        DP_reg_pipe11_n123), .ZN(DP_reg_pipe11_n75) );
  BUF_X1 DP_reg_pipe11_U3 ( .A(DP_n2), .Z(DP_reg_pipe11_n73) );
  BUF_X1 DP_reg_pipe11_U2 ( .A(DP_n2), .Z(DP_reg_pipe11_n74) );
  DFFR_X1 DP_reg_pipe11_Q_reg_0_ ( .D(DP_reg_pipe11_n98), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[0]), .QN(DP_reg_pipe11_n122) );
  DFFR_X1 DP_reg_pipe11_Q_reg_1_ ( .D(DP_reg_pipe11_n97), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[1]), .QN(DP_reg_pipe11_n121) );
  DFFR_X1 DP_reg_pipe11_Q_reg_2_ ( .D(DP_reg_pipe11_n96), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[2]), .QN(DP_reg_pipe11_n120) );
  DFFR_X1 DP_reg_pipe11_Q_reg_3_ ( .D(DP_reg_pipe11_n95), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[3]), .QN(DP_reg_pipe11_n119) );
  DFFR_X1 DP_reg_pipe11_Q_reg_4_ ( .D(DP_reg_pipe11_n94), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[4]), .QN(DP_reg_pipe11_n118) );
  DFFR_X1 DP_reg_pipe11_Q_reg_5_ ( .D(DP_reg_pipe11_n93), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[5]), .QN(DP_reg_pipe11_n117) );
  DFFR_X1 DP_reg_pipe11_Q_reg_6_ ( .D(DP_reg_pipe11_n92), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[6]), .QN(DP_reg_pipe11_n116) );
  DFFR_X1 DP_reg_pipe11_Q_reg_7_ ( .D(DP_reg_pipe11_n91), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[7]), .QN(DP_reg_pipe11_n115) );
  DFFR_X1 DP_reg_pipe11_Q_reg_8_ ( .D(DP_reg_pipe11_n90), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[8]), .QN(DP_reg_pipe11_n114) );
  DFFR_X1 DP_reg_pipe11_Q_reg_9_ ( .D(DP_reg_pipe11_n89), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[9]), .QN(DP_reg_pipe11_n113) );
  DFFR_X1 DP_reg_pipe11_Q_reg_10_ ( .D(DP_reg_pipe11_n88), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[10]), .QN(DP_reg_pipe11_n112) );
  DFFR_X1 DP_reg_pipe11_Q_reg_11_ ( .D(DP_reg_pipe11_n87), .CK(clk), .RN(
        DP_reg_pipe11_n74), .Q(DP_pipe11[11]), .QN(DP_reg_pipe11_n111) );
  DFFR_X1 DP_reg_pipe11_Q_reg_12_ ( .D(DP_reg_pipe11_n86), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[12]), .QN(DP_reg_pipe11_n110) );
  DFFR_X1 DP_reg_pipe11_Q_reg_13_ ( .D(DP_reg_pipe11_n85), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[13]), .QN(DP_reg_pipe11_n109) );
  DFFR_X1 DP_reg_pipe11_Q_reg_14_ ( .D(DP_reg_pipe11_n84), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[14]), .QN(DP_reg_pipe11_n108) );
  DFFR_X1 DP_reg_pipe11_Q_reg_15_ ( .D(DP_reg_pipe11_n83), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[15]), .QN(DP_reg_pipe11_n107) );
  DFFR_X1 DP_reg_pipe11_Q_reg_16_ ( .D(DP_reg_pipe11_n82), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[16]), .QN(DP_reg_pipe11_n106) );
  DFFR_X1 DP_reg_pipe11_Q_reg_17_ ( .D(DP_reg_pipe11_n81), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[17]), .QN(DP_reg_pipe11_n105) );
  DFFR_X1 DP_reg_pipe11_Q_reg_18_ ( .D(DP_reg_pipe11_n80), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[18]), .QN(DP_reg_pipe11_n104) );
  DFFR_X1 DP_reg_pipe11_Q_reg_19_ ( .D(DP_reg_pipe11_n79), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[19]), .QN(DP_reg_pipe11_n103) );
  DFFR_X1 DP_reg_pipe11_Q_reg_20_ ( .D(DP_reg_pipe11_n78), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[20]), .QN(DP_reg_pipe11_n102) );
  DFFR_X1 DP_reg_pipe11_Q_reg_21_ ( .D(DP_reg_pipe11_n77), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[21]), .QN(DP_reg_pipe11_n101) );
  DFFR_X1 DP_reg_pipe11_Q_reg_22_ ( .D(DP_reg_pipe11_n76), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[22]), .QN(DP_reg_pipe11_n100) );
  DFFR_X1 DP_reg_pipe11_Q_reg_23_ ( .D(DP_reg_pipe11_n75), .CK(clk), .RN(
        DP_reg_pipe11_n73), .Q(DP_pipe11[23]), .QN(DP_reg_pipe11_n99) );
  NAND2_X1 DP_reg_pipe12_U51 ( .A1(DP_pipe0_coeff_pipe02[6]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n140) );
  OAI21_X1 DP_reg_pipe12_U50 ( .B1(1'b1), .B2(DP_reg_pipe12_n116), .A(
        DP_reg_pipe12_n140), .ZN(DP_reg_pipe12_n92) );
  NAND2_X1 DP_reg_pipe12_U49 ( .A1(DP_pipe0_coeff_pipe02[5]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n141) );
  OAI21_X1 DP_reg_pipe12_U48 ( .B1(1'b1), .B2(DP_reg_pipe12_n117), .A(
        DP_reg_pipe12_n141), .ZN(DP_reg_pipe12_n93) );
  NAND2_X1 DP_reg_pipe12_U47 ( .A1(DP_pipe0_coeff_pipe02[4]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n142) );
  OAI21_X1 DP_reg_pipe12_U46 ( .B1(1'b1), .B2(DP_reg_pipe12_n118), .A(
        DP_reg_pipe12_n142), .ZN(DP_reg_pipe12_n94) );
  NAND2_X1 DP_reg_pipe12_U45 ( .A1(DP_pipe0_coeff_pipe02[3]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n143) );
  OAI21_X1 DP_reg_pipe12_U44 ( .B1(1'b1), .B2(DP_reg_pipe12_n119), .A(
        DP_reg_pipe12_n143), .ZN(DP_reg_pipe12_n95) );
  NAND2_X1 DP_reg_pipe12_U43 ( .A1(DP_pipe0_coeff_pipe02[2]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n144) );
  OAI21_X1 DP_reg_pipe12_U42 ( .B1(1'b1), .B2(DP_reg_pipe12_n120), .A(
        DP_reg_pipe12_n144), .ZN(DP_reg_pipe12_n96) );
  NAND2_X1 DP_reg_pipe12_U41 ( .A1(DP_pipe0_coeff_pipe02[1]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n145) );
  OAI21_X1 DP_reg_pipe12_U40 ( .B1(1'b1), .B2(DP_reg_pipe12_n121), .A(
        DP_reg_pipe12_n145), .ZN(DP_reg_pipe12_n97) );
  NAND2_X1 DP_reg_pipe12_U39 ( .A1(1'b1), .A2(DP_pipe0_coeff_pipe02[0]), .ZN(
        DP_reg_pipe12_n146) );
  OAI21_X1 DP_reg_pipe12_U38 ( .B1(1'b1), .B2(DP_reg_pipe12_n122), .A(
        DP_reg_pipe12_n146), .ZN(DP_reg_pipe12_n98) );
  NAND2_X1 DP_reg_pipe12_U37 ( .A1(DP_pipe0_coeff_pipe02[17]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n129) );
  OAI21_X1 DP_reg_pipe12_U36 ( .B1(1'b1), .B2(DP_reg_pipe12_n105), .A(
        DP_reg_pipe12_n129), .ZN(DP_reg_pipe12_n81) );
  NAND2_X1 DP_reg_pipe12_U35 ( .A1(DP_pipe0_coeff_pipe02[16]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n130) );
  OAI21_X1 DP_reg_pipe12_U34 ( .B1(1'b1), .B2(DP_reg_pipe12_n106), .A(
        DP_reg_pipe12_n130), .ZN(DP_reg_pipe12_n82) );
  NAND2_X1 DP_reg_pipe12_U33 ( .A1(DP_pipe0_coeff_pipe02[15]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n131) );
  OAI21_X1 DP_reg_pipe12_U32 ( .B1(1'b1), .B2(DP_reg_pipe12_n107), .A(
        DP_reg_pipe12_n131), .ZN(DP_reg_pipe12_n83) );
  NAND2_X1 DP_reg_pipe12_U31 ( .A1(DP_pipe0_coeff_pipe02[14]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n132) );
  OAI21_X1 DP_reg_pipe12_U30 ( .B1(1'b1), .B2(DP_reg_pipe12_n108), .A(
        DP_reg_pipe12_n132), .ZN(DP_reg_pipe12_n84) );
  NAND2_X1 DP_reg_pipe12_U29 ( .A1(DP_pipe0_coeff_pipe02[13]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n133) );
  OAI21_X1 DP_reg_pipe12_U28 ( .B1(1'b1), .B2(DP_reg_pipe12_n109), .A(
        DP_reg_pipe12_n133), .ZN(DP_reg_pipe12_n85) );
  NAND2_X1 DP_reg_pipe12_U27 ( .A1(DP_pipe0_coeff_pipe02[12]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n134) );
  OAI21_X1 DP_reg_pipe12_U26 ( .B1(1'b1), .B2(DP_reg_pipe12_n110), .A(
        DP_reg_pipe12_n134), .ZN(DP_reg_pipe12_n86) );
  NAND2_X1 DP_reg_pipe12_U25 ( .A1(DP_pipe0_coeff_pipe02[11]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n135) );
  OAI21_X1 DP_reg_pipe12_U24 ( .B1(1'b1), .B2(DP_reg_pipe12_n111), .A(
        DP_reg_pipe12_n135), .ZN(DP_reg_pipe12_n87) );
  NAND2_X1 DP_reg_pipe12_U23 ( .A1(DP_pipe0_coeff_pipe02[10]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n136) );
  OAI21_X1 DP_reg_pipe12_U22 ( .B1(1'b1), .B2(DP_reg_pipe12_n112), .A(
        DP_reg_pipe12_n136), .ZN(DP_reg_pipe12_n88) );
  NAND2_X1 DP_reg_pipe12_U21 ( .A1(DP_pipe0_coeff_pipe02[9]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n137) );
  OAI21_X1 DP_reg_pipe12_U20 ( .B1(1'b1), .B2(DP_reg_pipe12_n113), .A(
        DP_reg_pipe12_n137), .ZN(DP_reg_pipe12_n89) );
  NAND2_X1 DP_reg_pipe12_U19 ( .A1(DP_pipe0_coeff_pipe02[8]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n138) );
  OAI21_X1 DP_reg_pipe12_U18 ( .B1(1'b1), .B2(DP_reg_pipe12_n114), .A(
        DP_reg_pipe12_n138), .ZN(DP_reg_pipe12_n90) );
  NAND2_X1 DP_reg_pipe12_U17 ( .A1(DP_pipe0_coeff_pipe02[7]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n139) );
  OAI21_X1 DP_reg_pipe12_U16 ( .B1(1'b1), .B2(DP_reg_pipe12_n115), .A(
        DP_reg_pipe12_n139), .ZN(DP_reg_pipe12_n91) );
  NAND2_X1 DP_reg_pipe12_U15 ( .A1(DP_pipe0_coeff_pipe02[22]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n124) );
  OAI21_X1 DP_reg_pipe12_U14 ( .B1(1'b1), .B2(DP_reg_pipe12_n100), .A(
        DP_reg_pipe12_n124), .ZN(DP_reg_pipe12_n76) );
  NAND2_X1 DP_reg_pipe12_U13 ( .A1(DP_pipe0_coeff_pipe02[21]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n125) );
  OAI21_X1 DP_reg_pipe12_U12 ( .B1(1'b1), .B2(DP_reg_pipe12_n101), .A(
        DP_reg_pipe12_n125), .ZN(DP_reg_pipe12_n77) );
  NAND2_X1 DP_reg_pipe12_U11 ( .A1(DP_pipe0_coeff_pipe02[20]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n126) );
  OAI21_X1 DP_reg_pipe12_U10 ( .B1(1'b1), .B2(DP_reg_pipe12_n102), .A(
        DP_reg_pipe12_n126), .ZN(DP_reg_pipe12_n78) );
  NAND2_X1 DP_reg_pipe12_U9 ( .A1(DP_pipe0_coeff_pipe02[19]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n127) );
  OAI21_X1 DP_reg_pipe12_U8 ( .B1(1'b1), .B2(DP_reg_pipe12_n103), .A(
        DP_reg_pipe12_n127), .ZN(DP_reg_pipe12_n79) );
  NAND2_X1 DP_reg_pipe12_U7 ( .A1(DP_pipe0_coeff_pipe02[18]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n128) );
  OAI21_X1 DP_reg_pipe12_U6 ( .B1(1'b1), .B2(DP_reg_pipe12_n104), .A(
        DP_reg_pipe12_n128), .ZN(DP_reg_pipe12_n80) );
  NAND2_X1 DP_reg_pipe12_U5 ( .A1(DP_pipe0_coeff_pipe02[23]), .A2(1'b1), .ZN(
        DP_reg_pipe12_n123) );
  OAI21_X1 DP_reg_pipe12_U4 ( .B1(1'b1), .B2(DP_reg_pipe12_n99), .A(
        DP_reg_pipe12_n123), .ZN(DP_reg_pipe12_n75) );
  BUF_X1 DP_reg_pipe12_U3 ( .A(DP_n2), .Z(DP_reg_pipe12_n73) );
  BUF_X1 DP_reg_pipe12_U2 ( .A(DP_n2), .Z(DP_reg_pipe12_n74) );
  DFFR_X1 DP_reg_pipe12_Q_reg_0_ ( .D(DP_reg_pipe12_n98), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[0]), .QN(DP_reg_pipe12_n122) );
  DFFR_X1 DP_reg_pipe12_Q_reg_1_ ( .D(DP_reg_pipe12_n97), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[1]), .QN(DP_reg_pipe12_n121) );
  DFFR_X1 DP_reg_pipe12_Q_reg_2_ ( .D(DP_reg_pipe12_n96), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[2]), .QN(DP_reg_pipe12_n120) );
  DFFR_X1 DP_reg_pipe12_Q_reg_3_ ( .D(DP_reg_pipe12_n95), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[3]), .QN(DP_reg_pipe12_n119) );
  DFFR_X1 DP_reg_pipe12_Q_reg_4_ ( .D(DP_reg_pipe12_n94), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[4]), .QN(DP_reg_pipe12_n118) );
  DFFR_X1 DP_reg_pipe12_Q_reg_5_ ( .D(DP_reg_pipe12_n93), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[5]), .QN(DP_reg_pipe12_n117) );
  DFFR_X1 DP_reg_pipe12_Q_reg_6_ ( .D(DP_reg_pipe12_n92), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[6]), .QN(DP_reg_pipe12_n116) );
  DFFR_X1 DP_reg_pipe12_Q_reg_7_ ( .D(DP_reg_pipe12_n91), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[7]), .QN(DP_reg_pipe12_n115) );
  DFFR_X1 DP_reg_pipe12_Q_reg_8_ ( .D(DP_reg_pipe12_n90), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[8]), .QN(DP_reg_pipe12_n114) );
  DFFR_X1 DP_reg_pipe12_Q_reg_9_ ( .D(DP_reg_pipe12_n89), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[9]), .QN(DP_reg_pipe12_n113) );
  DFFR_X1 DP_reg_pipe12_Q_reg_10_ ( .D(DP_reg_pipe12_n88), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[10]), .QN(DP_reg_pipe12_n112) );
  DFFR_X1 DP_reg_pipe12_Q_reg_11_ ( .D(DP_reg_pipe12_n87), .CK(clk), .RN(
        DP_reg_pipe12_n74), .Q(DP_pipe12[11]), .QN(DP_reg_pipe12_n111) );
  DFFR_X1 DP_reg_pipe12_Q_reg_12_ ( .D(DP_reg_pipe12_n86), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[12]), .QN(DP_reg_pipe12_n110) );
  DFFR_X1 DP_reg_pipe12_Q_reg_13_ ( .D(DP_reg_pipe12_n85), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[13]), .QN(DP_reg_pipe12_n109) );
  DFFR_X1 DP_reg_pipe12_Q_reg_14_ ( .D(DP_reg_pipe12_n84), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[14]), .QN(DP_reg_pipe12_n108) );
  DFFR_X1 DP_reg_pipe12_Q_reg_15_ ( .D(DP_reg_pipe12_n83), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[15]), .QN(DP_reg_pipe12_n107) );
  DFFR_X1 DP_reg_pipe12_Q_reg_16_ ( .D(DP_reg_pipe12_n82), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[16]), .QN(DP_reg_pipe12_n106) );
  DFFR_X1 DP_reg_pipe12_Q_reg_17_ ( .D(DP_reg_pipe12_n81), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[17]), .QN(DP_reg_pipe12_n105) );
  DFFR_X1 DP_reg_pipe12_Q_reg_18_ ( .D(DP_reg_pipe12_n80), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[18]), .QN(DP_reg_pipe12_n104) );
  DFFR_X1 DP_reg_pipe12_Q_reg_19_ ( .D(DP_reg_pipe12_n79), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[19]), .QN(DP_reg_pipe12_n103) );
  DFFR_X1 DP_reg_pipe12_Q_reg_20_ ( .D(DP_reg_pipe12_n78), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[20]), .QN(DP_reg_pipe12_n102) );
  DFFR_X1 DP_reg_pipe12_Q_reg_21_ ( .D(DP_reg_pipe12_n77), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[21]), .QN(DP_reg_pipe12_n101) );
  DFFR_X1 DP_reg_pipe12_Q_reg_22_ ( .D(DP_reg_pipe12_n76), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[22]), .QN(DP_reg_pipe12_n100) );
  DFFR_X1 DP_reg_pipe12_Q_reg_23_ ( .D(DP_reg_pipe12_n75), .CK(clk), .RN(
        DP_reg_pipe12_n73), .Q(DP_pipe12[23]), .QN(DP_reg_pipe12_n99) );
  NAND2_X1 DP_reg_pipe13_U51 ( .A1(DP_pipe0_coeff_pipe03[7]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n139) );
  OAI21_X1 DP_reg_pipe13_U50 ( .B1(1'b1), .B2(DP_reg_pipe13_n115), .A(
        DP_reg_pipe13_n139), .ZN(DP_reg_pipe13_n91) );
  NAND2_X1 DP_reg_pipe13_U49 ( .A1(DP_pipe0_coeff_pipe03[6]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n140) );
  OAI21_X1 DP_reg_pipe13_U48 ( .B1(1'b1), .B2(DP_reg_pipe13_n116), .A(
        DP_reg_pipe13_n140), .ZN(DP_reg_pipe13_n92) );
  NAND2_X1 DP_reg_pipe13_U47 ( .A1(DP_pipe0_coeff_pipe03[5]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n141) );
  OAI21_X1 DP_reg_pipe13_U46 ( .B1(1'b1), .B2(DP_reg_pipe13_n117), .A(
        DP_reg_pipe13_n141), .ZN(DP_reg_pipe13_n93) );
  NAND2_X1 DP_reg_pipe13_U45 ( .A1(DP_pipe0_coeff_pipe03[4]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n142) );
  OAI21_X1 DP_reg_pipe13_U44 ( .B1(1'b1), .B2(DP_reg_pipe13_n118), .A(
        DP_reg_pipe13_n142), .ZN(DP_reg_pipe13_n94) );
  NAND2_X1 DP_reg_pipe13_U43 ( .A1(DP_pipe0_coeff_pipe03[3]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n143) );
  OAI21_X1 DP_reg_pipe13_U42 ( .B1(1'b1), .B2(DP_reg_pipe13_n119), .A(
        DP_reg_pipe13_n143), .ZN(DP_reg_pipe13_n95) );
  NAND2_X1 DP_reg_pipe13_U41 ( .A1(DP_pipe0_coeff_pipe03[2]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n144) );
  OAI21_X1 DP_reg_pipe13_U40 ( .B1(1'b1), .B2(DP_reg_pipe13_n120), .A(
        DP_reg_pipe13_n144), .ZN(DP_reg_pipe13_n96) );
  NAND2_X1 DP_reg_pipe13_U39 ( .A1(DP_pipe0_coeff_pipe03[1]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n145) );
  OAI21_X1 DP_reg_pipe13_U38 ( .B1(1'b1), .B2(DP_reg_pipe13_n121), .A(
        DP_reg_pipe13_n145), .ZN(DP_reg_pipe13_n97) );
  NAND2_X1 DP_reg_pipe13_U37 ( .A1(1'b1), .A2(DP_pipe0_coeff_pipe03[0]), .ZN(
        DP_reg_pipe13_n146) );
  OAI21_X1 DP_reg_pipe13_U36 ( .B1(1'b1), .B2(DP_reg_pipe13_n122), .A(
        DP_reg_pipe13_n146), .ZN(DP_reg_pipe13_n98) );
  NAND2_X1 DP_reg_pipe13_U35 ( .A1(DP_pipe0_coeff_pipe03[18]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n128) );
  OAI21_X1 DP_reg_pipe13_U34 ( .B1(1'b1), .B2(DP_reg_pipe13_n104), .A(
        DP_reg_pipe13_n128), .ZN(DP_reg_pipe13_n80) );
  NAND2_X1 DP_reg_pipe13_U33 ( .A1(DP_pipe0_coeff_pipe03[17]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n129) );
  OAI21_X1 DP_reg_pipe13_U32 ( .B1(1'b1), .B2(DP_reg_pipe13_n105), .A(
        DP_reg_pipe13_n129), .ZN(DP_reg_pipe13_n81) );
  NAND2_X1 DP_reg_pipe13_U31 ( .A1(DP_pipe0_coeff_pipe03[16]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n130) );
  OAI21_X1 DP_reg_pipe13_U30 ( .B1(1'b1), .B2(DP_reg_pipe13_n106), .A(
        DP_reg_pipe13_n130), .ZN(DP_reg_pipe13_n82) );
  NAND2_X1 DP_reg_pipe13_U29 ( .A1(DP_pipe0_coeff_pipe03[15]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n131) );
  OAI21_X1 DP_reg_pipe13_U28 ( .B1(1'b1), .B2(DP_reg_pipe13_n107), .A(
        DP_reg_pipe13_n131), .ZN(DP_reg_pipe13_n83) );
  NAND2_X1 DP_reg_pipe13_U27 ( .A1(DP_pipe0_coeff_pipe03[14]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n132) );
  OAI21_X1 DP_reg_pipe13_U26 ( .B1(1'b1), .B2(DP_reg_pipe13_n108), .A(
        DP_reg_pipe13_n132), .ZN(DP_reg_pipe13_n84) );
  NAND2_X1 DP_reg_pipe13_U25 ( .A1(DP_pipe0_coeff_pipe03[13]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n133) );
  OAI21_X1 DP_reg_pipe13_U24 ( .B1(1'b1), .B2(DP_reg_pipe13_n109), .A(
        DP_reg_pipe13_n133), .ZN(DP_reg_pipe13_n85) );
  NAND2_X1 DP_reg_pipe13_U23 ( .A1(DP_pipe0_coeff_pipe03[12]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n134) );
  OAI21_X1 DP_reg_pipe13_U22 ( .B1(1'b1), .B2(DP_reg_pipe13_n110), .A(
        DP_reg_pipe13_n134), .ZN(DP_reg_pipe13_n86) );
  NAND2_X1 DP_reg_pipe13_U21 ( .A1(DP_pipe0_coeff_pipe03[11]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n135) );
  OAI21_X1 DP_reg_pipe13_U20 ( .B1(1'b1), .B2(DP_reg_pipe13_n111), .A(
        DP_reg_pipe13_n135), .ZN(DP_reg_pipe13_n87) );
  NAND2_X1 DP_reg_pipe13_U19 ( .A1(DP_pipe0_coeff_pipe03[10]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n136) );
  OAI21_X1 DP_reg_pipe13_U18 ( .B1(1'b1), .B2(DP_reg_pipe13_n112), .A(
        DP_reg_pipe13_n136), .ZN(DP_reg_pipe13_n88) );
  NAND2_X1 DP_reg_pipe13_U17 ( .A1(DP_pipe0_coeff_pipe03[9]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n137) );
  OAI21_X1 DP_reg_pipe13_U16 ( .B1(1'b1), .B2(DP_reg_pipe13_n113), .A(
        DP_reg_pipe13_n137), .ZN(DP_reg_pipe13_n89) );
  NAND2_X1 DP_reg_pipe13_U15 ( .A1(DP_pipe0_coeff_pipe03[8]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n138) );
  OAI21_X1 DP_reg_pipe13_U14 ( .B1(1'b1), .B2(DP_reg_pipe13_n114), .A(
        DP_reg_pipe13_n138), .ZN(DP_reg_pipe13_n90) );
  NAND2_X1 DP_reg_pipe13_U13 ( .A1(DP_pipe0_coeff_pipe03[22]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n124) );
  OAI21_X1 DP_reg_pipe13_U12 ( .B1(1'b1), .B2(DP_reg_pipe13_n100), .A(
        DP_reg_pipe13_n124), .ZN(DP_reg_pipe13_n76) );
  NAND2_X1 DP_reg_pipe13_U11 ( .A1(DP_pipe0_coeff_pipe03[21]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n125) );
  OAI21_X1 DP_reg_pipe13_U10 ( .B1(1'b1), .B2(DP_reg_pipe13_n101), .A(
        DP_reg_pipe13_n125), .ZN(DP_reg_pipe13_n77) );
  NAND2_X1 DP_reg_pipe13_U9 ( .A1(DP_pipe0_coeff_pipe03[20]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n126) );
  OAI21_X1 DP_reg_pipe13_U8 ( .B1(1'b1), .B2(DP_reg_pipe13_n102), .A(
        DP_reg_pipe13_n126), .ZN(DP_reg_pipe13_n78) );
  NAND2_X1 DP_reg_pipe13_U7 ( .A1(DP_pipe0_coeff_pipe03[19]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n127) );
  OAI21_X1 DP_reg_pipe13_U6 ( .B1(1'b1), .B2(DP_reg_pipe13_n103), .A(
        DP_reg_pipe13_n127), .ZN(DP_reg_pipe13_n79) );
  NAND2_X1 DP_reg_pipe13_U5 ( .A1(DP_pipe0_coeff_pipe03[23]), .A2(1'b1), .ZN(
        DP_reg_pipe13_n123) );
  OAI21_X1 DP_reg_pipe13_U4 ( .B1(1'b1), .B2(DP_reg_pipe13_n99), .A(
        DP_reg_pipe13_n123), .ZN(DP_reg_pipe13_n75) );
  BUF_X1 DP_reg_pipe13_U3 ( .A(DP_n1), .Z(DP_reg_pipe13_n73) );
  BUF_X1 DP_reg_pipe13_U2 ( .A(DP_n1), .Z(DP_reg_pipe13_n74) );
  DFFR_X1 DP_reg_pipe13_Q_reg_0_ ( .D(DP_reg_pipe13_n98), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[0]), .QN(DP_reg_pipe13_n122) );
  DFFR_X1 DP_reg_pipe13_Q_reg_1_ ( .D(DP_reg_pipe13_n97), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[1]), .QN(DP_reg_pipe13_n121) );
  DFFR_X1 DP_reg_pipe13_Q_reg_2_ ( .D(DP_reg_pipe13_n96), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[2]), .QN(DP_reg_pipe13_n120) );
  DFFR_X1 DP_reg_pipe13_Q_reg_3_ ( .D(DP_reg_pipe13_n95), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[3]), .QN(DP_reg_pipe13_n119) );
  DFFR_X1 DP_reg_pipe13_Q_reg_4_ ( .D(DP_reg_pipe13_n94), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[4]), .QN(DP_reg_pipe13_n118) );
  DFFR_X1 DP_reg_pipe13_Q_reg_5_ ( .D(DP_reg_pipe13_n93), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[5]), .QN(DP_reg_pipe13_n117) );
  DFFR_X1 DP_reg_pipe13_Q_reg_6_ ( .D(DP_reg_pipe13_n92), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[6]), .QN(DP_reg_pipe13_n116) );
  DFFR_X1 DP_reg_pipe13_Q_reg_7_ ( .D(DP_reg_pipe13_n91), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[7]), .QN(DP_reg_pipe13_n115) );
  DFFR_X1 DP_reg_pipe13_Q_reg_8_ ( .D(DP_reg_pipe13_n90), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[8]), .QN(DP_reg_pipe13_n114) );
  DFFR_X1 DP_reg_pipe13_Q_reg_9_ ( .D(DP_reg_pipe13_n89), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[9]), .QN(DP_reg_pipe13_n113) );
  DFFR_X1 DP_reg_pipe13_Q_reg_10_ ( .D(DP_reg_pipe13_n88), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[10]), .QN(DP_reg_pipe13_n112) );
  DFFR_X1 DP_reg_pipe13_Q_reg_11_ ( .D(DP_reg_pipe13_n87), .CK(clk), .RN(
        DP_reg_pipe13_n74), .Q(DP_pipe13[11]), .QN(DP_reg_pipe13_n111) );
  DFFR_X1 DP_reg_pipe13_Q_reg_12_ ( .D(DP_reg_pipe13_n86), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[12]), .QN(DP_reg_pipe13_n110) );
  DFFR_X1 DP_reg_pipe13_Q_reg_13_ ( .D(DP_reg_pipe13_n85), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[13]), .QN(DP_reg_pipe13_n109) );
  DFFR_X1 DP_reg_pipe13_Q_reg_14_ ( .D(DP_reg_pipe13_n84), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[14]), .QN(DP_reg_pipe13_n108) );
  DFFR_X1 DP_reg_pipe13_Q_reg_15_ ( .D(DP_reg_pipe13_n83), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[15]), .QN(DP_reg_pipe13_n107) );
  DFFR_X1 DP_reg_pipe13_Q_reg_16_ ( .D(DP_reg_pipe13_n82), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[16]), .QN(DP_reg_pipe13_n106) );
  DFFR_X1 DP_reg_pipe13_Q_reg_17_ ( .D(DP_reg_pipe13_n81), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[17]), .QN(DP_reg_pipe13_n105) );
  DFFR_X1 DP_reg_pipe13_Q_reg_18_ ( .D(DP_reg_pipe13_n80), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[18]), .QN(DP_reg_pipe13_n104) );
  DFFR_X1 DP_reg_pipe13_Q_reg_19_ ( .D(DP_reg_pipe13_n79), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[19]), .QN(DP_reg_pipe13_n103) );
  DFFR_X1 DP_reg_pipe13_Q_reg_20_ ( .D(DP_reg_pipe13_n78), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[20]), .QN(DP_reg_pipe13_n102) );
  DFFR_X1 DP_reg_pipe13_Q_reg_21_ ( .D(DP_reg_pipe13_n77), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[21]), .QN(DP_reg_pipe13_n101) );
  DFFR_X1 DP_reg_pipe13_Q_reg_22_ ( .D(DP_reg_pipe13_n76), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[22]), .QN(DP_reg_pipe13_n100) );
  DFFR_X1 DP_reg_pipe13_Q_reg_23_ ( .D(DP_reg_pipe13_n75), .CK(clk), .RN(
        DP_reg_pipe13_n73), .Q(DP_pipe13[23]), .QN(DP_reg_pipe13_n99) );
  BUF_X1 DP_reg_out_U28 ( .A(delayed_controls_2__0_), .Z(DP_reg_out_n38) );
  BUF_X1 DP_reg_out_U27 ( .A(delayed_controls_2__0_), .Z(DP_reg_out_n37) );
  NAND2_X1 DP_reg_out_U26 ( .A1(DP_reg_out_n38), .A2(DP_y_out[0]), .ZN(
        DP_reg_out_n75) );
  OAI21_X1 DP_reg_out_U25 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n63), .A(
        DP_reg_out_n75), .ZN(DP_reg_out_n51) );
  NAND2_X1 DP_reg_out_U24 ( .A1(DP_y_out[10]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n65) );
  OAI21_X1 DP_reg_out_U23 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n53), .A(
        DP_reg_out_n65), .ZN(DP_reg_out_n41) );
  NAND2_X1 DP_reg_out_U22 ( .A1(DP_y_out[9]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n66) );
  OAI21_X1 DP_reg_out_U21 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n54), .A(
        DP_reg_out_n66), .ZN(DP_reg_out_n42) );
  NAND2_X1 DP_reg_out_U20 ( .A1(DP_y_out[8]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n67) );
  OAI21_X1 DP_reg_out_U19 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n55), .A(
        DP_reg_out_n67), .ZN(DP_reg_out_n43) );
  NAND2_X1 DP_reg_out_U18 ( .A1(DP_y_out[7]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n68) );
  OAI21_X1 DP_reg_out_U17 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n56), .A(
        DP_reg_out_n68), .ZN(DP_reg_out_n44) );
  NAND2_X1 DP_reg_out_U16 ( .A1(DP_y_out[6]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n69) );
  OAI21_X1 DP_reg_out_U15 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n57), .A(
        DP_reg_out_n69), .ZN(DP_reg_out_n45) );
  NAND2_X1 DP_reg_out_U14 ( .A1(DP_y_out[5]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n70) );
  OAI21_X1 DP_reg_out_U13 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n58), .A(
        DP_reg_out_n70), .ZN(DP_reg_out_n46) );
  NAND2_X1 DP_reg_out_U12 ( .A1(DP_y_out[4]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n71) );
  OAI21_X1 DP_reg_out_U11 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n59), .A(
        DP_reg_out_n71), .ZN(DP_reg_out_n47) );
  NAND2_X1 DP_reg_out_U10 ( .A1(DP_y_out[3]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n72) );
  OAI21_X1 DP_reg_out_U9 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n60), .A(
        DP_reg_out_n72), .ZN(DP_reg_out_n48) );
  NAND2_X1 DP_reg_out_U8 ( .A1(DP_y_out[2]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n73) );
  OAI21_X1 DP_reg_out_U7 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n61), .A(
        DP_reg_out_n73), .ZN(DP_reg_out_n49) );
  NAND2_X1 DP_reg_out_U6 ( .A1(DP_y_out[1]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n74) );
  OAI21_X1 DP_reg_out_U5 ( .B1(DP_reg_out_n38), .B2(DP_reg_out_n62), .A(
        DP_reg_out_n74), .ZN(DP_reg_out_n50) );
  NAND2_X1 DP_reg_out_U4 ( .A1(DP_y_out[11]), .A2(DP_reg_out_n37), .ZN(
        DP_reg_out_n64) );
  OAI21_X1 DP_reg_out_U3 ( .B1(DP_reg_out_n37), .B2(DP_reg_out_n52), .A(
        DP_reg_out_n64), .ZN(DP_reg_out_n40) );
  BUF_X1 DP_reg_out_U2 ( .A(DP_n6), .Z(DP_reg_out_n39) );
  DFFR_X1 DP_reg_out_Q_reg_0_ ( .D(DP_reg_out_n51), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[0]), .QN(DP_reg_out_n63) );
  DFFR_X1 DP_reg_out_Q_reg_1_ ( .D(DP_reg_out_n50), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[1]), .QN(DP_reg_out_n62) );
  DFFR_X1 DP_reg_out_Q_reg_2_ ( .D(DP_reg_out_n49), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[2]), .QN(DP_reg_out_n61) );
  DFFR_X1 DP_reg_out_Q_reg_3_ ( .D(DP_reg_out_n48), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[3]), .QN(DP_reg_out_n60) );
  DFFR_X1 DP_reg_out_Q_reg_4_ ( .D(DP_reg_out_n47), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[4]), .QN(DP_reg_out_n59) );
  DFFR_X1 DP_reg_out_Q_reg_5_ ( .D(DP_reg_out_n46), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[5]), .QN(DP_reg_out_n58) );
  DFFR_X1 DP_reg_out_Q_reg_6_ ( .D(DP_reg_out_n45), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[6]), .QN(DP_reg_out_n57) );
  DFFR_X1 DP_reg_out_Q_reg_7_ ( .D(DP_reg_out_n44), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[7]), .QN(DP_reg_out_n56) );
  DFFR_X1 DP_reg_out_Q_reg_8_ ( .D(DP_reg_out_n43), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[8]), .QN(DP_reg_out_n55) );
  DFFR_X1 DP_reg_out_Q_reg_9_ ( .D(DP_reg_out_n42), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[9]), .QN(DP_reg_out_n54) );
  DFFR_X1 DP_reg_out_Q_reg_10_ ( .D(DP_reg_out_n41), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[10]), .QN(DP_reg_out_n53) );
  DFFR_X1 DP_reg_out_Q_reg_11_ ( .D(DP_reg_out_n40), .CK(clk), .RN(
        DP_reg_out_n39), .Q(dOut[11]), .QN(DP_reg_out_n52) );
  XOR2_X1 DP_add_1_root_add_0_root_add_233_U2 ( .A(DP_pipe12[0]), .B(
        DP_pipe10[0]), .Z(DP_ff_part_0_) );
  AND2_X1 DP_add_1_root_add_0_root_add_233_U1 ( .A1(DP_pipe10[0]), .A2(
        DP_pipe12[0]), .ZN(DP_add_1_root_add_0_root_add_233_carry_1_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_1 ( .A(DP_pipe10[1]), .B(
        DP_pipe12[1]), .CI(DP_add_1_root_add_0_root_add_233_carry_1_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_2_), .S(DP_ff_part_1_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_2 ( .A(DP_pipe10[2]), .B(
        DP_pipe12[2]), .CI(DP_add_1_root_add_0_root_add_233_carry_2_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_3_), .S(DP_ff_part_2_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_3 ( .A(DP_pipe10[3]), .B(
        DP_pipe12[3]), .CI(DP_add_1_root_add_0_root_add_233_carry_3_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_4_), .S(DP_ff_part_3_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_4 ( .A(DP_pipe10[4]), .B(
        DP_pipe12[4]), .CI(DP_add_1_root_add_0_root_add_233_carry_4_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_5_), .S(DP_ff_part_4_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_5 ( .A(DP_pipe10[5]), .B(
        DP_pipe12[5]), .CI(DP_add_1_root_add_0_root_add_233_carry_5_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_6_), .S(DP_ff_part_5_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_6 ( .A(DP_pipe10[6]), .B(
        DP_pipe12[6]), .CI(DP_add_1_root_add_0_root_add_233_carry_6_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_7_), .S(DP_ff_part_6_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_7 ( .A(DP_pipe10[7]), .B(
        DP_pipe12[7]), .CI(DP_add_1_root_add_0_root_add_233_carry_7_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_8_), .S(DP_ff_part_7_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_8 ( .A(DP_pipe10[8]), .B(
        DP_pipe12[8]), .CI(DP_add_1_root_add_0_root_add_233_carry_8_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_9_), .S(DP_ff_part_8_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_9 ( .A(DP_pipe10[9]), .B(
        DP_pipe12[9]), .CI(DP_add_1_root_add_0_root_add_233_carry_9_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_10_), .S(DP_ff_part_9_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_10 ( .A(DP_pipe10[10]), .B(
        DP_pipe12[10]), .CI(DP_add_1_root_add_0_root_add_233_carry_10_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_11_), .S(DP_ff_part_10_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_11 ( .A(DP_pipe10[11]), .B(
        DP_pipe12[11]), .CI(DP_add_1_root_add_0_root_add_233_carry_11_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_12_), .S(DP_ff_part_11_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_12 ( .A(DP_pipe10[12]), .B(
        DP_pipe12[12]), .CI(DP_add_1_root_add_0_root_add_233_carry_12_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_13_), .S(DP_ff_part_12_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_13 ( .A(DP_pipe10[13]), .B(
        DP_pipe12[13]), .CI(DP_add_1_root_add_0_root_add_233_carry_13_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_14_), .S(DP_ff_part_13_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_14 ( .A(DP_pipe10[14]), .B(
        DP_pipe12[14]), .CI(DP_add_1_root_add_0_root_add_233_carry_14_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_15_), .S(DP_ff_part_14_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_15 ( .A(DP_pipe10[15]), .B(
        DP_pipe12[15]), .CI(DP_add_1_root_add_0_root_add_233_carry_15_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_16_), .S(DP_ff_part_15_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_16 ( .A(DP_pipe10[16]), .B(
        DP_pipe12[16]), .CI(DP_add_1_root_add_0_root_add_233_carry_16_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_17_), .S(DP_ff_part_16_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_17 ( .A(DP_pipe10[17]), .B(
        DP_pipe12[17]), .CI(DP_add_1_root_add_0_root_add_233_carry_17_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_18_), .S(DP_ff_part_17_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_18 ( .A(DP_pipe10[18]), .B(
        DP_pipe12[18]), .CI(DP_add_1_root_add_0_root_add_233_carry_18_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_19_), .S(DP_ff_part_18_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_19 ( .A(DP_pipe10[19]), .B(
        DP_pipe12[19]), .CI(DP_add_1_root_add_0_root_add_233_carry_19_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_20_), .S(DP_ff_part_19_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_20 ( .A(DP_pipe10[20]), .B(
        DP_pipe12[20]), .CI(DP_add_1_root_add_0_root_add_233_carry_20_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_21_), .S(DP_ff_part_20_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_21 ( .A(DP_pipe10[21]), .B(
        DP_pipe12[21]), .CI(DP_add_1_root_add_0_root_add_233_carry_21_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_22_), .S(DP_ff_part_21_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_22 ( .A(DP_pipe10[22]), .B(
        DP_pipe12[22]), .CI(DP_add_1_root_add_0_root_add_233_carry_22_), .CO(
        DP_add_1_root_add_0_root_add_233_carry_23_), .S(DP_ff_part_22_) );
  FA_X1 DP_add_1_root_add_0_root_add_233_U1_23 ( .A(DP_pipe10[23]), .B(
        DP_pipe12[23]), .CI(DP_add_1_root_add_0_root_add_233_carry_23_), .S(
        DP_ff_part_23_) );
  XOR2_X1 DP_add_2_root_add_0_root_add_233_U2 ( .A(DP_pipe13[0]), .B(
        DP_pipe11[0]), .Z(DP_ff_0_) );
  AND2_X1 DP_add_2_root_add_0_root_add_233_U1 ( .A1(DP_pipe11[0]), .A2(
        DP_pipe13[0]), .ZN(DP_add_2_root_add_0_root_add_233_carry_1_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_1 ( .A(DP_pipe11[1]), .B(
        DP_pipe13[1]), .CI(DP_add_2_root_add_0_root_add_233_carry_1_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_2_), .S(DP_ff_1_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_2 ( .A(DP_pipe11[2]), .B(
        DP_pipe13[2]), .CI(DP_add_2_root_add_0_root_add_233_carry_2_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_3_), .S(DP_ff_2_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_3 ( .A(DP_pipe11[3]), .B(
        DP_pipe13[3]), .CI(DP_add_2_root_add_0_root_add_233_carry_3_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_4_), .S(DP_ff_3_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_4 ( .A(DP_pipe11[4]), .B(
        DP_pipe13[4]), .CI(DP_add_2_root_add_0_root_add_233_carry_4_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_5_), .S(DP_ff_4_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_5 ( .A(DP_pipe11[5]), .B(
        DP_pipe13[5]), .CI(DP_add_2_root_add_0_root_add_233_carry_5_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_6_), .S(DP_ff_5_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_6 ( .A(DP_pipe11[6]), .B(
        DP_pipe13[6]), .CI(DP_add_2_root_add_0_root_add_233_carry_6_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_7_), .S(DP_ff_6_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_7 ( .A(DP_pipe11[7]), .B(
        DP_pipe13[7]), .CI(DP_add_2_root_add_0_root_add_233_carry_7_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_8_), .S(DP_ff_7_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_8 ( .A(DP_pipe11[8]), .B(
        DP_pipe13[8]), .CI(DP_add_2_root_add_0_root_add_233_carry_8_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_9_), .S(DP_ff_8_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_9 ( .A(DP_pipe11[9]), .B(
        DP_pipe13[9]), .CI(DP_add_2_root_add_0_root_add_233_carry_9_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_10_), .S(DP_ff_9_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_10 ( .A(DP_pipe11[10]), .B(
        DP_pipe13[10]), .CI(DP_add_2_root_add_0_root_add_233_carry_10_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_11_), .S(DP_ff_10_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_11 ( .A(DP_pipe11[11]), .B(
        DP_pipe13[11]), .CI(DP_add_2_root_add_0_root_add_233_carry_11_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_12_), .S(DP_ff_11_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_12 ( .A(DP_pipe11[12]), .B(
        DP_pipe13[12]), .CI(DP_add_2_root_add_0_root_add_233_carry_12_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_13_), .S(DP_ff_12_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_13 ( .A(DP_pipe11[13]), .B(
        DP_pipe13[13]), .CI(DP_add_2_root_add_0_root_add_233_carry_13_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_14_), .S(DP_ff_13_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_14 ( .A(DP_pipe11[14]), .B(
        DP_pipe13[14]), .CI(DP_add_2_root_add_0_root_add_233_carry_14_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_15_), .S(DP_ff_14_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_15 ( .A(DP_pipe11[15]), .B(
        DP_pipe13[15]), .CI(DP_add_2_root_add_0_root_add_233_carry_15_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_16_), .S(DP_ff_15_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_16 ( .A(DP_pipe11[16]), .B(
        DP_pipe13[16]), .CI(DP_add_2_root_add_0_root_add_233_carry_16_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_17_), .S(DP_ff_16_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_17 ( .A(DP_pipe11[17]), .B(
        DP_pipe13[17]), .CI(DP_add_2_root_add_0_root_add_233_carry_17_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_18_), .S(DP_ff_17_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_18 ( .A(DP_pipe11[18]), .B(
        DP_pipe13[18]), .CI(DP_add_2_root_add_0_root_add_233_carry_18_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_19_), .S(DP_ff_18_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_19 ( .A(DP_pipe11[19]), .B(
        DP_pipe13[19]), .CI(DP_add_2_root_add_0_root_add_233_carry_19_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_20_), .S(DP_ff_19_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_20 ( .A(DP_pipe11[20]), .B(
        DP_pipe13[20]), .CI(DP_add_2_root_add_0_root_add_233_carry_20_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_21_), .S(DP_ff_20_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_21 ( .A(DP_pipe11[21]), .B(
        DP_pipe13[21]), .CI(DP_add_2_root_add_0_root_add_233_carry_21_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_22_), .S(DP_ff_21_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_22 ( .A(DP_pipe11[22]), .B(
        DP_pipe13[22]), .CI(DP_add_2_root_add_0_root_add_233_carry_22_), .CO(
        DP_add_2_root_add_0_root_add_233_carry_23_), .S(DP_ff_22_) );
  FA_X1 DP_add_2_root_add_0_root_add_233_U1_23 ( .A(DP_pipe11[23]), .B(
        DP_pipe13[23]), .CI(DP_add_2_root_add_0_root_add_233_carry_23_), .S(
        DP_ff_23_) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U38 ( .A(DP_ff_1_), .ZN(
        DP_add_0_root_add_0_root_add_233_n35) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U37 ( .A(DP_ff_part_1_), .ZN(
        DP_add_0_root_add_0_root_add_233_n36) );
  OAI211_X1 DP_add_0_root_add_0_root_add_233_U36 ( .C1(DP_ff_1_), .C2(
        DP_ff_part_1_), .A(DP_ff_0_), .B(DP_ff_part_0_), .ZN(
        DP_add_0_root_add_0_root_add_233_n37) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U35 ( .B1(
        DP_add_0_root_add_0_root_add_233_n35), .B2(
        DP_add_0_root_add_0_root_add_233_n36), .A(
        DP_add_0_root_add_0_root_add_233_n37), .ZN(
        DP_add_0_root_add_0_root_add_233_n34) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U34 ( .A(
        DP_add_0_root_add_0_root_add_233_n34), .ZN(
        DP_add_0_root_add_0_root_add_233_n31) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U33 ( .A(DP_ff_2_), .ZN(
        DP_add_0_root_add_0_root_add_233_n32) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U32 ( .B1(DP_ff_2_), .B2(
        DP_add_0_root_add_0_root_add_233_n34), .A(DP_ff_part_2_), .ZN(
        DP_add_0_root_add_0_root_add_233_n33) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U31 ( .B1(
        DP_add_0_root_add_0_root_add_233_n31), .B2(
        DP_add_0_root_add_0_root_add_233_n32), .A(
        DP_add_0_root_add_0_root_add_233_n33), .ZN(
        DP_add_0_root_add_0_root_add_233_n30) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U30 ( .A(
        DP_add_0_root_add_0_root_add_233_n30), .ZN(
        DP_add_0_root_add_0_root_add_233_n27) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U29 ( .A(DP_ff_3_), .ZN(
        DP_add_0_root_add_0_root_add_233_n28) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U28 ( .B1(DP_ff_3_), .B2(
        DP_add_0_root_add_0_root_add_233_n30), .A(DP_ff_part_3_), .ZN(
        DP_add_0_root_add_0_root_add_233_n29) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U27 ( .B1(
        DP_add_0_root_add_0_root_add_233_n27), .B2(
        DP_add_0_root_add_0_root_add_233_n28), .A(
        DP_add_0_root_add_0_root_add_233_n29), .ZN(
        DP_add_0_root_add_0_root_add_233_n26) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U26 ( .A(
        DP_add_0_root_add_0_root_add_233_n26), .ZN(
        DP_add_0_root_add_0_root_add_233_n23) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U25 ( .A(DP_ff_4_), .ZN(
        DP_add_0_root_add_0_root_add_233_n24) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U24 ( .B1(DP_ff_4_), .B2(
        DP_add_0_root_add_0_root_add_233_n26), .A(DP_ff_part_4_), .ZN(
        DP_add_0_root_add_0_root_add_233_n25) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U23 ( .B1(
        DP_add_0_root_add_0_root_add_233_n23), .B2(
        DP_add_0_root_add_0_root_add_233_n24), .A(
        DP_add_0_root_add_0_root_add_233_n25), .ZN(
        DP_add_0_root_add_0_root_add_233_n22) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U22 ( .A(
        DP_add_0_root_add_0_root_add_233_n22), .ZN(
        DP_add_0_root_add_0_root_add_233_n19) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U21 ( .A(DP_ff_5_), .ZN(
        DP_add_0_root_add_0_root_add_233_n20) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U20 ( .B1(DP_ff_5_), .B2(
        DP_add_0_root_add_0_root_add_233_n22), .A(DP_ff_part_5_), .ZN(
        DP_add_0_root_add_0_root_add_233_n21) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U19 ( .B1(
        DP_add_0_root_add_0_root_add_233_n19), .B2(
        DP_add_0_root_add_0_root_add_233_n20), .A(
        DP_add_0_root_add_0_root_add_233_n21), .ZN(
        DP_add_0_root_add_0_root_add_233_n18) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U18 ( .A(
        DP_add_0_root_add_0_root_add_233_n18), .ZN(
        DP_add_0_root_add_0_root_add_233_n15) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U17 ( .A(DP_ff_6_), .ZN(
        DP_add_0_root_add_0_root_add_233_n16) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U16 ( .B1(DP_ff_6_), .B2(
        DP_add_0_root_add_0_root_add_233_n18), .A(DP_ff_part_6_), .ZN(
        DP_add_0_root_add_0_root_add_233_n17) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U15 ( .B1(
        DP_add_0_root_add_0_root_add_233_n15), .B2(
        DP_add_0_root_add_0_root_add_233_n16), .A(
        DP_add_0_root_add_0_root_add_233_n17), .ZN(
        DP_add_0_root_add_0_root_add_233_n12) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U14 ( .B1(DP_ff_7_), .B2(
        DP_add_0_root_add_0_root_add_233_n12), .A(DP_ff_part_7_), .ZN(
        DP_add_0_root_add_0_root_add_233_n14) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U13 ( .A(
        DP_add_0_root_add_0_root_add_233_n14), .ZN(
        DP_add_0_root_add_0_root_add_233_n13) );
  AOI21_X1 DP_add_0_root_add_0_root_add_233_U12 ( .B1(
        DP_add_0_root_add_0_root_add_233_n12), .B2(DP_ff_7_), .A(
        DP_add_0_root_add_0_root_add_233_n13), .ZN(
        DP_add_0_root_add_0_root_add_233_n8) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U11 ( .A(DP_ff_8_), .ZN(
        DP_add_0_root_add_0_root_add_233_n9) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U10 ( .A(
        DP_add_0_root_add_0_root_add_233_n8), .ZN(
        DP_add_0_root_add_0_root_add_233_n11) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U9 ( .B1(DP_ff_8_), .B2(
        DP_add_0_root_add_0_root_add_233_n11), .A(DP_ff_part_8_), .ZN(
        DP_add_0_root_add_0_root_add_233_n10) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U8 ( .B1(
        DP_add_0_root_add_0_root_add_233_n8), .B2(
        DP_add_0_root_add_0_root_add_233_n9), .A(
        DP_add_0_root_add_0_root_add_233_n10), .ZN(
        DP_add_0_root_add_0_root_add_233_n5) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U7 ( .B1(DP_ff_9_), .B2(
        DP_add_0_root_add_0_root_add_233_n5), .A(DP_ff_part_9_), .ZN(
        DP_add_0_root_add_0_root_add_233_n7) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U6 ( .A(
        DP_add_0_root_add_0_root_add_233_n7), .ZN(
        DP_add_0_root_add_0_root_add_233_n6) );
  AOI21_X1 DP_add_0_root_add_0_root_add_233_U5 ( .B1(
        DP_add_0_root_add_0_root_add_233_n5), .B2(DP_ff_9_), .A(
        DP_add_0_root_add_0_root_add_233_n6), .ZN(
        DP_add_0_root_add_0_root_add_233_n1) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U4 ( .A(DP_ff_10_), .ZN(
        DP_add_0_root_add_0_root_add_233_n2) );
  INV_X1 DP_add_0_root_add_0_root_add_233_U3 ( .A(
        DP_add_0_root_add_0_root_add_233_n1), .ZN(
        DP_add_0_root_add_0_root_add_233_n4) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U2 ( .B1(DP_ff_10_), .B2(
        DP_add_0_root_add_0_root_add_233_n4), .A(DP_ff_part_10_), .ZN(
        DP_add_0_root_add_0_root_add_233_n3) );
  OAI21_X1 DP_add_0_root_add_0_root_add_233_U1 ( .B1(
        DP_add_0_root_add_0_root_add_233_n1), .B2(
        DP_add_0_root_add_0_root_add_233_n2), .A(
        DP_add_0_root_add_0_root_add_233_n3), .ZN(
        DP_add_0_root_add_0_root_add_233_carry_11_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_11 ( .A(DP_ff_11_), .B(
        DP_ff_part_11_), .CI(DP_add_0_root_add_0_root_add_233_carry_11_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_12_), .S(DP_y_0_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_12 ( .A(DP_ff_12_), .B(
        DP_ff_part_12_), .CI(DP_add_0_root_add_0_root_add_233_carry_12_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_13_), .S(DP_y_1_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_13 ( .A(DP_ff_13_), .B(
        DP_ff_part_13_), .CI(DP_add_0_root_add_0_root_add_233_carry_13_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_14_), .S(DP_y_2_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_14 ( .A(DP_ff_14_), .B(
        DP_ff_part_14_), .CI(DP_add_0_root_add_0_root_add_233_carry_14_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_15_), .S(DP_y_3_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_15 ( .A(DP_ff_15_), .B(
        DP_ff_part_15_), .CI(DP_add_0_root_add_0_root_add_233_carry_15_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_16_), .S(DP_y_4_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_16 ( .A(DP_ff_16_), .B(
        DP_ff_part_16_), .CI(DP_add_0_root_add_0_root_add_233_carry_16_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_17_), .S(DP_y_5_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_17 ( .A(DP_ff_17_), .B(
        DP_ff_part_17_), .CI(DP_add_0_root_add_0_root_add_233_carry_17_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_18_), .S(DP_y_6_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_18 ( .A(DP_ff_18_), .B(
        DP_ff_part_18_), .CI(DP_add_0_root_add_0_root_add_233_carry_18_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_19_), .S(DP_y_7_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_19 ( .A(DP_ff_19_), .B(
        DP_ff_part_19_), .CI(DP_add_0_root_add_0_root_add_233_carry_19_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_20_), .S(DP_y_8_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_20 ( .A(DP_ff_20_), .B(
        DP_ff_part_20_), .CI(DP_add_0_root_add_0_root_add_233_carry_20_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_21_), .S(DP_y_9_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_21 ( .A(DP_ff_21_), .B(
        DP_ff_part_21_), .CI(DP_add_0_root_add_0_root_add_233_carry_21_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_22_), .S(DP_y_10_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_22 ( .A(DP_ff_22_), .B(
        DP_ff_part_22_), .CI(DP_add_0_root_add_0_root_add_233_carry_22_), .CO(
        DP_add_0_root_add_0_root_add_233_carry_23_), .S(DP_y_11_) );
  FA_X1 DP_add_0_root_add_0_root_add_233_U1_23 ( .A(DP_ff_23_), .B(
        DP_ff_part_23_), .CI(DP_add_0_root_add_0_root_add_233_carry_23_), .S(
        DP_y_23) );
  INV_X1 DP_mult_219_U1959 ( .A(DP_coeff_pipe03[1]), .ZN(DP_mult_219_n2159) );
  NOR2_X1 DP_mult_219_U1958 ( .A1(DP_mult_219_n2159), .A2(DP_coeff_pipe03[0]), 
        .ZN(DP_mult_219_n1636) );
  INV_X1 DP_mult_219_U1957 ( .A(DP_coeff_pipe03[2]), .ZN(DP_mult_219_n1742) );
  XNOR2_X1 DP_mult_219_U1956 ( .A(DP_coeff_pipe03[1]), .B(DP_mult_219_n1742), 
        .ZN(DP_mult_219_n2157) );
  AOI221_X1 DP_mult_219_U1955 ( .B1(DP_pipe03[1]), .B2(DP_mult_219_n1563), 
        .C1(DP_mult_219_n1396), .C2(DP_mult_219_n1555), .A(DP_mult_219_n1742), 
        .ZN(DP_mult_219_n2160) );
  INV_X1 DP_mult_219_U1954 ( .A(DP_coeff_pipe03[0]), .ZN(DP_mult_219_n2158) );
  INV_X1 DP_mult_219_U1953 ( .A(DP_pipe03[2]), .ZN(DP_mult_219_n1661) );
  INV_X1 DP_mult_219_U1952 ( .A(DP_mult_219_n1397), .ZN(DP_mult_219_n1650) );
  OAI22_X1 DP_mult_219_U1951 ( .A1(DP_mult_219_n1554), .A2(DP_mult_219_n1661), 
        .B1(DP_mult_219_n1564), .B2(DP_mult_219_n1650), .ZN(DP_mult_219_n2162)
         );
  AOI211_X1 DP_mult_219_U1950 ( .C1(DP_pipe03[1]), .C2(DP_mult_219_n1561), .A(
        DP_mult_219_n2162), .B(DP_pipe03[0]), .ZN(DP_mult_219_n2161) );
  AND2_X1 DP_mult_219_U1949 ( .A1(DP_mult_219_n2160), .A2(DP_mult_219_n2161), 
        .ZN(DP_mult_219_n2153) );
  INV_X1 DP_mult_219_U1948 ( .A(DP_mult_219_n1395), .ZN(DP_mult_219_n1657) );
  INV_X1 DP_mult_219_U1947 ( .A(DP_pipe03[1]), .ZN(DP_mult_219_n1649) );
  OAI22_X1 DP_mult_219_U1946 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1657), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1649), .ZN(DP_mult_219_n2156)
         );
  AOI221_X1 DP_mult_219_U1945 ( .B1(DP_pipe03[3]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[2]), .C2(DP_mult_219_n1563), .A(DP_mult_219_n2156), .ZN(
        DP_mult_219_n2155) );
  XNOR2_X1 DP_mult_219_U1944 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2155), 
        .ZN(DP_mult_219_n2154) );
  AOI222_X1 DP_mult_219_U1943 ( .A1(DP_mult_219_n2153), .A2(DP_mult_219_n2154), 
        .B1(DP_mult_219_n2153), .B2(DP_mult_219_n688), .C1(DP_mult_219_n688), 
        .C2(DP_mult_219_n2154), .ZN(DP_mult_219_n2148) );
  INV_X1 DP_mult_219_U1942 ( .A(DP_mult_219_n1394), .ZN(DP_mult_219_n1660) );
  OAI22_X1 DP_mult_219_U1941 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1660), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1661), .ZN(DP_mult_219_n2152)
         );
  AOI221_X1 DP_mult_219_U1940 ( .B1(DP_pipe03[4]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[3]), .C2(DP_mult_219_n1563), .A(DP_mult_219_n2152), .ZN(
        DP_mult_219_n2151) );
  XNOR2_X1 DP_mult_219_U1939 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2151), 
        .ZN(DP_mult_219_n2149) );
  INV_X1 DP_mult_219_U1938 ( .A(DP_mult_219_n686), .ZN(DP_mult_219_n2150) );
  OAI222_X1 DP_mult_219_U1937 ( .A1(DP_mult_219_n2148), .A2(DP_mult_219_n2149), 
        .B1(DP_mult_219_n2148), .B2(DP_mult_219_n2150), .C1(DP_mult_219_n2150), 
        .C2(DP_mult_219_n2149), .ZN(DP_mult_219_n2144) );
  INV_X1 DP_mult_219_U1936 ( .A(DP_mult_219_n1393), .ZN(DP_mult_219_n1664) );
  INV_X1 DP_mult_219_U1935 ( .A(DP_pipe03[3]), .ZN(DP_mult_219_n1665) );
  OAI22_X1 DP_mult_219_U1934 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1664), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1665), .ZN(DP_mult_219_n2147)
         );
  AOI221_X1 DP_mult_219_U1933 ( .B1(DP_pipe03[5]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[4]), .C2(DP_mult_219_n1563), .A(DP_mult_219_n2147), .ZN(
        DP_mult_219_n2146) );
  XNOR2_X1 DP_mult_219_U1932 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2146), 
        .ZN(DP_mult_219_n2145) );
  AOI222_X1 DP_mult_219_U1931 ( .A1(DP_mult_219_n2144), .A2(DP_mult_219_n2145), 
        .B1(DP_mult_219_n2144), .B2(DP_mult_219_n684), .C1(DP_mult_219_n684), 
        .C2(DP_mult_219_n2145), .ZN(DP_mult_219_n2139) );
  INV_X1 DP_mult_219_U1930 ( .A(DP_mult_219_n1392), .ZN(DP_mult_219_n1668) );
  INV_X1 DP_mult_219_U1929 ( .A(DP_pipe03[4]), .ZN(DP_mult_219_n1669) );
  OAI22_X1 DP_mult_219_U1928 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1668), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1669), .ZN(DP_mult_219_n2143)
         );
  AOI221_X1 DP_mult_219_U1927 ( .B1(DP_pipe03[6]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[5]), .C2(DP_mult_219_n1563), .A(DP_mult_219_n2143), .ZN(
        DP_mult_219_n2142) );
  XNOR2_X1 DP_mult_219_U1926 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2142), 
        .ZN(DP_mult_219_n2140) );
  INV_X1 DP_mult_219_U1925 ( .A(DP_mult_219_n680), .ZN(DP_mult_219_n2141) );
  OAI222_X1 DP_mult_219_U1924 ( .A1(DP_mult_219_n2139), .A2(DP_mult_219_n2140), 
        .B1(DP_mult_219_n2139), .B2(DP_mult_219_n2141), .C1(DP_mult_219_n2141), 
        .C2(DP_mult_219_n2140), .ZN(DP_mult_219_n2135) );
  INV_X1 DP_mult_219_U1923 ( .A(DP_mult_219_n1391), .ZN(DP_mult_219_n1672) );
  INV_X1 DP_mult_219_U1922 ( .A(DP_pipe03[5]), .ZN(DP_mult_219_n1673) );
  OAI22_X1 DP_mult_219_U1921 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1672), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1673), .ZN(DP_mult_219_n2138)
         );
  AOI221_X1 DP_mult_219_U1920 ( .B1(DP_pipe03[7]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[6]), .C2(DP_mult_219_n1563), .A(DP_mult_219_n2138), .ZN(
        DP_mult_219_n2137) );
  XNOR2_X1 DP_mult_219_U1919 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2137), 
        .ZN(DP_mult_219_n2136) );
  AOI222_X1 DP_mult_219_U1918 ( .A1(DP_mult_219_n2135), .A2(DP_mult_219_n2136), 
        .B1(DP_mult_219_n2135), .B2(DP_mult_219_n676), .C1(DP_mult_219_n676), 
        .C2(DP_mult_219_n2136), .ZN(DP_mult_219_n2130) );
  INV_X1 DP_mult_219_U1917 ( .A(DP_mult_219_n1390), .ZN(DP_mult_219_n1676) );
  INV_X1 DP_mult_219_U1916 ( .A(DP_pipe03[6]), .ZN(DP_mult_219_n1677) );
  OAI22_X1 DP_mult_219_U1915 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1676), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1677), .ZN(DP_mult_219_n2134)
         );
  AOI221_X1 DP_mult_219_U1914 ( .B1(DP_pipe03[8]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[7]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2134), .ZN(
        DP_mult_219_n2133) );
  XNOR2_X1 DP_mult_219_U1913 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2133), 
        .ZN(DP_mult_219_n2131) );
  INV_X1 DP_mult_219_U1912 ( .A(DP_mult_219_n672), .ZN(DP_mult_219_n2132) );
  OAI222_X1 DP_mult_219_U1911 ( .A1(DP_mult_219_n2130), .A2(DP_mult_219_n2131), 
        .B1(DP_mult_219_n2130), .B2(DP_mult_219_n2132), .C1(DP_mult_219_n2132), 
        .C2(DP_mult_219_n2131), .ZN(DP_mult_219_n2126) );
  INV_X1 DP_mult_219_U1910 ( .A(DP_mult_219_n1389), .ZN(DP_mult_219_n1680) );
  INV_X1 DP_mult_219_U1909 ( .A(DP_pipe03[7]), .ZN(DP_mult_219_n1681) );
  OAI22_X1 DP_mult_219_U1908 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1680), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1681), .ZN(DP_mult_219_n2129)
         );
  AOI221_X1 DP_mult_219_U1907 ( .B1(DP_pipe03[9]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[8]), .C2(DP_mult_219_n1563), .A(DP_mult_219_n2129), .ZN(
        DP_mult_219_n2128) );
  XNOR2_X1 DP_mult_219_U1906 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2128), 
        .ZN(DP_mult_219_n2127) );
  AOI222_X1 DP_mult_219_U1905 ( .A1(DP_mult_219_n2126), .A2(DP_mult_219_n2127), 
        .B1(DP_mult_219_n2126), .B2(DP_mult_219_n666), .C1(DP_mult_219_n666), 
        .C2(DP_mult_219_n2127), .ZN(DP_mult_219_n2121) );
  INV_X1 DP_mult_219_U1904 ( .A(DP_mult_219_n1388), .ZN(DP_mult_219_n1684) );
  INV_X1 DP_mult_219_U1903 ( .A(DP_pipe03[8]), .ZN(DP_mult_219_n1685) );
  OAI22_X1 DP_mult_219_U1902 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1684), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1685), .ZN(DP_mult_219_n2125)
         );
  AOI221_X1 DP_mult_219_U1901 ( .B1(DP_pipe03[10]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[9]), .C2(DP_mult_219_n1563), .A(DP_mult_219_n2125), .ZN(
        DP_mult_219_n2124) );
  XNOR2_X1 DP_mult_219_U1900 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2124), 
        .ZN(DP_mult_219_n2122) );
  INV_X1 DP_mult_219_U1899 ( .A(DP_mult_219_n660), .ZN(DP_mult_219_n2123) );
  OAI222_X1 DP_mult_219_U1898 ( .A1(DP_mult_219_n2121), .A2(DP_mult_219_n2122), 
        .B1(DP_mult_219_n2121), .B2(DP_mult_219_n2123), .C1(DP_mult_219_n2123), 
        .C2(DP_mult_219_n2122), .ZN(DP_mult_219_n2117) );
  INV_X1 DP_mult_219_U1897 ( .A(DP_mult_219_n1387), .ZN(DP_mult_219_n1688) );
  INV_X1 DP_mult_219_U1896 ( .A(DP_pipe03[9]), .ZN(DP_mult_219_n1689) );
  OAI22_X1 DP_mult_219_U1895 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1688), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1689), .ZN(DP_mult_219_n2120)
         );
  AOI221_X1 DP_mult_219_U1894 ( .B1(DP_pipe03[11]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[10]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2120), 
        .ZN(DP_mult_219_n2119) );
  XNOR2_X1 DP_mult_219_U1893 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2119), 
        .ZN(DP_mult_219_n2118) );
  AOI222_X1 DP_mult_219_U1892 ( .A1(DP_mult_219_n2117), .A2(DP_mult_219_n2118), 
        .B1(DP_mult_219_n2117), .B2(DP_mult_219_n654), .C1(DP_mult_219_n654), 
        .C2(DP_mult_219_n2118), .ZN(DP_mult_219_n2112) );
  INV_X1 DP_mult_219_U1891 ( .A(DP_mult_219_n1386), .ZN(DP_mult_219_n1692) );
  INV_X1 DP_mult_219_U1890 ( .A(DP_pipe03[10]), .ZN(DP_mult_219_n1693) );
  OAI22_X1 DP_mult_219_U1889 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1692), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1693), .ZN(DP_mult_219_n2116)
         );
  AOI221_X1 DP_mult_219_U1888 ( .B1(DP_pipe03[12]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[11]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2116), 
        .ZN(DP_mult_219_n2115) );
  XNOR2_X1 DP_mult_219_U1887 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2115), 
        .ZN(DP_mult_219_n2113) );
  INV_X1 DP_mult_219_U1886 ( .A(DP_mult_219_n646), .ZN(DP_mult_219_n2114) );
  OAI222_X1 DP_mult_219_U1885 ( .A1(DP_mult_219_n2112), .A2(DP_mult_219_n2113), 
        .B1(DP_mult_219_n2112), .B2(DP_mult_219_n2114), .C1(DP_mult_219_n2114), 
        .C2(DP_mult_219_n2113), .ZN(DP_mult_219_n2108) );
  INV_X1 DP_mult_219_U1884 ( .A(DP_mult_219_n1385), .ZN(DP_mult_219_n1696) );
  INV_X1 DP_mult_219_U1883 ( .A(DP_pipe03[11]), .ZN(DP_mult_219_n1697) );
  OAI22_X1 DP_mult_219_U1882 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1696), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1697), .ZN(DP_mult_219_n2111)
         );
  AOI221_X1 DP_mult_219_U1881 ( .B1(DP_pipe03[13]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[12]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2111), 
        .ZN(DP_mult_219_n2110) );
  XNOR2_X1 DP_mult_219_U1880 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2110), 
        .ZN(DP_mult_219_n2109) );
  AOI222_X1 DP_mult_219_U1879 ( .A1(DP_mult_219_n2108), .A2(DP_mult_219_n2109), 
        .B1(DP_mult_219_n2108), .B2(DP_mult_219_n638), .C1(DP_mult_219_n638), 
        .C2(DP_mult_219_n2109), .ZN(DP_mult_219_n2103) );
  INV_X1 DP_mult_219_U1878 ( .A(DP_mult_219_n1384), .ZN(DP_mult_219_n1700) );
  INV_X1 DP_mult_219_U1877 ( .A(DP_pipe03[12]), .ZN(DP_mult_219_n1701) );
  OAI22_X1 DP_mult_219_U1876 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1700), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1701), .ZN(DP_mult_219_n2107)
         );
  AOI221_X1 DP_mult_219_U1875 ( .B1(DP_pipe03[14]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[13]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2107), 
        .ZN(DP_mult_219_n2106) );
  XNOR2_X1 DP_mult_219_U1874 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2106), 
        .ZN(DP_mult_219_n2104) );
  INV_X1 DP_mult_219_U1873 ( .A(DP_mult_219_n630), .ZN(DP_mult_219_n2105) );
  OAI222_X1 DP_mult_219_U1872 ( .A1(DP_mult_219_n2103), .A2(DP_mult_219_n2104), 
        .B1(DP_mult_219_n2103), .B2(DP_mult_219_n2105), .C1(DP_mult_219_n2105), 
        .C2(DP_mult_219_n2104), .ZN(DP_mult_219_n2099) );
  INV_X1 DP_mult_219_U1871 ( .A(DP_mult_219_n1383), .ZN(DP_mult_219_n1704) );
  INV_X1 DP_mult_219_U1870 ( .A(DP_pipe03[13]), .ZN(DP_mult_219_n1705) );
  OAI22_X1 DP_mult_219_U1869 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1704), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1705), .ZN(DP_mult_219_n2102)
         );
  AOI221_X1 DP_mult_219_U1868 ( .B1(DP_pipe03[15]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[14]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2102), 
        .ZN(DP_mult_219_n2101) );
  XNOR2_X1 DP_mult_219_U1867 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2101), 
        .ZN(DP_mult_219_n2100) );
  AOI222_X1 DP_mult_219_U1866 ( .A1(DP_mult_219_n2099), .A2(DP_mult_219_n2100), 
        .B1(DP_mult_219_n2099), .B2(DP_mult_219_n620), .C1(DP_mult_219_n620), 
        .C2(DP_mult_219_n2100), .ZN(DP_mult_219_n2094) );
  INV_X1 DP_mult_219_U1865 ( .A(DP_mult_219_n1382), .ZN(DP_mult_219_n1708) );
  INV_X1 DP_mult_219_U1864 ( .A(DP_pipe03[14]), .ZN(DP_mult_219_n1709) );
  OAI22_X1 DP_mult_219_U1863 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1708), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1709), .ZN(DP_mult_219_n2098)
         );
  AOI221_X1 DP_mult_219_U1862 ( .B1(DP_pipe03[16]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[15]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2098), 
        .ZN(DP_mult_219_n2097) );
  XNOR2_X1 DP_mult_219_U1861 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2097), 
        .ZN(DP_mult_219_n2095) );
  INV_X1 DP_mult_219_U1860 ( .A(DP_mult_219_n610), .ZN(DP_mult_219_n2096) );
  OAI222_X1 DP_mult_219_U1859 ( .A1(DP_mult_219_n2094), .A2(DP_mult_219_n2095), 
        .B1(DP_mult_219_n2094), .B2(DP_mult_219_n2096), .C1(DP_mult_219_n2096), 
        .C2(DP_mult_219_n2095), .ZN(DP_mult_219_n2090) );
  INV_X1 DP_mult_219_U1858 ( .A(DP_mult_219_n1381), .ZN(DP_mult_219_n1712) );
  INV_X1 DP_mult_219_U1857 ( .A(DP_pipe03[15]), .ZN(DP_mult_219_n1713) );
  OAI22_X1 DP_mult_219_U1856 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1712), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1713), .ZN(DP_mult_219_n2093)
         );
  AOI221_X1 DP_mult_219_U1855 ( .B1(DP_pipe03[17]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[16]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2093), 
        .ZN(DP_mult_219_n2092) );
  XNOR2_X1 DP_mult_219_U1854 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2092), 
        .ZN(DP_mult_219_n2091) );
  AOI222_X1 DP_mult_219_U1853 ( .A1(DP_mult_219_n2090), .A2(DP_mult_219_n2091), 
        .B1(DP_mult_219_n2090), .B2(DP_mult_219_n600), .C1(DP_mult_219_n600), 
        .C2(DP_mult_219_n2091), .ZN(DP_mult_219_n2085) );
  INV_X1 DP_mult_219_U1852 ( .A(DP_mult_219_n1380), .ZN(DP_mult_219_n1716) );
  INV_X1 DP_mult_219_U1851 ( .A(DP_pipe03[16]), .ZN(DP_mult_219_n1717) );
  OAI22_X1 DP_mult_219_U1850 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1716), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1717), .ZN(DP_mult_219_n2089)
         );
  AOI221_X1 DP_mult_219_U1849 ( .B1(DP_pipe03[18]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[17]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2089), 
        .ZN(DP_mult_219_n2088) );
  XNOR2_X1 DP_mult_219_U1848 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2088), 
        .ZN(DP_mult_219_n2086) );
  INV_X1 DP_mult_219_U1847 ( .A(DP_mult_219_n588), .ZN(DP_mult_219_n2087) );
  OAI222_X1 DP_mult_219_U1846 ( .A1(DP_mult_219_n2085), .A2(DP_mult_219_n2086), 
        .B1(DP_mult_219_n2085), .B2(DP_mult_219_n2087), .C1(DP_mult_219_n2087), 
        .C2(DP_mult_219_n2086), .ZN(DP_mult_219_n2081) );
  INV_X1 DP_mult_219_U1845 ( .A(DP_mult_219_n1379), .ZN(DP_mult_219_n1720) );
  INV_X1 DP_mult_219_U1844 ( .A(DP_pipe03[17]), .ZN(DP_mult_219_n1721) );
  OAI22_X1 DP_mult_219_U1843 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1720), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1721), .ZN(DP_mult_219_n2084)
         );
  AOI221_X1 DP_mult_219_U1842 ( .B1(DP_pipe03[19]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[18]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2084), 
        .ZN(DP_mult_219_n2083) );
  XNOR2_X1 DP_mult_219_U1841 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2083), 
        .ZN(DP_mult_219_n2082) );
  AOI222_X1 DP_mult_219_U1840 ( .A1(DP_mult_219_n2081), .A2(DP_mult_219_n2082), 
        .B1(DP_mult_219_n2081), .B2(DP_mult_219_n576), .C1(DP_mult_219_n576), 
        .C2(DP_mult_219_n2082), .ZN(DP_mult_219_n2080) );
  INV_X1 DP_mult_219_U1839 ( .A(DP_mult_219_n2080), .ZN(DP_mult_219_n2076) );
  INV_X1 DP_mult_219_U1838 ( .A(DP_mult_219_n1378), .ZN(DP_mult_219_n1724) );
  INV_X1 DP_mult_219_U1837 ( .A(DP_pipe03[18]), .ZN(DP_mult_219_n1725) );
  OAI22_X1 DP_mult_219_U1836 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1724), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1725), .ZN(DP_mult_219_n2079)
         );
  AOI221_X1 DP_mult_219_U1835 ( .B1(DP_pipe03[20]), .B2(DP_mult_219_n1561), 
        .C1(DP_pipe03[19]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2079), 
        .ZN(DP_mult_219_n2078) );
  XNOR2_X1 DP_mult_219_U1834 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n2078), 
        .ZN(DP_mult_219_n2077) );
  AOI222_X1 DP_mult_219_U1833 ( .A1(DP_mult_219_n2076), .A2(DP_mult_219_n2077), 
        .B1(DP_mult_219_n2076), .B2(DP_mult_219_n564), .C1(DP_mult_219_n564), 
        .C2(DP_mult_219_n2077), .ZN(DP_mult_219_n2071) );
  INV_X1 DP_mult_219_U1832 ( .A(DP_mult_219_n1377), .ZN(DP_mult_219_n1728) );
  INV_X1 DP_mult_219_U1831 ( .A(DP_pipe03[19]), .ZN(DP_mult_219_n1729) );
  OAI22_X1 DP_mult_219_U1830 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1728), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1729), .ZN(DP_mult_219_n2075)
         );
  AOI221_X1 DP_mult_219_U1829 ( .B1(DP_mult_219_n1561), .B2(DP_pipe03[21]), 
        .C1(DP_pipe03[20]), .C2(DP_mult_219_n1562), .A(DP_mult_219_n2075), 
        .ZN(DP_mult_219_n2074) );
  XNOR2_X1 DP_mult_219_U1828 ( .A(DP_mult_219_n1742), .B(DP_mult_219_n2074), 
        .ZN(DP_mult_219_n2072) );
  INV_X1 DP_mult_219_U1827 ( .A(DP_mult_219_n550), .ZN(DP_mult_219_n2073) );
  OAI222_X1 DP_mult_219_U1826 ( .A1(DP_mult_219_n2071), .A2(DP_mult_219_n2072), 
        .B1(DP_mult_219_n2071), .B2(DP_mult_219_n2073), .C1(DP_mult_219_n2073), 
        .C2(DP_mult_219_n2072), .ZN(DP_mult_219_n326) );
  XNOR2_X1 DP_mult_219_U1825 ( .A(DP_coeff_pipe03[21]), .B(DP_mult_219_n1608), 
        .ZN(DP_mult_219_n2067) );
  INV_X1 DP_mult_219_U1824 ( .A(DP_mult_219_n2067), .ZN(DP_mult_219_n2070) );
  XNOR2_X1 DP_mult_219_U1823 ( .A(DP_coeff_pipe03[21]), .B(DP_coeff_pipe03[22]), .ZN(DP_mult_219_n2069) );
  XNOR2_X1 DP_mult_219_U1822 ( .A(DP_coeff_pipe03[22]), .B(DP_mult_219_n1611), 
        .ZN(DP_mult_219_n2068) );
  NAND3_X1 DP_mult_219_U1821 ( .A1(DP_mult_219_n2067), .A2(DP_mult_219_n2068), 
        .A3(DP_mult_219_n2069), .ZN(DP_mult_219_n1629) );
  INV_X1 DP_mult_219_U1820 ( .A(DP_pipe03[21]), .ZN(DP_mult_219_n1643) );
  OAI22_X1 DP_mult_219_U1819 ( .A1(DP_mult_219_n1548), .A2(DP_mult_219_n1619), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1643), .ZN(DP_mult_219_n2066)
         );
  AOI221_X1 DP_mult_219_U1818 ( .B1(DP_pipe03[22]), .B2(DP_mult_219_n1560), 
        .C1(DP_mult_219_n1375), .C2(DP_mult_219_n1549), .A(DP_mult_219_n2066), 
        .ZN(DP_mult_219_n2065) );
  XOR2_X1 DP_mult_219_U1817 ( .A(DP_mult_219_n1611), .B(DP_mult_219_n2065), 
        .Z(DP_mult_219_n1627) );
  INV_X1 DP_mult_219_U1816 ( .A(DP_mult_219_n1627), .ZN(DP_mult_219_n351) );
  INV_X1 DP_mult_219_U1815 ( .A(DP_mult_219_n356), .ZN(DP_mult_219_n360) );
  OAI22_X1 DP_mult_219_U1814 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1712), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1713), .ZN(DP_mult_219_n2064)
         );
  AOI221_X1 DP_mult_219_U1813 ( .B1(DP_pipe03[17]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[16]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2064), 
        .ZN(DP_mult_219_n2063) );
  XOR2_X1 DP_mult_219_U1812 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2063), 
        .Z(DP_mult_219_n374) );
  INV_X1 DP_mult_219_U1811 ( .A(DP_mult_219_n374), .ZN(DP_mult_219_n368) );
  INV_X1 DP_mult_219_U1810 ( .A(DP_mult_219_n387), .ZN(DP_mult_219_n395) );
  OAI22_X1 DP_mult_219_U1809 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1688), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1689), .ZN(DP_mult_219_n2062)
         );
  AOI221_X1 DP_mult_219_U1808 ( .B1(DP_pipe03[11]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[10]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2062), 
        .ZN(DP_mult_219_n2061) );
  XOR2_X1 DP_mult_219_U1807 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2061), 
        .Z(DP_mult_219_n421) );
  INV_X1 DP_mult_219_U1806 ( .A(DP_mult_219_n421), .ZN(DP_mult_219_n411) );
  OAI22_X1 DP_mult_219_U1805 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1676), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1677), .ZN(DP_mult_219_n2060)
         );
  AOI221_X1 DP_mult_219_U1804 ( .B1(DP_pipe03[8]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[7]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2060), .ZN(
        DP_mult_219_n2059) );
  XOR2_X1 DP_mult_219_U1803 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2059), 
        .Z(DP_mult_219_n454) );
  INV_X1 DP_mult_219_U1802 ( .A(DP_mult_219_n454), .ZN(DP_mult_219_n442) );
  OAI21_X1 DP_mult_219_U1801 ( .B1(DP_mult_219_n1561), .B2(DP_mult_219_n1563), 
        .A(DP_mult_219_n1615), .ZN(DP_mult_219_n2058) );
  OAI221_X1 DP_mult_219_U1800 ( .B1(DP_mult_219_n1619), .B2(DP_mult_219_n1639), 
        .C1(DP_mult_219_n1620), .C2(DP_mult_219_n1564), .A(DP_mult_219_n2058), 
        .ZN(DP_mult_219_n2057) );
  XOR2_X1 DP_mult_219_U1799 ( .A(DP_mult_219_n2057), .B(DP_mult_219_n1742), 
        .Z(DP_mult_219_n2056) );
  NOR2_X1 DP_mult_219_U1798 ( .A1(DP_mult_219_n2056), .A2(DP_mult_219_n519), 
        .ZN(DP_mult_219_n493) );
  INV_X1 DP_mult_219_U1797 ( .A(DP_mult_219_n493), .ZN(DP_mult_219_n479) );
  XNOR2_X1 DP_mult_219_U1796 ( .A(DP_mult_219_n519), .B(DP_mult_219_n2056), 
        .ZN(DP_mult_219_n506) );
  INV_X1 DP_mult_219_U1795 ( .A(DP_pipe03[20]), .ZN(DP_mult_219_n1640) );
  OAI22_X1 DP_mult_219_U1794 ( .A1(DP_mult_219_n1556), .A2(DP_mult_219_n1640), 
        .B1(DP_mult_219_n1550), .B2(DP_mult_219_n1643), .ZN(DP_mult_219_n2055)
         );
  AOI221_X1 DP_mult_219_U1793 ( .B1(DP_pipe03[22]), .B2(DP_mult_219_n1559), 
        .C1(DP_mult_219_n1376), .C2(DP_mult_219_n1549), .A(DP_mult_219_n2055), 
        .ZN(DP_mult_219_n2054) );
  XNOR2_X1 DP_mult_219_U1792 ( .A(DP_coeff_pipe03[23]), .B(DP_mult_219_n2054), 
        .ZN(DP_mult_219_n729) );
  OAI22_X1 DP_mult_219_U1791 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1728), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1729), .ZN(DP_mult_219_n2053)
         );
  AOI221_X1 DP_mult_219_U1790 ( .B1(DP_pipe03[21]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[20]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2053), 
        .ZN(DP_mult_219_n2052) );
  XNOR2_X1 DP_mult_219_U1789 ( .A(DP_coeff_pipe03[23]), .B(DP_mult_219_n2052), 
        .ZN(DP_mult_219_n730) );
  OAI22_X1 DP_mult_219_U1788 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1724), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1725), .ZN(DP_mult_219_n2051)
         );
  AOI221_X1 DP_mult_219_U1787 ( .B1(DP_pipe03[20]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[19]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2051), 
        .ZN(DP_mult_219_n2050) );
  XNOR2_X1 DP_mult_219_U1786 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2050), 
        .ZN(DP_mult_219_n731) );
  OAI22_X1 DP_mult_219_U1785 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1720), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1721), .ZN(DP_mult_219_n2049)
         );
  AOI221_X1 DP_mult_219_U1784 ( .B1(DP_pipe03[19]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[18]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2049), 
        .ZN(DP_mult_219_n2048) );
  XNOR2_X1 DP_mult_219_U1783 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2048), 
        .ZN(DP_mult_219_n732) );
  OAI22_X1 DP_mult_219_U1782 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1716), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1717), .ZN(DP_mult_219_n2047)
         );
  AOI221_X1 DP_mult_219_U1781 ( .B1(DP_pipe03[18]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[17]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2047), 
        .ZN(DP_mult_219_n2046) );
  XNOR2_X1 DP_mult_219_U1780 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2046), 
        .ZN(DP_mult_219_n733) );
  OAI22_X1 DP_mult_219_U1779 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1708), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1709), .ZN(DP_mult_219_n2045)
         );
  AOI221_X1 DP_mult_219_U1778 ( .B1(DP_pipe03[16]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[15]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2045), 
        .ZN(DP_mult_219_n2044) );
  XNOR2_X1 DP_mult_219_U1777 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2044), 
        .ZN(DP_mult_219_n734) );
  OAI22_X1 DP_mult_219_U1776 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1704), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1705), .ZN(DP_mult_219_n2043)
         );
  AOI221_X1 DP_mult_219_U1775 ( .B1(DP_pipe03[15]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[14]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2043), 
        .ZN(DP_mult_219_n2042) );
  XNOR2_X1 DP_mult_219_U1774 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2042), 
        .ZN(DP_mult_219_n735) );
  OAI22_X1 DP_mult_219_U1773 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1700), 
        .B1(DP_mult_219_n1556), .B2(DP_mult_219_n1701), .ZN(DP_mult_219_n2041)
         );
  AOI221_X1 DP_mult_219_U1772 ( .B1(DP_pipe03[14]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[13]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2041), 
        .ZN(DP_mult_219_n2040) );
  XNOR2_X1 DP_mult_219_U1771 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2040), 
        .ZN(DP_mult_219_n736) );
  OAI22_X1 DP_mult_219_U1770 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1696), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1697), .ZN(DP_mult_219_n2039)
         );
  AOI221_X1 DP_mult_219_U1769 ( .B1(DP_pipe03[13]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[12]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2039), 
        .ZN(DP_mult_219_n2038) );
  XNOR2_X1 DP_mult_219_U1768 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2038), 
        .ZN(DP_mult_219_n737) );
  OAI22_X1 DP_mult_219_U1767 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1692), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1693), .ZN(DP_mult_219_n2037)
         );
  AOI221_X1 DP_mult_219_U1766 ( .B1(DP_pipe03[12]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[11]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2037), 
        .ZN(DP_mult_219_n2036) );
  XNOR2_X1 DP_mult_219_U1765 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2036), 
        .ZN(DP_mult_219_n738) );
  OAI22_X1 DP_mult_219_U1764 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1684), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1685), .ZN(DP_mult_219_n2035)
         );
  AOI221_X1 DP_mult_219_U1763 ( .B1(DP_pipe03[10]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[9]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2035), .ZN(
        DP_mult_219_n2034) );
  XNOR2_X1 DP_mult_219_U1762 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2034), 
        .ZN(DP_mult_219_n739) );
  OAI22_X1 DP_mult_219_U1761 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1680), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1681), .ZN(DP_mult_219_n2033)
         );
  AOI221_X1 DP_mult_219_U1760 ( .B1(DP_pipe03[9]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[8]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2033), .ZN(
        DP_mult_219_n2032) );
  XNOR2_X1 DP_mult_219_U1759 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2032), 
        .ZN(DP_mult_219_n740) );
  OAI22_X1 DP_mult_219_U1758 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1672), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1673), .ZN(DP_mult_219_n2031)
         );
  AOI221_X1 DP_mult_219_U1757 ( .B1(DP_pipe03[7]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[6]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2031), .ZN(
        DP_mult_219_n2030) );
  XNOR2_X1 DP_mult_219_U1756 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2030), 
        .ZN(DP_mult_219_n741) );
  OAI22_X1 DP_mult_219_U1755 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1668), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1669), .ZN(DP_mult_219_n2029)
         );
  AOI221_X1 DP_mult_219_U1754 ( .B1(DP_pipe03[6]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[5]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2029), .ZN(
        DP_mult_219_n2028) );
  XNOR2_X1 DP_mult_219_U1753 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2028), 
        .ZN(DP_mult_219_n742) );
  OAI22_X1 DP_mult_219_U1752 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1664), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1665), .ZN(DP_mult_219_n2027)
         );
  AOI221_X1 DP_mult_219_U1751 ( .B1(DP_pipe03[5]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[4]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2027), .ZN(
        DP_mult_219_n2026) );
  XNOR2_X1 DP_mult_219_U1750 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2026), 
        .ZN(DP_mult_219_n743) );
  OAI22_X1 DP_mult_219_U1749 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1660), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1661), .ZN(DP_mult_219_n2025)
         );
  AOI221_X1 DP_mult_219_U1748 ( .B1(DP_pipe03[4]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[3]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2025), .ZN(
        DP_mult_219_n2024) );
  XNOR2_X1 DP_mult_219_U1747 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2024), 
        .ZN(DP_mult_219_n744) );
  OAI22_X1 DP_mult_219_U1746 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1657), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1649), .ZN(DP_mult_219_n2023)
         );
  AOI221_X1 DP_mult_219_U1745 ( .B1(DP_pipe03[3]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[2]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2023), .ZN(
        DP_mult_219_n2022) );
  XNOR2_X1 DP_mult_219_U1744 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2022), 
        .ZN(DP_mult_219_n745) );
  INV_X1 DP_mult_219_U1743 ( .A(DP_mult_219_n1396), .ZN(DP_mult_219_n1653) );
  INV_X1 DP_mult_219_U1742 ( .A(DP_pipe03[0]), .ZN(DP_mult_219_n1647) );
  OAI22_X1 DP_mult_219_U1741 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1653), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1567), .ZN(DP_mult_219_n2021)
         );
  AOI221_X1 DP_mult_219_U1740 ( .B1(DP_pipe03[2]), .B2(DP_mult_219_n1559), 
        .C1(DP_pipe03[1]), .C2(DP_mult_219_n1560), .A(DP_mult_219_n2021), .ZN(
        DP_mult_219_n2020) );
  XNOR2_X1 DP_mult_219_U1739 ( .A(DP_mult_219_n1610), .B(DP_mult_219_n2020), 
        .ZN(DP_mult_219_n746) );
  OAI222_X1 DP_mult_219_U1738 ( .A1(DP_mult_219_n1548), .A2(DP_mult_219_n1649), 
        .B1(DP_mult_219_n1550), .B2(DP_mult_219_n1566), .C1(DP_mult_219_n1558), 
        .C2(DP_mult_219_n1650), .ZN(DP_mult_219_n2019) );
  XNOR2_X1 DP_mult_219_U1737 ( .A(DP_mult_219_n2019), .B(DP_mult_219_n1611), 
        .ZN(DP_mult_219_n747) );
  OAI22_X1 DP_mult_219_U1736 ( .A1(DP_mult_219_n1548), .A2(DP_mult_219_n1567), 
        .B1(DP_mult_219_n1558), .B2(DP_mult_219_n1567), .ZN(DP_mult_219_n2018)
         );
  XNOR2_X1 DP_mult_219_U1735 ( .A(DP_mult_219_n2018), .B(DP_mult_219_n1611), 
        .ZN(DP_mult_219_n748) );
  XOR2_X1 DP_mult_219_U1734 ( .A(DP_coeff_pipe03[18]), .B(DP_mult_219_n1607), 
        .Z(DP_mult_219_n2017) );
  XOR2_X1 DP_mult_219_U1733 ( .A(DP_coeff_pipe03[19]), .B(DP_mult_219_n1608), 
        .Z(DP_mult_219_n2016) );
  XNOR2_X1 DP_mult_219_U1732 ( .A(DP_coeff_pipe03[18]), .B(DP_coeff_pipe03[19]), .ZN(DP_mult_219_n2015) );
  NAND3_X1 DP_mult_219_U1731 ( .A1(DP_mult_219_n2017), .A2(DP_mult_219_n2016), 
        .A3(DP_mult_219_n2015), .ZN(DP_mult_219_n1967) );
  INV_X1 DP_mult_219_U1730 ( .A(DP_mult_219_n2017), .ZN(DP_mult_219_n2014) );
  OAI21_X1 DP_mult_219_U1729 ( .B1(DP_mult_219_n1594), .B2(DP_mult_219_n1595), 
        .A(DP_mult_219_n1615), .ZN(DP_mult_219_n2013) );
  OAI221_X1 DP_mult_219_U1728 ( .B1(DP_mult_219_n1617), .B2(DP_mult_219_n1597), 
        .C1(DP_mult_219_n1620), .C2(DP_mult_219_n1593), .A(DP_mult_219_n2013), 
        .ZN(DP_mult_219_n2012) );
  XNOR2_X1 DP_mult_219_U1727 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n2012), 
        .ZN(DP_mult_219_n749) );
  INV_X1 DP_mult_219_U1726 ( .A(DP_mult_219_n1374), .ZN(DP_mult_219_n1633) );
  INV_X1 DP_mult_219_U1725 ( .A(DP_pipe03[22]), .ZN(DP_mult_219_n1634) );
  OAI22_X1 DP_mult_219_U1724 ( .A1(DP_mult_219_n1633), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1634), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n2011)
         );
  AOI221_X1 DP_mult_219_U1723 ( .B1(DP_mult_219_n1594), .B2(DP_mult_219_n1614), 
        .C1(DP_mult_219_n1595), .C2(DP_mult_219_n1615), .A(DP_mult_219_n2011), 
        .ZN(DP_mult_219_n2010) );
  XNOR2_X1 DP_mult_219_U1722 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n2010), 
        .ZN(DP_mult_219_n750) );
  OAI22_X1 DP_mult_219_U1721 ( .A1(DP_mult_219_n1617), .A2(DP_mult_219_n1541), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n2009)
         );
  AOI221_X1 DP_mult_219_U1720 ( .B1(DP_mult_219_n1595), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1542), .C2(DP_mult_219_n1375), .A(DP_mult_219_n2009), 
        .ZN(DP_mult_219_n2008) );
  XNOR2_X1 DP_mult_219_U1719 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n2008), 
        .ZN(DP_mult_219_n751) );
  OAI22_X1 DP_mult_219_U1718 ( .A1(DP_mult_219_n1640), .A2(DP_mult_219_n1597), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1543), .ZN(DP_mult_219_n2007)
         );
  AOI221_X1 DP_mult_219_U1717 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1542), .C2(DP_mult_219_n1376), .A(DP_mult_219_n2007), 
        .ZN(DP_mult_219_n2006) );
  XNOR2_X1 DP_mult_219_U1716 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n2006), 
        .ZN(DP_mult_219_n752) );
  OAI22_X1 DP_mult_219_U1715 ( .A1(DP_mult_219_n1728), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1729), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n2005)
         );
  AOI221_X1 DP_mult_219_U1714 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[21]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[20]), .A(DP_mult_219_n2005), 
        .ZN(DP_mult_219_n2004) );
  XNOR2_X1 DP_mult_219_U1713 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n2004), 
        .ZN(DP_mult_219_n753) );
  OAI22_X1 DP_mult_219_U1712 ( .A1(DP_mult_219_n1724), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1725), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n2003)
         );
  AOI221_X1 DP_mult_219_U1711 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[20]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[19]), .A(DP_mult_219_n2003), 
        .ZN(DP_mult_219_n2002) );
  XNOR2_X1 DP_mult_219_U1710 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n2002), 
        .ZN(DP_mult_219_n754) );
  OAI22_X1 DP_mult_219_U1709 ( .A1(DP_mult_219_n1720), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1721), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n2001)
         );
  AOI221_X1 DP_mult_219_U1708 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[19]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[18]), .A(DP_mult_219_n2001), 
        .ZN(DP_mult_219_n2000) );
  XNOR2_X1 DP_mult_219_U1707 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n2000), 
        .ZN(DP_mult_219_n755) );
  OAI22_X1 DP_mult_219_U1706 ( .A1(DP_mult_219_n1716), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1717), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n1999)
         );
  AOI221_X1 DP_mult_219_U1705 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[18]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[17]), .A(DP_mult_219_n1999), 
        .ZN(DP_mult_219_n1998) );
  XNOR2_X1 DP_mult_219_U1704 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n1998), 
        .ZN(DP_mult_219_n756) );
  OAI22_X1 DP_mult_219_U1703 ( .A1(DP_mult_219_n1712), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1713), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n1997)
         );
  AOI221_X1 DP_mult_219_U1702 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[17]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[16]), .A(DP_mult_219_n1997), 
        .ZN(DP_mult_219_n1996) );
  XNOR2_X1 DP_mult_219_U1701 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n1996), 
        .ZN(DP_mult_219_n757) );
  OAI22_X1 DP_mult_219_U1700 ( .A1(DP_mult_219_n1708), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1709), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n1995)
         );
  AOI221_X1 DP_mult_219_U1699 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[16]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[15]), .A(DP_mult_219_n1995), 
        .ZN(DP_mult_219_n1994) );
  XNOR2_X1 DP_mult_219_U1698 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n1994), 
        .ZN(DP_mult_219_n758) );
  OAI22_X1 DP_mult_219_U1697 ( .A1(DP_mult_219_n1704), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1705), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n1993)
         );
  AOI221_X1 DP_mult_219_U1696 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[15]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[14]), .A(DP_mult_219_n1993), 
        .ZN(DP_mult_219_n1992) );
  XNOR2_X1 DP_mult_219_U1695 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n1992), 
        .ZN(DP_mult_219_n759) );
  OAI22_X1 DP_mult_219_U1694 ( .A1(DP_mult_219_n1700), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1701), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n1991)
         );
  AOI221_X1 DP_mult_219_U1693 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[14]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[13]), .A(DP_mult_219_n1991), 
        .ZN(DP_mult_219_n1990) );
  XNOR2_X1 DP_mult_219_U1692 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n1990), 
        .ZN(DP_mult_219_n760) );
  OAI22_X1 DP_mult_219_U1691 ( .A1(DP_mult_219_n1696), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1697), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n1989)
         );
  AOI221_X1 DP_mult_219_U1690 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[13]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[12]), .A(DP_mult_219_n1989), 
        .ZN(DP_mult_219_n1988) );
  XNOR2_X1 DP_mult_219_U1689 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n1988), 
        .ZN(DP_mult_219_n761) );
  OAI22_X1 DP_mult_219_U1688 ( .A1(DP_mult_219_n1692), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1693), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1987)
         );
  AOI221_X1 DP_mult_219_U1687 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[12]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[11]), .A(DP_mult_219_n1987), 
        .ZN(DP_mult_219_n1986) );
  XNOR2_X1 DP_mult_219_U1686 ( .A(DP_mult_219_n1609), .B(DP_mult_219_n1986), 
        .ZN(DP_mult_219_n762) );
  OAI22_X1 DP_mult_219_U1685 ( .A1(DP_mult_219_n1688), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1689), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1985)
         );
  AOI221_X1 DP_mult_219_U1684 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[11]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[10]), .A(DP_mult_219_n1985), 
        .ZN(DP_mult_219_n1984) );
  XNOR2_X1 DP_mult_219_U1683 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1984), 
        .ZN(DP_mult_219_n763) );
  OAI22_X1 DP_mult_219_U1682 ( .A1(DP_mult_219_n1684), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1685), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1983)
         );
  AOI221_X1 DP_mult_219_U1681 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[10]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[9]), .A(DP_mult_219_n1983), .ZN(
        DP_mult_219_n1982) );
  XNOR2_X1 DP_mult_219_U1680 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1982), 
        .ZN(DP_mult_219_n764) );
  OAI22_X1 DP_mult_219_U1679 ( .A1(DP_mult_219_n1680), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1681), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1981)
         );
  AOI221_X1 DP_mult_219_U1678 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[9]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[8]), .A(DP_mult_219_n1981), .ZN(
        DP_mult_219_n1980) );
  XNOR2_X1 DP_mult_219_U1677 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1980), 
        .ZN(DP_mult_219_n765) );
  OAI22_X1 DP_mult_219_U1676 ( .A1(DP_mult_219_n1676), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1677), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1979)
         );
  AOI221_X1 DP_mult_219_U1675 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[8]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[7]), .A(DP_mult_219_n1979), .ZN(
        DP_mult_219_n1978) );
  XNOR2_X1 DP_mult_219_U1674 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1978), 
        .ZN(DP_mult_219_n766) );
  OAI22_X1 DP_mult_219_U1673 ( .A1(DP_mult_219_n1672), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1673), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1977)
         );
  AOI221_X1 DP_mult_219_U1672 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[7]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[6]), .A(DP_mult_219_n1977), .ZN(
        DP_mult_219_n1976) );
  XNOR2_X1 DP_mult_219_U1671 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1976), 
        .ZN(DP_mult_219_n767) );
  OAI22_X1 DP_mult_219_U1670 ( .A1(DP_mult_219_n1668), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1669), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1975)
         );
  AOI221_X1 DP_mult_219_U1669 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[6]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[5]), .A(DP_mult_219_n1975), .ZN(
        DP_mult_219_n1974) );
  XNOR2_X1 DP_mult_219_U1668 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1974), 
        .ZN(DP_mult_219_n768) );
  OAI22_X1 DP_mult_219_U1667 ( .A1(DP_mult_219_n1664), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1665), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1973)
         );
  AOI221_X1 DP_mult_219_U1666 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[5]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[4]), .A(DP_mult_219_n1973), .ZN(
        DP_mult_219_n1972) );
  XNOR2_X1 DP_mult_219_U1665 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1972), 
        .ZN(DP_mult_219_n769) );
  OAI22_X1 DP_mult_219_U1664 ( .A1(DP_mult_219_n1660), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1661), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1971)
         );
  AOI221_X1 DP_mult_219_U1663 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[4]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[3]), .A(DP_mult_219_n1971), .ZN(
        DP_mult_219_n1970) );
  XNOR2_X1 DP_mult_219_U1662 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1970), 
        .ZN(DP_mult_219_n770) );
  OAI22_X1 DP_mult_219_U1661 ( .A1(DP_mult_219_n1657), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1649), .B2(DP_mult_219_n1597), .ZN(DP_mult_219_n1969)
         );
  AOI221_X1 DP_mult_219_U1660 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[3]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[2]), .A(DP_mult_219_n1969), .ZN(
        DP_mult_219_n1968) );
  XNOR2_X1 DP_mult_219_U1659 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1968), 
        .ZN(DP_mult_219_n771) );
  OAI22_X1 DP_mult_219_U1658 ( .A1(DP_mult_219_n1653), .A2(DP_mult_219_n1593), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1596), .ZN(DP_mult_219_n1966)
         );
  AOI221_X1 DP_mult_219_U1657 ( .B1(DP_mult_219_n1594), .B2(DP_pipe03[2]), 
        .C1(DP_mult_219_n1595), .C2(DP_pipe03[1]), .A(DP_mult_219_n1966), .ZN(
        DP_mult_219_n1965) );
  XNOR2_X1 DP_mult_219_U1656 ( .A(DP_mult_219_n1608), .B(DP_mult_219_n1965), 
        .ZN(DP_mult_219_n772) );
  OAI222_X1 DP_mult_219_U1655 ( .A1(DP_mult_219_n1649), .A2(DP_mult_219_n1541), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1543), .C1(DP_mult_219_n1650), 
        .C2(DP_mult_219_n1593), .ZN(DP_mult_219_n1964) );
  XOR2_X1 DP_mult_219_U1654 ( .A(DP_mult_219_n1964), .B(DP_mult_219_n1608), 
        .Z(DP_mult_219_n773) );
  OAI22_X1 DP_mult_219_U1653 ( .A1(DP_mult_219_n1565), .A2(DP_mult_219_n1541), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1593), .ZN(DP_mult_219_n1963)
         );
  XOR2_X1 DP_mult_219_U1652 ( .A(DP_mult_219_n1963), .B(DP_mult_219_n1608), 
        .Z(DP_mult_219_n774) );
  XOR2_X1 DP_mult_219_U1651 ( .A(DP_coeff_pipe03[15]), .B(DP_mult_219_n1605), 
        .Z(DP_mult_219_n1962) );
  XNOR2_X1 DP_mult_219_U1650 ( .A(DP_coeff_pipe03[16]), .B(DP_mult_219_n1607), 
        .ZN(DP_mult_219_n1961) );
  XNOR2_X1 DP_mult_219_U1649 ( .A(DP_coeff_pipe03[15]), .B(DP_coeff_pipe03[16]), .ZN(DP_mult_219_n1960) );
  NAND3_X1 DP_mult_219_U1648 ( .A1(DP_mult_219_n1962), .A2(DP_mult_219_n1961), 
        .A3(DP_mult_219_n1960), .ZN(DP_mult_219_n1912) );
  INV_X1 DP_mult_219_U1647 ( .A(DP_mult_219_n1962), .ZN(DP_mult_219_n1959) );
  OAI21_X1 DP_mult_219_U1646 ( .B1(DP_mult_219_n1589), .B2(DP_mult_219_n1590), 
        .A(DP_mult_219_n1615), .ZN(DP_mult_219_n1958) );
  OAI221_X1 DP_mult_219_U1645 ( .B1(DP_mult_219_n1619), .B2(DP_mult_219_n1592), 
        .C1(DP_mult_219_n1617), .C2(DP_mult_219_n1588), .A(DP_mult_219_n1958), 
        .ZN(DP_mult_219_n1957) );
  XNOR2_X1 DP_mult_219_U1644 ( .A(DP_coeff_pipe03[17]), .B(DP_mult_219_n1957), 
        .ZN(DP_mult_219_n775) );
  OAI22_X1 DP_mult_219_U1643 ( .A1(DP_mult_219_n1633), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1634), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1956)
         );
  AOI221_X1 DP_mult_219_U1642 ( .B1(DP_mult_219_n1589), .B2(DP_mult_219_n1614), 
        .C1(DP_mult_219_n1590), .C2(DP_mult_219_n1615), .A(DP_mult_219_n1956), 
        .ZN(DP_mult_219_n1955) );
  XNOR2_X1 DP_mult_219_U1641 ( .A(DP_coeff_pipe03[17]), .B(DP_mult_219_n1955), 
        .ZN(DP_mult_219_n776) );
  OAI22_X1 DP_mult_219_U1640 ( .A1(DP_mult_219_n1617), .A2(DP_mult_219_n1534), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1954)
         );
  AOI221_X1 DP_mult_219_U1639 ( .B1(DP_mult_219_n1590), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1537), .C2(DP_mult_219_n1375), .A(DP_mult_219_n1954), 
        .ZN(DP_mult_219_n1953) );
  XNOR2_X1 DP_mult_219_U1638 ( .A(DP_coeff_pipe03[17]), .B(DP_mult_219_n1953), 
        .ZN(DP_mult_219_n777) );
  OAI22_X1 DP_mult_219_U1637 ( .A1(DP_mult_219_n1640), .A2(DP_mult_219_n1592), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1540), .ZN(DP_mult_219_n1952)
         );
  AOI221_X1 DP_mult_219_U1636 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1537), .C2(DP_mult_219_n1376), .A(DP_mult_219_n1952), 
        .ZN(DP_mult_219_n1951) );
  XNOR2_X1 DP_mult_219_U1635 ( .A(DP_coeff_pipe03[17]), .B(DP_mult_219_n1951), 
        .ZN(DP_mult_219_n778) );
  OAI22_X1 DP_mult_219_U1634 ( .A1(DP_mult_219_n1728), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1729), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1950)
         );
  AOI221_X1 DP_mult_219_U1633 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[21]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[20]), .A(DP_mult_219_n1950), 
        .ZN(DP_mult_219_n1949) );
  XNOR2_X1 DP_mult_219_U1632 ( .A(DP_coeff_pipe03[17]), .B(DP_mult_219_n1949), 
        .ZN(DP_mult_219_n779) );
  OAI22_X1 DP_mult_219_U1631 ( .A1(DP_mult_219_n1724), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1725), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1948)
         );
  AOI221_X1 DP_mult_219_U1630 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[20]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[19]), .A(DP_mult_219_n1948), 
        .ZN(DP_mult_219_n1947) );
  XNOR2_X1 DP_mult_219_U1629 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1947), 
        .ZN(DP_mult_219_n780) );
  OAI22_X1 DP_mult_219_U1628 ( .A1(DP_mult_219_n1720), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1721), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1946)
         );
  AOI221_X1 DP_mult_219_U1627 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[19]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[18]), .A(DP_mult_219_n1946), 
        .ZN(DP_mult_219_n1945) );
  XNOR2_X1 DP_mult_219_U1626 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1945), 
        .ZN(DP_mult_219_n781) );
  OAI22_X1 DP_mult_219_U1625 ( .A1(DP_mult_219_n1716), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1717), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1944)
         );
  AOI221_X1 DP_mult_219_U1624 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[18]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[17]), .A(DP_mult_219_n1944), 
        .ZN(DP_mult_219_n1943) );
  XNOR2_X1 DP_mult_219_U1623 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1943), 
        .ZN(DP_mult_219_n782) );
  OAI22_X1 DP_mult_219_U1622 ( .A1(DP_mult_219_n1712), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1713), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1942)
         );
  AOI221_X1 DP_mult_219_U1621 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[17]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[16]), .A(DP_mult_219_n1942), 
        .ZN(DP_mult_219_n1941) );
  XNOR2_X1 DP_mult_219_U1620 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1941), 
        .ZN(DP_mult_219_n783) );
  OAI22_X1 DP_mult_219_U1619 ( .A1(DP_mult_219_n1708), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1709), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1940)
         );
  AOI221_X1 DP_mult_219_U1618 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[16]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[15]), .A(DP_mult_219_n1940), 
        .ZN(DP_mult_219_n1939) );
  XNOR2_X1 DP_mult_219_U1617 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1939), 
        .ZN(DP_mult_219_n784) );
  OAI22_X1 DP_mult_219_U1616 ( .A1(DP_mult_219_n1704), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1705), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1938)
         );
  AOI221_X1 DP_mult_219_U1615 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[15]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[14]), .A(DP_mult_219_n1938), 
        .ZN(DP_mult_219_n1937) );
  XNOR2_X1 DP_mult_219_U1614 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1937), 
        .ZN(DP_mult_219_n785) );
  OAI22_X1 DP_mult_219_U1613 ( .A1(DP_mult_219_n1700), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1701), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1936)
         );
  AOI221_X1 DP_mult_219_U1612 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[14]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[13]), .A(DP_mult_219_n1936), 
        .ZN(DP_mult_219_n1935) );
  XNOR2_X1 DP_mult_219_U1611 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1935), 
        .ZN(DP_mult_219_n786) );
  OAI22_X1 DP_mult_219_U1610 ( .A1(DP_mult_219_n1696), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1697), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1934)
         );
  AOI221_X1 DP_mult_219_U1609 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[13]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[12]), .A(DP_mult_219_n1934), 
        .ZN(DP_mult_219_n1933) );
  XNOR2_X1 DP_mult_219_U1608 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1933), 
        .ZN(DP_mult_219_n787) );
  OAI22_X1 DP_mult_219_U1607 ( .A1(DP_mult_219_n1692), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1693), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1932)
         );
  AOI221_X1 DP_mult_219_U1606 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[12]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[11]), .A(DP_mult_219_n1932), 
        .ZN(DP_mult_219_n1931) );
  XNOR2_X1 DP_mult_219_U1605 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1931), 
        .ZN(DP_mult_219_n788) );
  OAI22_X1 DP_mult_219_U1604 ( .A1(DP_mult_219_n1688), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1689), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1930)
         );
  AOI221_X1 DP_mult_219_U1603 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[11]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[10]), .A(DP_mult_219_n1930), 
        .ZN(DP_mult_219_n1929) );
  XNOR2_X1 DP_mult_219_U1602 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1929), 
        .ZN(DP_mult_219_n789) );
  OAI22_X1 DP_mult_219_U1601 ( .A1(DP_mult_219_n1684), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1685), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1928)
         );
  AOI221_X1 DP_mult_219_U1600 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[10]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[9]), .A(DP_mult_219_n1928), .ZN(
        DP_mult_219_n1927) );
  XNOR2_X1 DP_mult_219_U1599 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1927), 
        .ZN(DP_mult_219_n790) );
  OAI22_X1 DP_mult_219_U1598 ( .A1(DP_mult_219_n1680), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1681), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1926)
         );
  AOI221_X1 DP_mult_219_U1597 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[9]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[8]), .A(DP_mult_219_n1926), .ZN(
        DP_mult_219_n1925) );
  XNOR2_X1 DP_mult_219_U1596 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1925), 
        .ZN(DP_mult_219_n791) );
  OAI22_X1 DP_mult_219_U1595 ( .A1(DP_mult_219_n1676), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1677), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1924)
         );
  AOI221_X1 DP_mult_219_U1594 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[8]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[7]), .A(DP_mult_219_n1924), .ZN(
        DP_mult_219_n1923) );
  XNOR2_X1 DP_mult_219_U1593 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1923), 
        .ZN(DP_mult_219_n792) );
  OAI22_X1 DP_mult_219_U1592 ( .A1(DP_mult_219_n1672), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1673), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1922)
         );
  AOI221_X1 DP_mult_219_U1591 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[7]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[6]), .A(DP_mult_219_n1922), .ZN(
        DP_mult_219_n1921) );
  XNOR2_X1 DP_mult_219_U1590 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1921), 
        .ZN(DP_mult_219_n793) );
  OAI22_X1 DP_mult_219_U1589 ( .A1(DP_mult_219_n1668), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1669), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1920)
         );
  AOI221_X1 DP_mult_219_U1588 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[6]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[5]), .A(DP_mult_219_n1920), .ZN(
        DP_mult_219_n1919) );
  XNOR2_X1 DP_mult_219_U1587 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1919), 
        .ZN(DP_mult_219_n794) );
  OAI22_X1 DP_mult_219_U1586 ( .A1(DP_mult_219_n1664), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1665), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1918)
         );
  AOI221_X1 DP_mult_219_U1585 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[5]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[4]), .A(DP_mult_219_n1918), .ZN(
        DP_mult_219_n1917) );
  XNOR2_X1 DP_mult_219_U1584 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1917), 
        .ZN(DP_mult_219_n795) );
  OAI22_X1 DP_mult_219_U1583 ( .A1(DP_mult_219_n1660), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1661), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1916)
         );
  AOI221_X1 DP_mult_219_U1582 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[4]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[3]), .A(DP_mult_219_n1916), .ZN(
        DP_mult_219_n1915) );
  XNOR2_X1 DP_mult_219_U1581 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1915), 
        .ZN(DP_mult_219_n796) );
  OAI22_X1 DP_mult_219_U1580 ( .A1(DP_mult_219_n1657), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1649), .B2(DP_mult_219_n1592), .ZN(DP_mult_219_n1914)
         );
  AOI221_X1 DP_mult_219_U1579 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[3]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[2]), .A(DP_mult_219_n1914), .ZN(
        DP_mult_219_n1913) );
  XNOR2_X1 DP_mult_219_U1578 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1913), 
        .ZN(DP_mult_219_n797) );
  OAI22_X1 DP_mult_219_U1577 ( .A1(DP_mult_219_n1653), .A2(DP_mult_219_n1588), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1591), .ZN(DP_mult_219_n1911)
         );
  AOI221_X1 DP_mult_219_U1576 ( .B1(DP_mult_219_n1589), .B2(DP_pipe03[2]), 
        .C1(DP_mult_219_n1590), .C2(DP_pipe03[1]), .A(DP_mult_219_n1911), .ZN(
        DP_mult_219_n1910) );
  XNOR2_X1 DP_mult_219_U1575 ( .A(DP_mult_219_n1606), .B(DP_mult_219_n1910), 
        .ZN(DP_mult_219_n798) );
  OAI222_X1 DP_mult_219_U1574 ( .A1(DP_mult_219_n1649), .A2(DP_mult_219_n1534), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1540), .C1(DP_mult_219_n1650), 
        .C2(DP_mult_219_n1588), .ZN(DP_mult_219_n1909) );
  XNOR2_X1 DP_mult_219_U1573 ( .A(DP_mult_219_n1909), .B(DP_mult_219_n1607), 
        .ZN(DP_mult_219_n799) );
  OAI22_X1 DP_mult_219_U1572 ( .A1(DP_mult_219_n1565), .A2(DP_mult_219_n1534), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1588), .ZN(DP_mult_219_n1908)
         );
  XNOR2_X1 DP_mult_219_U1571 ( .A(DP_mult_219_n1908), .B(DP_mult_219_n1607), 
        .ZN(DP_mult_219_n800) );
  XOR2_X1 DP_mult_219_U1570 ( .A(DP_coeff_pipe03[12]), .B(DP_mult_219_n1603), 
        .Z(DP_mult_219_n1907) );
  XNOR2_X1 DP_mult_219_U1569 ( .A(DP_coeff_pipe03[13]), .B(DP_mult_219_n1605), 
        .ZN(DP_mult_219_n1906) );
  XNOR2_X1 DP_mult_219_U1568 ( .A(DP_coeff_pipe03[12]), .B(DP_coeff_pipe03[13]), .ZN(DP_mult_219_n1905) );
  NAND3_X1 DP_mult_219_U1567 ( .A1(DP_mult_219_n1907), .A2(DP_mult_219_n1906), 
        .A3(DP_mult_219_n1905), .ZN(DP_mult_219_n1857) );
  INV_X1 DP_mult_219_U1566 ( .A(DP_mult_219_n1907), .ZN(DP_mult_219_n1904) );
  OAI21_X1 DP_mult_219_U1565 ( .B1(DP_mult_219_n1584), .B2(DP_mult_219_n1585), 
        .A(DP_mult_219_n1615), .ZN(DP_mult_219_n1903) );
  OAI221_X1 DP_mult_219_U1564 ( .B1(DP_mult_219_n1617), .B2(DP_mult_219_n1587), 
        .C1(DP_mult_219_n1620), .C2(DP_mult_219_n1583), .A(DP_mult_219_n1903), 
        .ZN(DP_mult_219_n1902) );
  XNOR2_X1 DP_mult_219_U1563 ( .A(DP_coeff_pipe03[14]), .B(DP_mult_219_n1902), 
        .ZN(DP_mult_219_n801) );
  OAI22_X1 DP_mult_219_U1562 ( .A1(DP_mult_219_n1633), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1634), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1901)
         );
  AOI221_X1 DP_mult_219_U1561 ( .B1(DP_mult_219_n1584), .B2(DP_mult_219_n1615), 
        .C1(DP_mult_219_n1585), .C2(DP_mult_219_n1615), .A(DP_mult_219_n1901), 
        .ZN(DP_mult_219_n1900) );
  XNOR2_X1 DP_mult_219_U1560 ( .A(DP_coeff_pipe03[14]), .B(DP_mult_219_n1900), 
        .ZN(DP_mult_219_n802) );
  OAI22_X1 DP_mult_219_U1559 ( .A1(DP_mult_219_n1617), .A2(DP_mult_219_n1533), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1899)
         );
  AOI221_X1 DP_mult_219_U1558 ( .B1(DP_mult_219_n1585), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1536), .C2(DP_mult_219_n1375), .A(DP_mult_219_n1899), 
        .ZN(DP_mult_219_n1898) );
  XNOR2_X1 DP_mult_219_U1557 ( .A(DP_coeff_pipe03[14]), .B(DP_mult_219_n1898), 
        .ZN(DP_mult_219_n803) );
  OAI22_X1 DP_mult_219_U1556 ( .A1(DP_mult_219_n1640), .A2(DP_mult_219_n1587), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1539), .ZN(DP_mult_219_n1897)
         );
  AOI221_X1 DP_mult_219_U1555 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1536), .C2(DP_mult_219_n1376), .A(DP_mult_219_n1897), 
        .ZN(DP_mult_219_n1896) );
  XNOR2_X1 DP_mult_219_U1554 ( .A(DP_coeff_pipe03[14]), .B(DP_mult_219_n1896), 
        .ZN(DP_mult_219_n804) );
  OAI22_X1 DP_mult_219_U1553 ( .A1(DP_mult_219_n1728), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1729), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1895)
         );
  AOI221_X1 DP_mult_219_U1552 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[21]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[20]), .A(DP_mult_219_n1895), 
        .ZN(DP_mult_219_n1894) );
  XNOR2_X1 DP_mult_219_U1551 ( .A(DP_coeff_pipe03[14]), .B(DP_mult_219_n1894), 
        .ZN(DP_mult_219_n805) );
  OAI22_X1 DP_mult_219_U1550 ( .A1(DP_mult_219_n1724), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1725), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1893)
         );
  AOI221_X1 DP_mult_219_U1549 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[20]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[19]), .A(DP_mult_219_n1893), 
        .ZN(DP_mult_219_n1892) );
  XNOR2_X1 DP_mult_219_U1548 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1892), 
        .ZN(DP_mult_219_n806) );
  OAI22_X1 DP_mult_219_U1547 ( .A1(DP_mult_219_n1720), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1721), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1891)
         );
  AOI221_X1 DP_mult_219_U1546 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[19]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[18]), .A(DP_mult_219_n1891), 
        .ZN(DP_mult_219_n1890) );
  XNOR2_X1 DP_mult_219_U1545 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1890), 
        .ZN(DP_mult_219_n807) );
  OAI22_X1 DP_mult_219_U1544 ( .A1(DP_mult_219_n1716), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1717), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1889)
         );
  AOI221_X1 DP_mult_219_U1543 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[18]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[17]), .A(DP_mult_219_n1889), 
        .ZN(DP_mult_219_n1888) );
  XNOR2_X1 DP_mult_219_U1542 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1888), 
        .ZN(DP_mult_219_n808) );
  OAI22_X1 DP_mult_219_U1541 ( .A1(DP_mult_219_n1712), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1713), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1887)
         );
  AOI221_X1 DP_mult_219_U1540 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[17]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[16]), .A(DP_mult_219_n1887), 
        .ZN(DP_mult_219_n1886) );
  XNOR2_X1 DP_mult_219_U1539 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1886), 
        .ZN(DP_mult_219_n809) );
  OAI22_X1 DP_mult_219_U1538 ( .A1(DP_mult_219_n1708), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1709), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1885)
         );
  AOI221_X1 DP_mult_219_U1537 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[16]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[15]), .A(DP_mult_219_n1885), 
        .ZN(DP_mult_219_n1884) );
  XNOR2_X1 DP_mult_219_U1536 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1884), 
        .ZN(DP_mult_219_n810) );
  OAI22_X1 DP_mult_219_U1535 ( .A1(DP_mult_219_n1704), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1705), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1883)
         );
  AOI221_X1 DP_mult_219_U1534 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[15]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[14]), .A(DP_mult_219_n1883), 
        .ZN(DP_mult_219_n1882) );
  XNOR2_X1 DP_mult_219_U1533 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1882), 
        .ZN(DP_mult_219_n811) );
  OAI22_X1 DP_mult_219_U1532 ( .A1(DP_mult_219_n1700), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1701), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1881)
         );
  AOI221_X1 DP_mult_219_U1531 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[14]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[13]), .A(DP_mult_219_n1881), 
        .ZN(DP_mult_219_n1880) );
  XNOR2_X1 DP_mult_219_U1530 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1880), 
        .ZN(DP_mult_219_n812) );
  OAI22_X1 DP_mult_219_U1529 ( .A1(DP_mult_219_n1696), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1697), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1879)
         );
  AOI221_X1 DP_mult_219_U1528 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[13]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[12]), .A(DP_mult_219_n1879), 
        .ZN(DP_mult_219_n1878) );
  XNOR2_X1 DP_mult_219_U1527 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1878), 
        .ZN(DP_mult_219_n813) );
  OAI22_X1 DP_mult_219_U1526 ( .A1(DP_mult_219_n1692), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1693), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1877)
         );
  AOI221_X1 DP_mult_219_U1525 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[12]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[11]), .A(DP_mult_219_n1877), 
        .ZN(DP_mult_219_n1876) );
  XNOR2_X1 DP_mult_219_U1524 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1876), 
        .ZN(DP_mult_219_n814) );
  OAI22_X1 DP_mult_219_U1523 ( .A1(DP_mult_219_n1688), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1689), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1875)
         );
  AOI221_X1 DP_mult_219_U1522 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[11]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[10]), .A(DP_mult_219_n1875), 
        .ZN(DP_mult_219_n1874) );
  XNOR2_X1 DP_mult_219_U1521 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1874), 
        .ZN(DP_mult_219_n815) );
  OAI22_X1 DP_mult_219_U1520 ( .A1(DP_mult_219_n1684), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1685), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1873)
         );
  AOI221_X1 DP_mult_219_U1519 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[10]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[9]), .A(DP_mult_219_n1873), .ZN(
        DP_mult_219_n1872) );
  XNOR2_X1 DP_mult_219_U1518 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1872), 
        .ZN(DP_mult_219_n816) );
  OAI22_X1 DP_mult_219_U1517 ( .A1(DP_mult_219_n1680), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1681), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1871)
         );
  AOI221_X1 DP_mult_219_U1516 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[9]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[8]), .A(DP_mult_219_n1871), .ZN(
        DP_mult_219_n1870) );
  XNOR2_X1 DP_mult_219_U1515 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1870), 
        .ZN(DP_mult_219_n817) );
  OAI22_X1 DP_mult_219_U1514 ( .A1(DP_mult_219_n1676), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1677), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1869)
         );
  AOI221_X1 DP_mult_219_U1513 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[8]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[7]), .A(DP_mult_219_n1869), .ZN(
        DP_mult_219_n1868) );
  XNOR2_X1 DP_mult_219_U1512 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1868), 
        .ZN(DP_mult_219_n818) );
  OAI22_X1 DP_mult_219_U1511 ( .A1(DP_mult_219_n1672), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1673), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1867)
         );
  AOI221_X1 DP_mult_219_U1510 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[7]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[6]), .A(DP_mult_219_n1867), .ZN(
        DP_mult_219_n1866) );
  XNOR2_X1 DP_mult_219_U1509 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1866), 
        .ZN(DP_mult_219_n819) );
  OAI22_X1 DP_mult_219_U1508 ( .A1(DP_mult_219_n1668), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1669), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1865)
         );
  AOI221_X1 DP_mult_219_U1507 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[6]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[5]), .A(DP_mult_219_n1865), .ZN(
        DP_mult_219_n1864) );
  XNOR2_X1 DP_mult_219_U1506 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1864), 
        .ZN(DP_mult_219_n820) );
  OAI22_X1 DP_mult_219_U1505 ( .A1(DP_mult_219_n1664), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1665), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1863)
         );
  AOI221_X1 DP_mult_219_U1504 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[5]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[4]), .A(DP_mult_219_n1863), .ZN(
        DP_mult_219_n1862) );
  XNOR2_X1 DP_mult_219_U1503 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1862), 
        .ZN(DP_mult_219_n821) );
  OAI22_X1 DP_mult_219_U1502 ( .A1(DP_mult_219_n1660), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1661), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1861)
         );
  AOI221_X1 DP_mult_219_U1501 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[4]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[3]), .A(DP_mult_219_n1861), .ZN(
        DP_mult_219_n1860) );
  XNOR2_X1 DP_mult_219_U1500 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1860), 
        .ZN(DP_mult_219_n822) );
  OAI22_X1 DP_mult_219_U1499 ( .A1(DP_mult_219_n1657), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1649), .B2(DP_mult_219_n1587), .ZN(DP_mult_219_n1859)
         );
  AOI221_X1 DP_mult_219_U1498 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[3]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[2]), .A(DP_mult_219_n1859), .ZN(
        DP_mult_219_n1858) );
  XNOR2_X1 DP_mult_219_U1497 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1858), 
        .ZN(DP_mult_219_n823) );
  OAI22_X1 DP_mult_219_U1496 ( .A1(DP_mult_219_n1653), .A2(DP_mult_219_n1583), 
        .B1(DP_mult_219_n1565), .B2(DP_mult_219_n1586), .ZN(DP_mult_219_n1856)
         );
  AOI221_X1 DP_mult_219_U1495 ( .B1(DP_mult_219_n1584), .B2(DP_pipe03[2]), 
        .C1(DP_mult_219_n1585), .C2(DP_pipe03[1]), .A(DP_mult_219_n1856), .ZN(
        DP_mult_219_n1855) );
  XNOR2_X1 DP_mult_219_U1494 ( .A(DP_mult_219_n1604), .B(DP_mult_219_n1855), 
        .ZN(DP_mult_219_n824) );
  OAI222_X1 DP_mult_219_U1493 ( .A1(DP_mult_219_n1649), .A2(DP_mult_219_n1533), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1539), .C1(DP_mult_219_n1650), 
        .C2(DP_mult_219_n1583), .ZN(DP_mult_219_n1854) );
  XNOR2_X1 DP_mult_219_U1492 ( .A(DP_mult_219_n1854), .B(DP_mult_219_n1605), 
        .ZN(DP_mult_219_n825) );
  OAI22_X1 DP_mult_219_U1491 ( .A1(DP_mult_219_n1565), .A2(DP_mult_219_n1533), 
        .B1(DP_mult_219_n1565), .B2(DP_mult_219_n1583), .ZN(DP_mult_219_n1853)
         );
  XNOR2_X1 DP_mult_219_U1490 ( .A(DP_mult_219_n1853), .B(DP_mult_219_n1605), 
        .ZN(DP_mult_219_n826) );
  XOR2_X1 DP_mult_219_U1489 ( .A(DP_coeff_pipe03[9]), .B(DP_mult_219_n1601), 
        .Z(DP_mult_219_n1852) );
  XNOR2_X1 DP_mult_219_U1488 ( .A(DP_coeff_pipe03[10]), .B(DP_mult_219_n1603), 
        .ZN(DP_mult_219_n1851) );
  XNOR2_X1 DP_mult_219_U1487 ( .A(DP_coeff_pipe03[10]), .B(DP_coeff_pipe03[9]), 
        .ZN(DP_mult_219_n1850) );
  NAND3_X1 DP_mult_219_U1486 ( .A1(DP_mult_219_n1852), .A2(DP_mult_219_n1851), 
        .A3(DP_mult_219_n1850), .ZN(DP_mult_219_n1802) );
  INV_X1 DP_mult_219_U1485 ( .A(DP_mult_219_n1852), .ZN(DP_mult_219_n1849) );
  OAI21_X1 DP_mult_219_U1484 ( .B1(DP_mult_219_n1579), .B2(DP_mult_219_n1580), 
        .A(DP_mult_219_n1615), .ZN(DP_mult_219_n1848) );
  OAI221_X1 DP_mult_219_U1483 ( .B1(DP_mult_219_n1618), .B2(DP_mult_219_n1582), 
        .C1(DP_mult_219_n1617), .C2(DP_mult_219_n1578), .A(DP_mult_219_n1848), 
        .ZN(DP_mult_219_n1847) );
  XNOR2_X1 DP_mult_219_U1482 ( .A(DP_coeff_pipe03[11]), .B(DP_mult_219_n1847), 
        .ZN(DP_mult_219_n827) );
  OAI22_X1 DP_mult_219_U1481 ( .A1(DP_mult_219_n1633), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1634), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1846)
         );
  AOI221_X1 DP_mult_219_U1480 ( .B1(DP_mult_219_n1579), .B2(DP_mult_219_n1615), 
        .C1(DP_mult_219_n1580), .C2(DP_mult_219_n1615), .A(DP_mult_219_n1846), 
        .ZN(DP_mult_219_n1845) );
  XNOR2_X1 DP_mult_219_U1479 ( .A(DP_coeff_pipe03[11]), .B(DP_mult_219_n1845), 
        .ZN(DP_mult_219_n828) );
  OAI22_X1 DP_mult_219_U1478 ( .A1(DP_mult_219_n1617), .A2(DP_mult_219_n1545), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1844)
         );
  AOI221_X1 DP_mult_219_U1477 ( .B1(DP_mult_219_n1580), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1535), .C2(DP_mult_219_n1375), .A(DP_mult_219_n1844), 
        .ZN(DP_mult_219_n1843) );
  XNOR2_X1 DP_mult_219_U1476 ( .A(DP_coeff_pipe03[11]), .B(DP_mult_219_n1843), 
        .ZN(DP_mult_219_n829) );
  OAI22_X1 DP_mult_219_U1475 ( .A1(DP_mult_219_n1640), .A2(DP_mult_219_n1582), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1538), .ZN(DP_mult_219_n1842)
         );
  AOI221_X1 DP_mult_219_U1474 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1535), .C2(DP_mult_219_n1376), .A(DP_mult_219_n1842), 
        .ZN(DP_mult_219_n1841) );
  XNOR2_X1 DP_mult_219_U1473 ( .A(DP_coeff_pipe03[11]), .B(DP_mult_219_n1841), 
        .ZN(DP_mult_219_n830) );
  OAI22_X1 DP_mult_219_U1472 ( .A1(DP_mult_219_n1728), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1729), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1840)
         );
  AOI221_X1 DP_mult_219_U1471 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[21]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[20]), .A(DP_mult_219_n1840), 
        .ZN(DP_mult_219_n1839) );
  XNOR2_X1 DP_mult_219_U1470 ( .A(DP_coeff_pipe03[11]), .B(DP_mult_219_n1839), 
        .ZN(DP_mult_219_n831) );
  OAI22_X1 DP_mult_219_U1469 ( .A1(DP_mult_219_n1724), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1725), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1838)
         );
  AOI221_X1 DP_mult_219_U1468 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[20]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[19]), .A(DP_mult_219_n1838), 
        .ZN(DP_mult_219_n1837) );
  XNOR2_X1 DP_mult_219_U1467 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1837), 
        .ZN(DP_mult_219_n832) );
  OAI22_X1 DP_mult_219_U1466 ( .A1(DP_mult_219_n1720), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1721), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1836)
         );
  AOI221_X1 DP_mult_219_U1465 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[19]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[18]), .A(DP_mult_219_n1836), 
        .ZN(DP_mult_219_n1835) );
  XNOR2_X1 DP_mult_219_U1464 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1835), 
        .ZN(DP_mult_219_n833) );
  OAI22_X1 DP_mult_219_U1463 ( .A1(DP_mult_219_n1716), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1717), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1834)
         );
  AOI221_X1 DP_mult_219_U1462 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[18]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[17]), .A(DP_mult_219_n1834), 
        .ZN(DP_mult_219_n1833) );
  XNOR2_X1 DP_mult_219_U1461 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1833), 
        .ZN(DP_mult_219_n834) );
  OAI22_X1 DP_mult_219_U1460 ( .A1(DP_mult_219_n1712), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1713), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1832)
         );
  AOI221_X1 DP_mult_219_U1459 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[17]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[16]), .A(DP_mult_219_n1832), 
        .ZN(DP_mult_219_n1831) );
  XNOR2_X1 DP_mult_219_U1458 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1831), 
        .ZN(DP_mult_219_n835) );
  OAI22_X1 DP_mult_219_U1457 ( .A1(DP_mult_219_n1708), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1709), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1830)
         );
  AOI221_X1 DP_mult_219_U1456 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[16]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[15]), .A(DP_mult_219_n1830), 
        .ZN(DP_mult_219_n1829) );
  XNOR2_X1 DP_mult_219_U1455 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1829), 
        .ZN(DP_mult_219_n836) );
  OAI22_X1 DP_mult_219_U1454 ( .A1(DP_mult_219_n1704), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1705), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1828)
         );
  AOI221_X1 DP_mult_219_U1453 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[15]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[14]), .A(DP_mult_219_n1828), 
        .ZN(DP_mult_219_n1827) );
  XNOR2_X1 DP_mult_219_U1452 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1827), 
        .ZN(DP_mult_219_n837) );
  OAI22_X1 DP_mult_219_U1451 ( .A1(DP_mult_219_n1700), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1701), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1826)
         );
  AOI221_X1 DP_mult_219_U1450 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[14]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[13]), .A(DP_mult_219_n1826), 
        .ZN(DP_mult_219_n1825) );
  XNOR2_X1 DP_mult_219_U1449 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1825), 
        .ZN(DP_mult_219_n838) );
  OAI22_X1 DP_mult_219_U1448 ( .A1(DP_mult_219_n1696), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1697), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1824)
         );
  AOI221_X1 DP_mult_219_U1447 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[13]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[12]), .A(DP_mult_219_n1824), 
        .ZN(DP_mult_219_n1823) );
  XNOR2_X1 DP_mult_219_U1446 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1823), 
        .ZN(DP_mult_219_n839) );
  OAI22_X1 DP_mult_219_U1445 ( .A1(DP_mult_219_n1692), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1693), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1822)
         );
  AOI221_X1 DP_mult_219_U1444 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[12]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[11]), .A(DP_mult_219_n1822), 
        .ZN(DP_mult_219_n1821) );
  XNOR2_X1 DP_mult_219_U1443 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1821), 
        .ZN(DP_mult_219_n840) );
  OAI22_X1 DP_mult_219_U1442 ( .A1(DP_mult_219_n1688), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1689), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1820)
         );
  AOI221_X1 DP_mult_219_U1441 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[11]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[10]), .A(DP_mult_219_n1820), 
        .ZN(DP_mult_219_n1819) );
  XNOR2_X1 DP_mult_219_U1440 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1819), 
        .ZN(DP_mult_219_n841) );
  OAI22_X1 DP_mult_219_U1439 ( .A1(DP_mult_219_n1684), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1685), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1818)
         );
  AOI221_X1 DP_mult_219_U1438 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[10]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[9]), .A(DP_mult_219_n1818), .ZN(
        DP_mult_219_n1817) );
  XNOR2_X1 DP_mult_219_U1437 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1817), 
        .ZN(DP_mult_219_n842) );
  OAI22_X1 DP_mult_219_U1436 ( .A1(DP_mult_219_n1680), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1681), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1816)
         );
  AOI221_X1 DP_mult_219_U1435 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[9]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[8]), .A(DP_mult_219_n1816), .ZN(
        DP_mult_219_n1815) );
  XNOR2_X1 DP_mult_219_U1434 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1815), 
        .ZN(DP_mult_219_n843) );
  OAI22_X1 DP_mult_219_U1433 ( .A1(DP_mult_219_n1676), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1677), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1814)
         );
  AOI221_X1 DP_mult_219_U1432 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[8]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[7]), .A(DP_mult_219_n1814), .ZN(
        DP_mult_219_n1813) );
  XNOR2_X1 DP_mult_219_U1431 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1813), 
        .ZN(DP_mult_219_n844) );
  OAI22_X1 DP_mult_219_U1430 ( .A1(DP_mult_219_n1672), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1673), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1812)
         );
  AOI221_X1 DP_mult_219_U1429 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[7]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[6]), .A(DP_mult_219_n1812), .ZN(
        DP_mult_219_n1811) );
  XNOR2_X1 DP_mult_219_U1428 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1811), 
        .ZN(DP_mult_219_n845) );
  OAI22_X1 DP_mult_219_U1427 ( .A1(DP_mult_219_n1668), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1669), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1810)
         );
  AOI221_X1 DP_mult_219_U1426 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[6]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[5]), .A(DP_mult_219_n1810), .ZN(
        DP_mult_219_n1809) );
  XNOR2_X1 DP_mult_219_U1425 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1809), 
        .ZN(DP_mult_219_n846) );
  OAI22_X1 DP_mult_219_U1424 ( .A1(DP_mult_219_n1664), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1665), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1808)
         );
  AOI221_X1 DP_mult_219_U1423 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[5]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[4]), .A(DP_mult_219_n1808), .ZN(
        DP_mult_219_n1807) );
  XNOR2_X1 DP_mult_219_U1422 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1807), 
        .ZN(DP_mult_219_n847) );
  OAI22_X1 DP_mult_219_U1421 ( .A1(DP_mult_219_n1660), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1661), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1806)
         );
  AOI221_X1 DP_mult_219_U1420 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[4]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[3]), .A(DP_mult_219_n1806), .ZN(
        DP_mult_219_n1805) );
  XNOR2_X1 DP_mult_219_U1419 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1805), 
        .ZN(DP_mult_219_n848) );
  OAI22_X1 DP_mult_219_U1418 ( .A1(DP_mult_219_n1657), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1649), .B2(DP_mult_219_n1582), .ZN(DP_mult_219_n1804)
         );
  AOI221_X1 DP_mult_219_U1417 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[3]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[2]), .A(DP_mult_219_n1804), .ZN(
        DP_mult_219_n1803) );
  XNOR2_X1 DP_mult_219_U1416 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1803), 
        .ZN(DP_mult_219_n849) );
  OAI22_X1 DP_mult_219_U1415 ( .A1(DP_mult_219_n1653), .A2(DP_mult_219_n1578), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1581), .ZN(DP_mult_219_n1801)
         );
  AOI221_X1 DP_mult_219_U1414 ( .B1(DP_mult_219_n1579), .B2(DP_pipe03[2]), 
        .C1(DP_mult_219_n1580), .C2(DP_pipe03[1]), .A(DP_mult_219_n1801), .ZN(
        DP_mult_219_n1800) );
  XNOR2_X1 DP_mult_219_U1413 ( .A(DP_mult_219_n1602), .B(DP_mult_219_n1800), 
        .ZN(DP_mult_219_n850) );
  OAI222_X1 DP_mult_219_U1412 ( .A1(DP_mult_219_n1649), .A2(DP_mult_219_n1545), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1538), .C1(DP_mult_219_n1650), 
        .C2(DP_mult_219_n1578), .ZN(DP_mult_219_n1799) );
  XNOR2_X1 DP_mult_219_U1411 ( .A(DP_mult_219_n1799), .B(DP_mult_219_n1603), 
        .ZN(DP_mult_219_n851) );
  OAI22_X1 DP_mult_219_U1410 ( .A1(DP_mult_219_n1565), .A2(DP_mult_219_n1545), 
        .B1(DP_mult_219_n1565), .B2(DP_mult_219_n1578), .ZN(DP_mult_219_n1798)
         );
  XNOR2_X1 DP_mult_219_U1409 ( .A(DP_mult_219_n1798), .B(DP_mult_219_n1603), 
        .ZN(DP_mult_219_n852) );
  XOR2_X1 DP_mult_219_U1408 ( .A(DP_coeff_pipe03[6]), .B(DP_mult_219_n1599), 
        .Z(DP_mult_219_n1797) );
  XNOR2_X1 DP_mult_219_U1407 ( .A(DP_coeff_pipe03[7]), .B(DP_mult_219_n1601), 
        .ZN(DP_mult_219_n1796) );
  XNOR2_X1 DP_mult_219_U1406 ( .A(DP_coeff_pipe03[6]), .B(DP_coeff_pipe03[7]), 
        .ZN(DP_mult_219_n1795) );
  NAND3_X1 DP_mult_219_U1405 ( .A1(DP_mult_219_n1797), .A2(DP_mult_219_n1796), 
        .A3(DP_mult_219_n1795), .ZN(DP_mult_219_n1747) );
  INV_X1 DP_mult_219_U1404 ( .A(DP_mult_219_n1797), .ZN(DP_mult_219_n1794) );
  OAI21_X1 DP_mult_219_U1403 ( .B1(DP_mult_219_n1574), .B2(DP_mult_219_n1575), 
        .A(DP_mult_219_n1615), .ZN(DP_mult_219_n1793) );
  OAI221_X1 DP_mult_219_U1402 ( .B1(DP_mult_219_n1618), .B2(DP_mult_219_n1577), 
        .C1(DP_mult_219_n1617), .C2(DP_mult_219_n1573), .A(DP_mult_219_n1793), 
        .ZN(DP_mult_219_n1792) );
  XNOR2_X1 DP_mult_219_U1401 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1792), 
        .ZN(DP_mult_219_n853) );
  OAI22_X1 DP_mult_219_U1400 ( .A1(DP_mult_219_n1633), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1634), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1791)
         );
  AOI221_X1 DP_mult_219_U1399 ( .B1(DP_mult_219_n1574), .B2(DP_mult_219_n1614), 
        .C1(DP_mult_219_n1575), .C2(DP_mult_219_n1615), .A(DP_mult_219_n1791), 
        .ZN(DP_mult_219_n1790) );
  XNOR2_X1 DP_mult_219_U1398 ( .A(DP_coeff_pipe03[8]), .B(DP_mult_219_n1790), 
        .ZN(DP_mult_219_n854) );
  OAI22_X1 DP_mult_219_U1397 ( .A1(DP_mult_219_n1617), .A2(DP_mult_219_n1544), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1789)
         );
  AOI221_X1 DP_mult_219_U1396 ( .B1(DP_mult_219_n1575), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1546), .C2(DP_mult_219_n1375), .A(DP_mult_219_n1789), 
        .ZN(DP_mult_219_n1788) );
  XNOR2_X1 DP_mult_219_U1395 ( .A(DP_coeff_pipe03[8]), .B(DP_mult_219_n1788), 
        .ZN(DP_mult_219_n855) );
  OAI22_X1 DP_mult_219_U1394 ( .A1(DP_mult_219_n1640), .A2(DP_mult_219_n1577), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1547), .ZN(DP_mult_219_n1787)
         );
  AOI221_X1 DP_mult_219_U1393 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1546), .C2(DP_mult_219_n1376), .A(DP_mult_219_n1787), 
        .ZN(DP_mult_219_n1786) );
  XNOR2_X1 DP_mult_219_U1392 ( .A(DP_coeff_pipe03[8]), .B(DP_mult_219_n1786), 
        .ZN(DP_mult_219_n856) );
  OAI22_X1 DP_mult_219_U1391 ( .A1(DP_mult_219_n1728), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1729), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1785)
         );
  AOI221_X1 DP_mult_219_U1390 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[21]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[20]), .A(DP_mult_219_n1785), 
        .ZN(DP_mult_219_n1784) );
  XNOR2_X1 DP_mult_219_U1389 ( .A(DP_coeff_pipe03[8]), .B(DP_mult_219_n1784), 
        .ZN(DP_mult_219_n857) );
  OAI22_X1 DP_mult_219_U1388 ( .A1(DP_mult_219_n1724), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1725), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1783)
         );
  AOI221_X1 DP_mult_219_U1387 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[20]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[19]), .A(DP_mult_219_n1783), 
        .ZN(DP_mult_219_n1782) );
  XNOR2_X1 DP_mult_219_U1386 ( .A(DP_coeff_pipe03[8]), .B(DP_mult_219_n1782), 
        .ZN(DP_mult_219_n858) );
  OAI22_X1 DP_mult_219_U1385 ( .A1(DP_mult_219_n1720), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1721), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1781)
         );
  AOI221_X1 DP_mult_219_U1384 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[19]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[18]), .A(DP_mult_219_n1781), 
        .ZN(DP_mult_219_n1780) );
  XNOR2_X1 DP_mult_219_U1383 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1780), 
        .ZN(DP_mult_219_n859) );
  OAI22_X1 DP_mult_219_U1382 ( .A1(DP_mult_219_n1716), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1717), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1779)
         );
  AOI221_X1 DP_mult_219_U1381 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[18]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[17]), .A(DP_mult_219_n1779), 
        .ZN(DP_mult_219_n1778) );
  XNOR2_X1 DP_mult_219_U1380 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1778), 
        .ZN(DP_mult_219_n860) );
  OAI22_X1 DP_mult_219_U1379 ( .A1(DP_mult_219_n1712), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1713), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1777)
         );
  AOI221_X1 DP_mult_219_U1378 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[17]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[16]), .A(DP_mult_219_n1777), 
        .ZN(DP_mult_219_n1776) );
  XNOR2_X1 DP_mult_219_U1377 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1776), 
        .ZN(DP_mult_219_n861) );
  OAI22_X1 DP_mult_219_U1376 ( .A1(DP_mult_219_n1708), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1709), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1775)
         );
  AOI221_X1 DP_mult_219_U1375 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[16]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[15]), .A(DP_mult_219_n1775), 
        .ZN(DP_mult_219_n1774) );
  XNOR2_X1 DP_mult_219_U1374 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1774), 
        .ZN(DP_mult_219_n862) );
  OAI22_X1 DP_mult_219_U1373 ( .A1(DP_mult_219_n1704), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1705), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1773)
         );
  AOI221_X1 DP_mult_219_U1372 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[15]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[14]), .A(DP_mult_219_n1773), 
        .ZN(DP_mult_219_n1772) );
  XNOR2_X1 DP_mult_219_U1371 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1772), 
        .ZN(DP_mult_219_n863) );
  OAI22_X1 DP_mult_219_U1370 ( .A1(DP_mult_219_n1700), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1701), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1771)
         );
  AOI221_X1 DP_mult_219_U1369 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[14]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[13]), .A(DP_mult_219_n1771), 
        .ZN(DP_mult_219_n1770) );
  XNOR2_X1 DP_mult_219_U1368 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1770), 
        .ZN(DP_mult_219_n864) );
  OAI22_X1 DP_mult_219_U1367 ( .A1(DP_mult_219_n1696), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1697), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1769)
         );
  AOI221_X1 DP_mult_219_U1366 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[13]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[12]), .A(DP_mult_219_n1769), 
        .ZN(DP_mult_219_n1768) );
  XNOR2_X1 DP_mult_219_U1365 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1768), 
        .ZN(DP_mult_219_n865) );
  OAI22_X1 DP_mult_219_U1364 ( .A1(DP_mult_219_n1692), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1693), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1767)
         );
  AOI221_X1 DP_mult_219_U1363 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[12]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[11]), .A(DP_mult_219_n1767), 
        .ZN(DP_mult_219_n1766) );
  XNOR2_X1 DP_mult_219_U1362 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1766), 
        .ZN(DP_mult_219_n866) );
  OAI22_X1 DP_mult_219_U1361 ( .A1(DP_mult_219_n1688), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1689), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1765)
         );
  AOI221_X1 DP_mult_219_U1360 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[11]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[10]), .A(DP_mult_219_n1765), 
        .ZN(DP_mult_219_n1764) );
  XNOR2_X1 DP_mult_219_U1359 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1764), 
        .ZN(DP_mult_219_n867) );
  OAI22_X1 DP_mult_219_U1358 ( .A1(DP_mult_219_n1684), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1685), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1763)
         );
  AOI221_X1 DP_mult_219_U1357 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[10]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[9]), .A(DP_mult_219_n1763), .ZN(
        DP_mult_219_n1762) );
  XNOR2_X1 DP_mult_219_U1356 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1762), 
        .ZN(DP_mult_219_n868) );
  OAI22_X1 DP_mult_219_U1355 ( .A1(DP_mult_219_n1680), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1681), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1761)
         );
  AOI221_X1 DP_mult_219_U1354 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[9]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[8]), .A(DP_mult_219_n1761), .ZN(
        DP_mult_219_n1760) );
  XNOR2_X1 DP_mult_219_U1353 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1760), 
        .ZN(DP_mult_219_n869) );
  OAI22_X1 DP_mult_219_U1352 ( .A1(DP_mult_219_n1676), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1677), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1759)
         );
  AOI221_X1 DP_mult_219_U1351 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[8]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[7]), .A(DP_mult_219_n1759), .ZN(
        DP_mult_219_n1758) );
  XNOR2_X1 DP_mult_219_U1350 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1758), 
        .ZN(DP_mult_219_n870) );
  OAI22_X1 DP_mult_219_U1349 ( .A1(DP_mult_219_n1672), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1673), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1757)
         );
  AOI221_X1 DP_mult_219_U1348 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[7]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[6]), .A(DP_mult_219_n1757), .ZN(
        DP_mult_219_n1756) );
  XNOR2_X1 DP_mult_219_U1347 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1756), 
        .ZN(DP_mult_219_n871) );
  OAI22_X1 DP_mult_219_U1346 ( .A1(DP_mult_219_n1668), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1669), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1755)
         );
  AOI221_X1 DP_mult_219_U1345 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[6]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[5]), .A(DP_mult_219_n1755), .ZN(
        DP_mult_219_n1754) );
  XNOR2_X1 DP_mult_219_U1344 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1754), 
        .ZN(DP_mult_219_n872) );
  OAI22_X1 DP_mult_219_U1343 ( .A1(DP_mult_219_n1664), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1665), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1753)
         );
  AOI221_X1 DP_mult_219_U1342 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[5]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[4]), .A(DP_mult_219_n1753), .ZN(
        DP_mult_219_n1752) );
  XNOR2_X1 DP_mult_219_U1341 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1752), 
        .ZN(DP_mult_219_n873) );
  OAI22_X1 DP_mult_219_U1340 ( .A1(DP_mult_219_n1660), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1661), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1751)
         );
  AOI221_X1 DP_mult_219_U1339 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[4]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[3]), .A(DP_mult_219_n1751), .ZN(
        DP_mult_219_n1750) );
  XNOR2_X1 DP_mult_219_U1338 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1750), 
        .ZN(DP_mult_219_n874) );
  OAI22_X1 DP_mult_219_U1337 ( .A1(DP_mult_219_n1657), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1649), .B2(DP_mult_219_n1577), .ZN(DP_mult_219_n1749)
         );
  AOI221_X1 DP_mult_219_U1336 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[3]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[2]), .A(DP_mult_219_n1749), .ZN(
        DP_mult_219_n1748) );
  XNOR2_X1 DP_mult_219_U1335 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1748), 
        .ZN(DP_mult_219_n875) );
  OAI22_X1 DP_mult_219_U1334 ( .A1(DP_mult_219_n1653), .A2(DP_mult_219_n1573), 
        .B1(DP_mult_219_n1565), .B2(DP_mult_219_n1576), .ZN(DP_mult_219_n1746)
         );
  AOI221_X1 DP_mult_219_U1333 ( .B1(DP_mult_219_n1574), .B2(DP_pipe03[2]), 
        .C1(DP_mult_219_n1575), .C2(DP_pipe03[1]), .A(DP_mult_219_n1746), .ZN(
        DP_mult_219_n1745) );
  XNOR2_X1 DP_mult_219_U1332 ( .A(DP_mult_219_n1600), .B(DP_mult_219_n1745), 
        .ZN(DP_mult_219_n876) );
  OAI222_X1 DP_mult_219_U1331 ( .A1(DP_mult_219_n1649), .A2(DP_mult_219_n1544), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1547), .C1(DP_mult_219_n1650), 
        .C2(DP_mult_219_n1573), .ZN(DP_mult_219_n1744) );
  XNOR2_X1 DP_mult_219_U1330 ( .A(DP_mult_219_n1744), .B(DP_mult_219_n1601), 
        .ZN(DP_mult_219_n877) );
  OAI22_X1 DP_mult_219_U1329 ( .A1(DP_mult_219_n1565), .A2(DP_mult_219_n1544), 
        .B1(DP_mult_219_n1565), .B2(DP_mult_219_n1573), .ZN(DP_mult_219_n1743)
         );
  XNOR2_X1 DP_mult_219_U1328 ( .A(DP_mult_219_n1743), .B(DP_mult_219_n1601), 
        .ZN(DP_mult_219_n878) );
  XOR2_X1 DP_mult_219_U1327 ( .A(DP_coeff_pipe03[3]), .B(DP_mult_219_n1742), 
        .Z(DP_mult_219_n1741) );
  XNOR2_X1 DP_mult_219_U1326 ( .A(DP_coeff_pipe03[4]), .B(DP_mult_219_n1599), 
        .ZN(DP_mult_219_n1740) );
  XNOR2_X1 DP_mult_219_U1325 ( .A(DP_coeff_pipe03[3]), .B(DP_coeff_pipe03[4]), 
        .ZN(DP_mult_219_n1739) );
  NAND3_X1 DP_mult_219_U1324 ( .A1(DP_mult_219_n1741), .A2(DP_mult_219_n1740), 
        .A3(DP_mult_219_n1739), .ZN(DP_mult_219_n1654) );
  INV_X1 DP_mult_219_U1323 ( .A(DP_mult_219_n1741), .ZN(DP_mult_219_n1738) );
  OAI21_X1 DP_mult_219_U1322 ( .B1(DP_mult_219_n1569), .B2(DP_mult_219_n1570), 
        .A(DP_mult_219_n1615), .ZN(DP_mult_219_n1737) );
  OAI221_X1 DP_mult_219_U1321 ( .B1(DP_mult_219_n1618), .B2(DP_mult_219_n1572), 
        .C1(DP_mult_219_n1618), .C2(DP_mult_219_n1568), .A(DP_mult_219_n1737), 
        .ZN(DP_mult_219_n1736) );
  XNOR2_X1 DP_mult_219_U1320 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1736), 
        .ZN(DP_mult_219_n879) );
  OAI22_X1 DP_mult_219_U1319 ( .A1(DP_mult_219_n1633), .A2(DP_mult_219_n1568), 
        .B1(DP_mult_219_n1634), .B2(DP_mult_219_n1572), .ZN(DP_mult_219_n1735)
         );
  AOI221_X1 DP_mult_219_U1318 ( .B1(DP_mult_219_n1569), .B2(DP_mult_219_n1614), 
        .C1(DP_mult_219_n1570), .C2(DP_mult_219_n1615), .A(DP_mult_219_n1735), 
        .ZN(DP_mult_219_n1734) );
  XNOR2_X1 DP_mult_219_U1317 ( .A(DP_coeff_pipe03[5]), .B(DP_mult_219_n1734), 
        .ZN(DP_mult_219_n880) );
  OAI22_X1 DP_mult_219_U1316 ( .A1(DP_mult_219_n1616), .A2(DP_mult_219_n1552), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1572), .ZN(DP_mult_219_n1733)
         );
  AOI221_X1 DP_mult_219_U1315 ( .B1(DP_mult_219_n1570), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1551), .C2(DP_mult_219_n1375), .A(DP_mult_219_n1733), 
        .ZN(DP_mult_219_n1732) );
  XNOR2_X1 DP_mult_219_U1314 ( .A(DP_coeff_pipe03[5]), .B(DP_mult_219_n1732), 
        .ZN(DP_mult_219_n881) );
  OAI22_X1 DP_mult_219_U1313 ( .A1(DP_mult_219_n1640), .A2(DP_mult_219_n1572), 
        .B1(DP_mult_219_n1643), .B2(DP_mult_219_n1553), .ZN(DP_mult_219_n1731)
         );
  AOI221_X1 DP_mult_219_U1312 ( .B1(DP_mult_219_n1569), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1551), .C2(DP_mult_219_n1376), .A(DP_mult_219_n1731), 
        .ZN(DP_mult_219_n1730) );
  XNOR2_X1 DP_mult_219_U1311 ( .A(DP_coeff_pipe03[5]), .B(DP_mult_219_n1730), 
        .ZN(DP_mult_219_n882) );
  OAI22_X1 DP_mult_219_U1310 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1728), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1729), .ZN(DP_mult_219_n1727)
         );
  AOI221_X1 DP_mult_219_U1309 ( .B1(DP_mult_219_n1569), .B2(DP_pipe03[21]), 
        .C1(DP_mult_219_n1570), .C2(DP_pipe03[20]), .A(DP_mult_219_n1727), 
        .ZN(DP_mult_219_n1726) );
  XNOR2_X1 DP_mult_219_U1308 ( .A(DP_coeff_pipe03[5]), .B(DP_mult_219_n1726), 
        .ZN(DP_mult_219_n883) );
  OAI22_X1 DP_mult_219_U1307 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1724), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1725), .ZN(DP_mult_219_n1723)
         );
  AOI221_X1 DP_mult_219_U1306 ( .B1(DP_mult_219_n1569), .B2(DP_pipe03[20]), 
        .C1(DP_pipe03[19]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1723), 
        .ZN(DP_mult_219_n1722) );
  XNOR2_X1 DP_mult_219_U1305 ( .A(DP_coeff_pipe03[5]), .B(DP_mult_219_n1722), 
        .ZN(DP_mult_219_n884) );
  OAI22_X1 DP_mult_219_U1304 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1720), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1721), .ZN(DP_mult_219_n1719)
         );
  AOI221_X1 DP_mult_219_U1303 ( .B1(DP_pipe03[19]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[18]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1719), 
        .ZN(DP_mult_219_n1718) );
  XNOR2_X1 DP_mult_219_U1302 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1718), 
        .ZN(DP_mult_219_n885) );
  OAI22_X1 DP_mult_219_U1301 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1716), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1717), .ZN(DP_mult_219_n1715)
         );
  AOI221_X1 DP_mult_219_U1300 ( .B1(DP_pipe03[18]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[17]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1715), 
        .ZN(DP_mult_219_n1714) );
  XNOR2_X1 DP_mult_219_U1299 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1714), 
        .ZN(DP_mult_219_n886) );
  OAI22_X1 DP_mult_219_U1298 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1712), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1713), .ZN(DP_mult_219_n1711)
         );
  AOI221_X1 DP_mult_219_U1297 ( .B1(DP_pipe03[17]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[16]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1711), 
        .ZN(DP_mult_219_n1710) );
  XNOR2_X1 DP_mult_219_U1296 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1710), 
        .ZN(DP_mult_219_n887) );
  OAI22_X1 DP_mult_219_U1295 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1708), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1709), .ZN(DP_mult_219_n1707)
         );
  AOI221_X1 DP_mult_219_U1294 ( .B1(DP_pipe03[16]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[15]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1707), 
        .ZN(DP_mult_219_n1706) );
  XNOR2_X1 DP_mult_219_U1293 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1706), 
        .ZN(DP_mult_219_n888) );
  OAI22_X1 DP_mult_219_U1292 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1704), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1705), .ZN(DP_mult_219_n1703)
         );
  AOI221_X1 DP_mult_219_U1291 ( .B1(DP_pipe03[15]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[14]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1703), 
        .ZN(DP_mult_219_n1702) );
  XNOR2_X1 DP_mult_219_U1290 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1702), 
        .ZN(DP_mult_219_n889) );
  OAI22_X1 DP_mult_219_U1289 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1700), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1701), .ZN(DP_mult_219_n1699)
         );
  AOI221_X1 DP_mult_219_U1288 ( .B1(DP_pipe03[14]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[13]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1699), 
        .ZN(DP_mult_219_n1698) );
  XNOR2_X1 DP_mult_219_U1287 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1698), 
        .ZN(DP_mult_219_n890) );
  OAI22_X1 DP_mult_219_U1286 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1696), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1697), .ZN(DP_mult_219_n1695)
         );
  AOI221_X1 DP_mult_219_U1285 ( .B1(DP_pipe03[13]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[12]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1695), 
        .ZN(DP_mult_219_n1694) );
  XNOR2_X1 DP_mult_219_U1284 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1694), 
        .ZN(DP_mult_219_n891) );
  OAI22_X1 DP_mult_219_U1283 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1692), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1693), .ZN(DP_mult_219_n1691)
         );
  AOI221_X1 DP_mult_219_U1282 ( .B1(DP_pipe03[12]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[11]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1691), 
        .ZN(DP_mult_219_n1690) );
  XNOR2_X1 DP_mult_219_U1281 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1690), 
        .ZN(DP_mult_219_n892) );
  OAI22_X1 DP_mult_219_U1280 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1688), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1689), .ZN(DP_mult_219_n1687)
         );
  AOI221_X1 DP_mult_219_U1279 ( .B1(DP_pipe03[11]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[10]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1687), 
        .ZN(DP_mult_219_n1686) );
  XNOR2_X1 DP_mult_219_U1278 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1686), 
        .ZN(DP_mult_219_n893) );
  OAI22_X1 DP_mult_219_U1277 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1684), 
        .B1(DP_mult_219_n1572), .B2(DP_mult_219_n1685), .ZN(DP_mult_219_n1683)
         );
  AOI221_X1 DP_mult_219_U1276 ( .B1(DP_pipe03[10]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[9]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1683), .ZN(
        DP_mult_219_n1682) );
  XNOR2_X1 DP_mult_219_U1275 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1682), 
        .ZN(DP_mult_219_n894) );
  OAI22_X1 DP_mult_219_U1274 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1680), 
        .B1(DP_mult_219_n1572), .B2(DP_mult_219_n1681), .ZN(DP_mult_219_n1679)
         );
  AOI221_X1 DP_mult_219_U1273 ( .B1(DP_pipe03[9]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[8]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1679), .ZN(
        DP_mult_219_n1678) );
  XNOR2_X1 DP_mult_219_U1272 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1678), 
        .ZN(DP_mult_219_n895) );
  OAI22_X1 DP_mult_219_U1271 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1676), 
        .B1(DP_mult_219_n1571), .B2(DP_mult_219_n1677), .ZN(DP_mult_219_n1675)
         );
  AOI221_X1 DP_mult_219_U1270 ( .B1(DP_pipe03[8]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[7]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1675), .ZN(
        DP_mult_219_n1674) );
  XNOR2_X1 DP_mult_219_U1269 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1674), 
        .ZN(DP_mult_219_n896) );
  OAI22_X1 DP_mult_219_U1268 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1672), 
        .B1(DP_mult_219_n1572), .B2(DP_mult_219_n1673), .ZN(DP_mult_219_n1671)
         );
  AOI221_X1 DP_mult_219_U1267 ( .B1(DP_pipe03[7]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[6]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1671), .ZN(
        DP_mult_219_n1670) );
  XNOR2_X1 DP_mult_219_U1266 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1670), 
        .ZN(DP_mult_219_n897) );
  OAI22_X1 DP_mult_219_U1265 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1668), 
        .B1(DP_mult_219_n1572), .B2(DP_mult_219_n1669), .ZN(DP_mult_219_n1667)
         );
  AOI221_X1 DP_mult_219_U1264 ( .B1(DP_pipe03[6]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[5]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1667), .ZN(
        DP_mult_219_n1666) );
  XNOR2_X1 DP_mult_219_U1263 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1666), 
        .ZN(DP_mult_219_n898) );
  OAI22_X1 DP_mult_219_U1262 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1664), 
        .B1(DP_mult_219_n1572), .B2(DP_mult_219_n1665), .ZN(DP_mult_219_n1663)
         );
  AOI221_X1 DP_mult_219_U1261 ( .B1(DP_pipe03[5]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[4]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1663), .ZN(
        DP_mult_219_n1662) );
  XNOR2_X1 DP_mult_219_U1260 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1662), 
        .ZN(DP_mult_219_n899) );
  OAI22_X1 DP_mult_219_U1259 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1660), 
        .B1(DP_mult_219_n1661), .B2(DP_mult_219_n1572), .ZN(DP_mult_219_n1659)
         );
  AOI221_X1 DP_mult_219_U1258 ( .B1(DP_pipe03[4]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[3]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1659), .ZN(
        DP_mult_219_n1658) );
  XNOR2_X1 DP_mult_219_U1257 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1658), 
        .ZN(DP_mult_219_n900) );
  OAI22_X1 DP_mult_219_U1256 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1657), 
        .B1(DP_mult_219_n1649), .B2(DP_mult_219_n1572), .ZN(DP_mult_219_n1656)
         );
  AOI221_X1 DP_mult_219_U1255 ( .B1(DP_pipe03[3]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[2]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1656), .ZN(
        DP_mult_219_n1655) );
  XNOR2_X1 DP_mult_219_U1254 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1655), 
        .ZN(DP_mult_219_n901) );
  OAI22_X1 DP_mult_219_U1253 ( .A1(DP_mult_219_n1568), .A2(DP_mult_219_n1653), 
        .B1(DP_mult_219_n1565), .B2(DP_mult_219_n1572), .ZN(DP_mult_219_n1652)
         );
  AOI221_X1 DP_mult_219_U1252 ( .B1(DP_pipe03[2]), .B2(DP_mult_219_n1569), 
        .C1(DP_pipe03[1]), .C2(DP_mult_219_n1570), .A(DP_mult_219_n1652), .ZN(
        DP_mult_219_n1651) );
  XNOR2_X1 DP_mult_219_U1251 ( .A(DP_mult_219_n1598), .B(DP_mult_219_n1651), 
        .ZN(DP_mult_219_n902) );
  OAI222_X1 DP_mult_219_U1250 ( .A1(DP_mult_219_n1552), .A2(DP_mult_219_n1649), 
        .B1(DP_mult_219_n1566), .B2(DP_mult_219_n1553), .C1(DP_mult_219_n1568), 
        .C2(DP_mult_219_n1650), .ZN(DP_mult_219_n1648) );
  XNOR2_X1 DP_mult_219_U1249 ( .A(DP_mult_219_n1648), .B(DP_mult_219_n1599), 
        .ZN(DP_mult_219_n903) );
  OAI22_X1 DP_mult_219_U1248 ( .A1(DP_mult_219_n1565), .A2(DP_mult_219_n1552), 
        .B1(DP_mult_219_n1568), .B2(DP_mult_219_n1567), .ZN(DP_mult_219_n1646)
         );
  XNOR2_X1 DP_mult_219_U1247 ( .A(DP_mult_219_n1646), .B(DP_mult_219_n1599), 
        .ZN(DP_mult_219_n904) );
  OAI22_X1 DP_mult_219_U1246 ( .A1(DP_mult_219_n1633), .A2(DP_mult_219_n1564), 
        .B1(DP_mult_219_n1634), .B2(DP_mult_219_n1639), .ZN(DP_mult_219_n1645)
         );
  AOI221_X1 DP_mult_219_U1245 ( .B1(DP_mult_219_n1561), .B2(DP_mult_219_n1614), 
        .C1(DP_mult_219_n1563), .C2(DP_mult_219_n1615), .A(DP_mult_219_n1645), 
        .ZN(DP_mult_219_n1644) );
  XNOR2_X1 DP_mult_219_U1244 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n1644), 
        .ZN(DP_mult_219_n906) );
  OAI22_X1 DP_mult_219_U1243 ( .A1(DP_mult_219_n1643), .A2(DP_mult_219_n1639), 
        .B1(DP_mult_219_n1617), .B2(DP_mult_219_n1554), .ZN(DP_mult_219_n1642)
         );
  AOI221_X1 DP_mult_219_U1242 ( .B1(DP_mult_219_n1563), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1555), .C2(DP_mult_219_n1375), .A(DP_mult_219_n1642), 
        .ZN(DP_mult_219_n1641) );
  XNOR2_X1 DP_mult_219_U1241 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n1641), 
        .ZN(DP_mult_219_n907) );
  INV_X1 DP_mult_219_U1240 ( .A(DP_mult_219_n1376), .ZN(DP_mult_219_n1638) );
  OAI22_X1 DP_mult_219_U1239 ( .A1(DP_mult_219_n1564), .A2(DP_mult_219_n1638), 
        .B1(DP_mult_219_n1639), .B2(DP_mult_219_n1640), .ZN(DP_mult_219_n1637)
         );
  AOI221_X1 DP_mult_219_U1238 ( .B1(DP_mult_219_n1561), .B2(DP_pipe03[22]), 
        .C1(DP_mult_219_n1563), .C2(DP_pipe03[21]), .A(DP_mult_219_n1637), 
        .ZN(DP_mult_219_n1635) );
  XNOR2_X1 DP_mult_219_U1237 ( .A(DP_coeff_pipe03[2]), .B(DP_mult_219_n1635), 
        .ZN(DP_mult_219_n908) );
  OAI22_X1 DP_mult_219_U1236 ( .A1(DP_mult_219_n1558), .A2(DP_mult_219_n1633), 
        .B1(DP_mult_219_n1557), .B2(DP_mult_219_n1634), .ZN(DP_mult_219_n1632)
         );
  AOI221_X1 DP_mult_219_U1235 ( .B1(DP_mult_219_n1613), .B2(DP_mult_219_n1559), 
        .C1(DP_mult_219_n1560), .C2(DP_mult_219_n1615), .A(DP_mult_219_n1632), 
        .ZN(DP_mult_219_n1631) );
  XOR2_X1 DP_mult_219_U1234 ( .A(DP_coeff_pipe03[23]), .B(DP_mult_219_n1631), 
        .Z(DP_mult_219_n1625) );
  INV_X1 DP_mult_219_U1233 ( .A(DP_mult_219_n1625), .ZN(DP_mult_219_n1621) );
  OAI21_X1 DP_mult_219_U1232 ( .B1(DP_mult_219_n1559), .B2(DP_mult_219_n1560), 
        .A(DP_mult_219_n1615), .ZN(DP_mult_219_n1630) );
  OAI221_X1 DP_mult_219_U1231 ( .B1(DP_mult_219_n1617), .B2(DP_mult_219_n1557), 
        .C1(DP_mult_219_n1617), .C2(DP_mult_219_n1558), .A(DP_mult_219_n1630), 
        .ZN(DP_mult_219_n1628) );
  XOR2_X1 DP_mult_219_U1230 ( .A(DP_mult_219_n1628), .B(DP_mult_219_n1611), 
        .Z(DP_mult_219_n1622) );
  AOI222_X1 DP_mult_219_U1229 ( .A1(DP_mult_219_n1627), .A2(DP_mult_219_n303), 
        .B1(DP_mult_219_n1625), .B2(DP_mult_219_n303), .C1(DP_mult_219_n1627), 
        .C2(DP_mult_219_n1625), .ZN(DP_mult_219_n1624) );
  INV_X1 DP_mult_219_U1228 ( .A(DP_mult_219_n1622), .ZN(DP_mult_219_n1626) );
  OAI22_X1 DP_mult_219_U1227 ( .A1(DP_mult_219_n1624), .A2(DP_mult_219_n1625), 
        .B1(DP_mult_219_n1624), .B2(DP_mult_219_n1626), .ZN(DP_mult_219_n1623)
         );
  AOI21_X1 DP_mult_219_U1226 ( .B1(DP_mult_219_n1621), .B2(DP_mult_219_n1622), 
        .A(DP_mult_219_n1623), .ZN(DP_pipe0_coeff_pipe03[23]) );
  INV_X1 DP_mult_219_U1225 ( .A(DP_mult_219_n1614), .ZN(DP_mult_219_n1620) );
  INV_X1 DP_mult_219_U1224 ( .A(DP_mult_219_n1613), .ZN(DP_mult_219_n1619) );
  INV_X1 DP_mult_219_U1223 ( .A(DP_mult_219_n1613), .ZN(DP_mult_219_n1618) );
  INV_X1 DP_mult_219_U1222 ( .A(DP_mult_219_n1612), .ZN(DP_mult_219_n1617) );
  INV_X1 DP_mult_219_U1221 ( .A(DP_mult_219_n1612), .ZN(DP_mult_219_n1616) );
  CLKBUF_X1 DP_mult_219_U1220 ( .A(DP_pipe03[23]), .Z(DP_mult_219_n1614) );
  CLKBUF_X1 DP_mult_219_U1219 ( .A(DP_pipe03[23]), .Z(DP_mult_219_n1613) );
  CLKBUF_X1 DP_mult_219_U1218 ( .A(DP_pipe03[23]), .Z(DP_mult_219_n1612) );
  BUF_X1 DP_mult_219_U1217 ( .A(DP_mult_219_n1647), .Z(DP_mult_219_n1567) );
  BUF_X1 DP_mult_219_U1216 ( .A(DP_mult_219_n1647), .Z(DP_mult_219_n1566) );
  BUF_X1 DP_mult_219_U1215 ( .A(DP_mult_219_n1647), .Z(DP_mult_219_n1565) );
  INV_X1 DP_mult_219_U1214 ( .A(DP_mult_219_n1616), .ZN(DP_mult_219_n1615) );
  AND2_X1 DP_mult_219_U1213 ( .A1(DP_coeff_pipe03[0]), .A2(DP_mult_219_n2157), 
        .ZN(DP_mult_219_n1555) );
  BUF_X1 DP_mult_219_U1212 ( .A(DP_mult_219_n1636), .Z(DP_mult_219_n1562) );
  OR2_X1 DP_mult_219_U1211 ( .A1(DP_mult_219_n2158), .A2(DP_mult_219_n2157), 
        .ZN(DP_mult_219_n1554) );
  BUF_X1 DP_mult_219_U1210 ( .A(DP_mult_219_n1636), .Z(DP_mult_219_n1563) );
  INV_X1 DP_mult_219_U1209 ( .A(DP_mult_219_n1555), .ZN(DP_mult_219_n1564) );
  NAND3_X1 DP_mult_219_U1208 ( .A1(DP_mult_219_n2157), .A2(DP_mult_219_n2158), 
        .A3(DP_mult_219_n2159), .ZN(DP_mult_219_n1639) );
  INV_X1 DP_mult_219_U1207 ( .A(DP_coeff_pipe03[23]), .ZN(DP_mult_219_n1611)
         );
  INV_X1 DP_mult_219_U1206 ( .A(DP_coeff_pipe03[8]), .ZN(DP_mult_219_n1601) );
  INV_X1 DP_mult_219_U1205 ( .A(DP_coeff_pipe03[5]), .ZN(DP_mult_219_n1599) );
  OR2_X1 DP_mult_219_U1204 ( .A1(DP_mult_219_n1738), .A2(DP_mult_219_n1739), 
        .ZN(DP_mult_219_n1553) );
  OR2_X1 DP_mult_219_U1203 ( .A1(DP_mult_219_n1740), .A2(DP_mult_219_n1741), 
        .ZN(DP_mult_219_n1552) );
  INV_X1 DP_mult_219_U1202 ( .A(DP_mult_219_n1554), .ZN(DP_mult_219_n1561) );
  INV_X1 DP_mult_219_U1201 ( .A(DP_mult_219_n1611), .ZN(DP_mult_219_n1610) );
  BUF_X1 DP_mult_219_U1200 ( .A(DP_coeff_pipe03[20]), .Z(DP_mult_219_n1609) );
  AND2_X1 DP_mult_219_U1199 ( .A1(DP_mult_219_n1738), .A2(DP_mult_219_n1740), 
        .ZN(DP_mult_219_n1551) );
  BUF_X1 DP_mult_219_U1198 ( .A(DP_mult_219_n1654), .Z(DP_mult_219_n1572) );
  BUF_X1 DP_mult_219_U1197 ( .A(DP_mult_219_n1654), .Z(DP_mult_219_n1571) );
  INV_X1 DP_mult_219_U1196 ( .A(DP_mult_219_n1552), .ZN(DP_mult_219_n1569) );
  INV_X1 DP_mult_219_U1195 ( .A(DP_mult_219_n1553), .ZN(DP_mult_219_n1570) );
  INV_X1 DP_mult_219_U1194 ( .A(DP_mult_219_n1601), .ZN(DP_mult_219_n1600) );
  INV_X1 DP_mult_219_U1193 ( .A(DP_mult_219_n1599), .ZN(DP_mult_219_n1598) );
  INV_X1 DP_mult_219_U1192 ( .A(DP_coeff_pipe03[17]), .ZN(DP_mult_219_n1607)
         );
  INV_X1 DP_mult_219_U1191 ( .A(DP_coeff_pipe03[11]), .ZN(DP_mult_219_n1603)
         );
  OR2_X1 DP_mult_219_U1190 ( .A1(DP_mult_219_n2070), .A2(DP_mult_219_n2069), 
        .ZN(DP_mult_219_n1550) );
  AND2_X1 DP_mult_219_U1189 ( .A1(DP_mult_219_n2070), .A2(DP_mult_219_n2068), 
        .ZN(DP_mult_219_n1549) );
  OR2_X1 DP_mult_219_U1188 ( .A1(DP_mult_219_n2068), .A2(DP_mult_219_n2067), 
        .ZN(DP_mult_219_n1548) );
  BUF_X1 DP_mult_219_U1187 ( .A(DP_coeff_pipe03[20]), .Z(DP_mult_219_n1608) );
  INV_X1 DP_mult_219_U1186 ( .A(DP_coeff_pipe03[14]), .ZN(DP_mult_219_n1605)
         );
  OR2_X1 DP_mult_219_U1185 ( .A1(DP_mult_219_n1794), .A2(DP_mult_219_n1795), 
        .ZN(DP_mult_219_n1547) );
  AND2_X1 DP_mult_219_U1184 ( .A1(DP_mult_219_n1794), .A2(DP_mult_219_n1796), 
        .ZN(DP_mult_219_n1546) );
  OR2_X1 DP_mult_219_U1183 ( .A1(DP_mult_219_n1851), .A2(DP_mult_219_n1852), 
        .ZN(DP_mult_219_n1545) );
  OR2_X1 DP_mult_219_U1182 ( .A1(DP_mult_219_n1796), .A2(DP_mult_219_n1797), 
        .ZN(DP_mult_219_n1544) );
  BUF_X1 DP_mult_219_U1181 ( .A(DP_mult_219_n1629), .Z(DP_mult_219_n1556) );
  INV_X1 DP_mult_219_U1180 ( .A(DP_mult_219_n1551), .ZN(DP_mult_219_n1568) );
  INV_X1 DP_mult_219_U1179 ( .A(DP_mult_219_n1605), .ZN(DP_mult_219_n1604) );
  INV_X1 DP_mult_219_U1178 ( .A(DP_mult_219_n1603), .ZN(DP_mult_219_n1602) );
  OR2_X1 DP_mult_219_U1177 ( .A1(DP_mult_219_n2014), .A2(DP_mult_219_n2015), 
        .ZN(DP_mult_219_n1543) );
  AND2_X1 DP_mult_219_U1176 ( .A1(DP_mult_219_n2014), .A2(DP_mult_219_n2016), 
        .ZN(DP_mult_219_n1542) );
  OR2_X1 DP_mult_219_U1175 ( .A1(DP_mult_219_n2016), .A2(DP_mult_219_n2017), 
        .ZN(DP_mult_219_n1541) );
  BUF_X1 DP_mult_219_U1174 ( .A(DP_mult_219_n1629), .Z(DP_mult_219_n1557) );
  INV_X1 DP_mult_219_U1173 ( .A(DP_mult_219_n1548), .ZN(DP_mult_219_n1559) );
  INV_X1 DP_mult_219_U1172 ( .A(DP_mult_219_n1549), .ZN(DP_mult_219_n1558) );
  INV_X1 DP_mult_219_U1171 ( .A(DP_mult_219_n1550), .ZN(DP_mult_219_n1560) );
  INV_X1 DP_mult_219_U1170 ( .A(DP_mult_219_n1607), .ZN(DP_mult_219_n1606) );
  INV_X1 DP_mult_219_U1169 ( .A(DP_mult_219_n1545), .ZN(DP_mult_219_n1579) );
  INV_X1 DP_mult_219_U1168 ( .A(DP_mult_219_n1544), .ZN(DP_mult_219_n1574) );
  OR2_X1 DP_mult_219_U1167 ( .A1(DP_mult_219_n1959), .A2(DP_mult_219_n1960), 
        .ZN(DP_mult_219_n1540) );
  OR2_X1 DP_mult_219_U1166 ( .A1(DP_mult_219_n1904), .A2(DP_mult_219_n1905), 
        .ZN(DP_mult_219_n1539) );
  OR2_X1 DP_mult_219_U1165 ( .A1(DP_mult_219_n1849), .A2(DP_mult_219_n1850), 
        .ZN(DP_mult_219_n1538) );
  BUF_X1 DP_mult_219_U1164 ( .A(DP_mult_219_n1802), .Z(DP_mult_219_n1582) );
  BUF_X1 DP_mult_219_U1163 ( .A(DP_mult_219_n1747), .Z(DP_mult_219_n1577) );
  BUF_X1 DP_mult_219_U1162 ( .A(DP_mult_219_n1802), .Z(DP_mult_219_n1581) );
  BUF_X1 DP_mult_219_U1161 ( .A(DP_mult_219_n1747), .Z(DP_mult_219_n1576) );
  INV_X1 DP_mult_219_U1160 ( .A(DP_mult_219_n1546), .ZN(DP_mult_219_n1573) );
  INV_X1 DP_mult_219_U1159 ( .A(DP_mult_219_n1541), .ZN(DP_mult_219_n1594) );
  INV_X1 DP_mult_219_U1158 ( .A(DP_mult_219_n1547), .ZN(DP_mult_219_n1575) );
  AND2_X1 DP_mult_219_U1157 ( .A1(DP_mult_219_n1959), .A2(DP_mult_219_n1961), 
        .ZN(DP_mult_219_n1537) );
  AND2_X1 DP_mult_219_U1156 ( .A1(DP_mult_219_n1904), .A2(DP_mult_219_n1906), 
        .ZN(DP_mult_219_n1536) );
  AND2_X1 DP_mult_219_U1155 ( .A1(DP_mult_219_n1849), .A2(DP_mult_219_n1851), 
        .ZN(DP_mult_219_n1535) );
  OR2_X1 DP_mult_219_U1154 ( .A1(DP_mult_219_n1961), .A2(DP_mult_219_n1962), 
        .ZN(DP_mult_219_n1534) );
  OR2_X1 DP_mult_219_U1153 ( .A1(DP_mult_219_n1906), .A2(DP_mult_219_n1907), 
        .ZN(DP_mult_219_n1533) );
  BUF_X1 DP_mult_219_U1152 ( .A(DP_mult_219_n1967), .Z(DP_mult_219_n1597) );
  BUF_X1 DP_mult_219_U1151 ( .A(DP_mult_219_n1967), .Z(DP_mult_219_n1596) );
  INV_X1 DP_mult_219_U1150 ( .A(DP_mult_219_n1542), .ZN(DP_mult_219_n1593) );
  INV_X1 DP_mult_219_U1149 ( .A(DP_mult_219_n1543), .ZN(DP_mult_219_n1595) );
  BUF_X1 DP_mult_219_U1148 ( .A(DP_mult_219_n1857), .Z(DP_mult_219_n1587) );
  INV_X1 DP_mult_219_U1147 ( .A(DP_mult_219_n1534), .ZN(DP_mult_219_n1589) );
  INV_X1 DP_mult_219_U1146 ( .A(DP_mult_219_n1533), .ZN(DP_mult_219_n1584) );
  INV_X1 DP_mult_219_U1145 ( .A(DP_mult_219_n1540), .ZN(DP_mult_219_n1590) );
  INV_X1 DP_mult_219_U1144 ( .A(DP_mult_219_n1539), .ZN(DP_mult_219_n1585) );
  INV_X1 DP_mult_219_U1143 ( .A(DP_mult_219_n1538), .ZN(DP_mult_219_n1580) );
  BUF_X1 DP_mult_219_U1142 ( .A(DP_mult_219_n1912), .Z(DP_mult_219_n1592) );
  BUF_X1 DP_mult_219_U1141 ( .A(DP_mult_219_n1912), .Z(DP_mult_219_n1591) );
  BUF_X1 DP_mult_219_U1140 ( .A(DP_mult_219_n1857), .Z(DP_mult_219_n1586) );
  INV_X1 DP_mult_219_U1139 ( .A(DP_mult_219_n1536), .ZN(DP_mult_219_n1583) );
  INV_X1 DP_mult_219_U1138 ( .A(DP_mult_219_n1537), .ZN(DP_mult_219_n1588) );
  INV_X1 DP_mult_219_U1137 ( .A(DP_mult_219_n1535), .ZN(DP_mult_219_n1578) );
  HA_X1 DP_mult_219_U1134 ( .A(DP_pipe03[0]), .B(DP_pipe03[1]), .CO(
        DP_mult_219_n727), .S(DP_mult_219_n1397) );
  FA_X1 DP_mult_219_U1133 ( .A(DP_pipe03[1]), .B(DP_pipe03[2]), .CI(
        DP_mult_219_n727), .CO(DP_mult_219_n726), .S(DP_mult_219_n1396) );
  FA_X1 DP_mult_219_U1132 ( .A(DP_pipe03[2]), .B(DP_pipe03[3]), .CI(
        DP_mult_219_n726), .CO(DP_mult_219_n725), .S(DP_mult_219_n1395) );
  FA_X1 DP_mult_219_U1131 ( .A(DP_pipe03[3]), .B(DP_pipe03[4]), .CI(
        DP_mult_219_n725), .CO(DP_mult_219_n724), .S(DP_mult_219_n1394) );
  FA_X1 DP_mult_219_U1130 ( .A(DP_pipe03[4]), .B(DP_pipe03[5]), .CI(
        DP_mult_219_n724), .CO(DP_mult_219_n723), .S(DP_mult_219_n1393) );
  FA_X1 DP_mult_219_U1129 ( .A(DP_pipe03[5]), .B(DP_pipe03[6]), .CI(
        DP_mult_219_n723), .CO(DP_mult_219_n722), .S(DP_mult_219_n1392) );
  FA_X1 DP_mult_219_U1128 ( .A(DP_pipe03[6]), .B(DP_pipe03[7]), .CI(
        DP_mult_219_n722), .CO(DP_mult_219_n721), .S(DP_mult_219_n1391) );
  FA_X1 DP_mult_219_U1127 ( .A(DP_pipe03[7]), .B(DP_pipe03[8]), .CI(
        DP_mult_219_n721), .CO(DP_mult_219_n720), .S(DP_mult_219_n1390) );
  FA_X1 DP_mult_219_U1126 ( .A(DP_pipe03[8]), .B(DP_pipe03[9]), .CI(
        DP_mult_219_n720), .CO(DP_mult_219_n719), .S(DP_mult_219_n1389) );
  FA_X1 DP_mult_219_U1125 ( .A(DP_pipe03[9]), .B(DP_pipe03[10]), .CI(
        DP_mult_219_n719), .CO(DP_mult_219_n718), .S(DP_mult_219_n1388) );
  FA_X1 DP_mult_219_U1124 ( .A(DP_pipe03[10]), .B(DP_pipe03[11]), .CI(
        DP_mult_219_n718), .CO(DP_mult_219_n717), .S(DP_mult_219_n1387) );
  FA_X1 DP_mult_219_U1123 ( .A(DP_pipe03[11]), .B(DP_pipe03[12]), .CI(
        DP_mult_219_n717), .CO(DP_mult_219_n716), .S(DP_mult_219_n1386) );
  FA_X1 DP_mult_219_U1122 ( .A(DP_pipe03[12]), .B(DP_pipe03[13]), .CI(
        DP_mult_219_n716), .CO(DP_mult_219_n715), .S(DP_mult_219_n1385) );
  FA_X1 DP_mult_219_U1121 ( .A(DP_pipe03[13]), .B(DP_pipe03[14]), .CI(
        DP_mult_219_n715), .CO(DP_mult_219_n714), .S(DP_mult_219_n1384) );
  FA_X1 DP_mult_219_U1120 ( .A(DP_pipe03[14]), .B(DP_pipe03[15]), .CI(
        DP_mult_219_n714), .CO(DP_mult_219_n713), .S(DP_mult_219_n1383) );
  FA_X1 DP_mult_219_U1119 ( .A(DP_pipe03[15]), .B(DP_pipe03[16]), .CI(
        DP_mult_219_n713), .CO(DP_mult_219_n712), .S(DP_mult_219_n1382) );
  FA_X1 DP_mult_219_U1118 ( .A(DP_pipe03[16]), .B(DP_pipe03[17]), .CI(
        DP_mult_219_n712), .CO(DP_mult_219_n711), .S(DP_mult_219_n1381) );
  FA_X1 DP_mult_219_U1117 ( .A(DP_pipe03[17]), .B(DP_pipe03[18]), .CI(
        DP_mult_219_n711), .CO(DP_mult_219_n710), .S(DP_mult_219_n1380) );
  FA_X1 DP_mult_219_U1116 ( .A(DP_pipe03[18]), .B(DP_pipe03[19]), .CI(
        DP_mult_219_n710), .CO(DP_mult_219_n709), .S(DP_mult_219_n1379) );
  FA_X1 DP_mult_219_U1115 ( .A(DP_pipe03[19]), .B(DP_pipe03[20]), .CI(
        DP_mult_219_n709), .CO(DP_mult_219_n708), .S(DP_mult_219_n1378) );
  FA_X1 DP_mult_219_U1114 ( .A(DP_pipe03[20]), .B(DP_pipe03[21]), .CI(
        DP_mult_219_n708), .CO(DP_mult_219_n707), .S(DP_mult_219_n1377) );
  FA_X1 DP_mult_219_U1113 ( .A(DP_pipe03[21]), .B(DP_pipe03[22]), .CI(
        DP_mult_219_n707), .CO(DP_mult_219_n706), .S(DP_mult_219_n1376) );
  FA_X1 DP_mult_219_U1112 ( .A(DP_pipe03[22]), .B(DP_mult_219_n1615), .CI(
        DP_mult_219_n706), .CO(DP_mult_219_n1374), .S(DP_mult_219_n1375) );
  HA_X1 DP_mult_219_U408 ( .A(DP_mult_219_n904), .B(DP_mult_219_n1598), .CO(
        DP_mult_219_n687), .S(DP_mult_219_n688) );
  HA_X1 DP_mult_219_U407 ( .A(DP_mult_219_n687), .B(DP_mult_219_n903), .CO(
        DP_mult_219_n685), .S(DP_mult_219_n686) );
  HA_X1 DP_mult_219_U406 ( .A(DP_mult_219_n685), .B(DP_mult_219_n902), .CO(
        DP_mult_219_n683), .S(DP_mult_219_n684) );
  HA_X1 DP_mult_219_U405 ( .A(DP_mult_219_n878), .B(DP_mult_219_n1600), .CO(
        DP_mult_219_n681), .S(DP_mult_219_n682) );
  FA_X1 DP_mult_219_U404 ( .A(DP_mult_219_n901), .B(DP_mult_219_n682), .CI(
        DP_mult_219_n683), .CO(DP_mult_219_n679), .S(DP_mult_219_n680) );
  HA_X1 DP_mult_219_U403 ( .A(DP_mult_219_n681), .B(DP_mult_219_n877), .CO(
        DP_mult_219_n677), .S(DP_mult_219_n678) );
  FA_X1 DP_mult_219_U402 ( .A(DP_mult_219_n900), .B(DP_mult_219_n678), .CI(
        DP_mult_219_n679), .CO(DP_mult_219_n675), .S(DP_mult_219_n676) );
  HA_X1 DP_mult_219_U401 ( .A(DP_mult_219_n677), .B(DP_mult_219_n876), .CO(
        DP_mult_219_n673), .S(DP_mult_219_n674) );
  FA_X1 DP_mult_219_U400 ( .A(DP_mult_219_n899), .B(DP_mult_219_n674), .CI(
        DP_mult_219_n675), .CO(DP_mult_219_n671), .S(DP_mult_219_n672) );
  HA_X1 DP_mult_219_U399 ( .A(DP_mult_219_n852), .B(DP_mult_219_n1602), .CO(
        DP_mult_219_n669), .S(DP_mult_219_n670) );
  FA_X1 DP_mult_219_U398 ( .A(DP_mult_219_n875), .B(DP_mult_219_n670), .CI(
        DP_mult_219_n673), .CO(DP_mult_219_n667), .S(DP_mult_219_n668) );
  FA_X1 DP_mult_219_U397 ( .A(DP_mult_219_n898), .B(DP_mult_219_n668), .CI(
        DP_mult_219_n671), .CO(DP_mult_219_n665), .S(DP_mult_219_n666) );
  HA_X1 DP_mult_219_U396 ( .A(DP_mult_219_n669), .B(DP_mult_219_n851), .CO(
        DP_mult_219_n663), .S(DP_mult_219_n664) );
  FA_X1 DP_mult_219_U395 ( .A(DP_mult_219_n874), .B(DP_mult_219_n664), .CI(
        DP_mult_219_n667), .CO(DP_mult_219_n661), .S(DP_mult_219_n662) );
  FA_X1 DP_mult_219_U394 ( .A(DP_mult_219_n897), .B(DP_mult_219_n662), .CI(
        DP_mult_219_n665), .CO(DP_mult_219_n659), .S(DP_mult_219_n660) );
  HA_X1 DP_mult_219_U393 ( .A(DP_mult_219_n663), .B(DP_mult_219_n850), .CO(
        DP_mult_219_n657), .S(DP_mult_219_n658) );
  FA_X1 DP_mult_219_U392 ( .A(DP_mult_219_n873), .B(DP_mult_219_n658), .CI(
        DP_mult_219_n661), .CO(DP_mult_219_n655), .S(DP_mult_219_n656) );
  FA_X1 DP_mult_219_U391 ( .A(DP_mult_219_n896), .B(DP_mult_219_n656), .CI(
        DP_mult_219_n659), .CO(DP_mult_219_n653), .S(DP_mult_219_n654) );
  HA_X1 DP_mult_219_U390 ( .A(DP_mult_219_n826), .B(DP_mult_219_n1604), .CO(
        DP_mult_219_n651), .S(DP_mult_219_n652) );
  FA_X1 DP_mult_219_U389 ( .A(DP_mult_219_n849), .B(DP_mult_219_n652), .CI(
        DP_mult_219_n657), .CO(DP_mult_219_n649), .S(DP_mult_219_n650) );
  FA_X1 DP_mult_219_U388 ( .A(DP_mult_219_n872), .B(DP_mult_219_n650), .CI(
        DP_mult_219_n655), .CO(DP_mult_219_n647), .S(DP_mult_219_n648) );
  FA_X1 DP_mult_219_U387 ( .A(DP_mult_219_n895), .B(DP_mult_219_n648), .CI(
        DP_mult_219_n653), .CO(DP_mult_219_n645), .S(DP_mult_219_n646) );
  HA_X1 DP_mult_219_U386 ( .A(DP_mult_219_n651), .B(DP_mult_219_n825), .CO(
        DP_mult_219_n643), .S(DP_mult_219_n644) );
  FA_X1 DP_mult_219_U385 ( .A(DP_mult_219_n848), .B(DP_mult_219_n644), .CI(
        DP_mult_219_n649), .CO(DP_mult_219_n641), .S(DP_mult_219_n642) );
  FA_X1 DP_mult_219_U384 ( .A(DP_mult_219_n871), .B(DP_mult_219_n642), .CI(
        DP_mult_219_n647), .CO(DP_mult_219_n639), .S(DP_mult_219_n640) );
  FA_X1 DP_mult_219_U383 ( .A(DP_mult_219_n894), .B(DP_mult_219_n640), .CI(
        DP_mult_219_n645), .CO(DP_mult_219_n637), .S(DP_mult_219_n638) );
  HA_X1 DP_mult_219_U382 ( .A(DP_mult_219_n643), .B(DP_mult_219_n824), .CO(
        DP_mult_219_n635), .S(DP_mult_219_n636) );
  FA_X1 DP_mult_219_U381 ( .A(DP_mult_219_n847), .B(DP_mult_219_n636), .CI(
        DP_mult_219_n641), .CO(DP_mult_219_n633), .S(DP_mult_219_n634) );
  FA_X1 DP_mult_219_U380 ( .A(DP_mult_219_n870), .B(DP_mult_219_n634), .CI(
        DP_mult_219_n639), .CO(DP_mult_219_n631), .S(DP_mult_219_n632) );
  FA_X1 DP_mult_219_U379 ( .A(DP_mult_219_n893), .B(DP_mult_219_n632), .CI(
        DP_mult_219_n637), .CO(DP_mult_219_n629), .S(DP_mult_219_n630) );
  HA_X1 DP_mult_219_U378 ( .A(DP_mult_219_n800), .B(DP_mult_219_n1606), .CO(
        DP_mult_219_n627), .S(DP_mult_219_n628) );
  FA_X1 DP_mult_219_U377 ( .A(DP_mult_219_n823), .B(DP_mult_219_n628), .CI(
        DP_mult_219_n635), .CO(DP_mult_219_n625), .S(DP_mult_219_n626) );
  FA_X1 DP_mult_219_U376 ( .A(DP_mult_219_n846), .B(DP_mult_219_n626), .CI(
        DP_mult_219_n633), .CO(DP_mult_219_n623), .S(DP_mult_219_n624) );
  FA_X1 DP_mult_219_U375 ( .A(DP_mult_219_n869), .B(DP_mult_219_n624), .CI(
        DP_mult_219_n631), .CO(DP_mult_219_n621), .S(DP_mult_219_n622) );
  FA_X1 DP_mult_219_U374 ( .A(DP_mult_219_n892), .B(DP_mult_219_n622), .CI(
        DP_mult_219_n629), .CO(DP_mult_219_n619), .S(DP_mult_219_n620) );
  HA_X1 DP_mult_219_U373 ( .A(DP_mult_219_n627), .B(DP_mult_219_n799), .CO(
        DP_mult_219_n617), .S(DP_mult_219_n618) );
  FA_X1 DP_mult_219_U372 ( .A(DP_mult_219_n822), .B(DP_mult_219_n618), .CI(
        DP_mult_219_n625), .CO(DP_mult_219_n615), .S(DP_mult_219_n616) );
  FA_X1 DP_mult_219_U371 ( .A(DP_mult_219_n845), .B(DP_mult_219_n616), .CI(
        DP_mult_219_n623), .CO(DP_mult_219_n613), .S(DP_mult_219_n614) );
  FA_X1 DP_mult_219_U370 ( .A(DP_mult_219_n868), .B(DP_mult_219_n614), .CI(
        DP_mult_219_n621), .CO(DP_mult_219_n611), .S(DP_mult_219_n612) );
  FA_X1 DP_mult_219_U369 ( .A(DP_mult_219_n891), .B(DP_mult_219_n612), .CI(
        DP_mult_219_n619), .CO(DP_mult_219_n609), .S(DP_mult_219_n610) );
  HA_X1 DP_mult_219_U368 ( .A(DP_mult_219_n617), .B(DP_mult_219_n798), .CO(
        DP_mult_219_n607), .S(DP_mult_219_n608) );
  FA_X1 DP_mult_219_U367 ( .A(DP_mult_219_n821), .B(DP_mult_219_n608), .CI(
        DP_mult_219_n615), .CO(DP_mult_219_n605), .S(DP_mult_219_n606) );
  FA_X1 DP_mult_219_U366 ( .A(DP_mult_219_n844), .B(DP_mult_219_n606), .CI(
        DP_mult_219_n613), .CO(DP_mult_219_n603), .S(DP_mult_219_n604) );
  FA_X1 DP_mult_219_U365 ( .A(DP_mult_219_n867), .B(DP_mult_219_n604), .CI(
        DP_mult_219_n611), .CO(DP_mult_219_n601), .S(DP_mult_219_n602) );
  FA_X1 DP_mult_219_U364 ( .A(DP_mult_219_n890), .B(DP_mult_219_n602), .CI(
        DP_mult_219_n609), .CO(DP_mult_219_n599), .S(DP_mult_219_n600) );
  HA_X1 DP_mult_219_U363 ( .A(DP_mult_219_n774), .B(DP_mult_219_n1608), .CO(
        DP_mult_219_n597), .S(DP_mult_219_n598) );
  FA_X1 DP_mult_219_U362 ( .A(DP_mult_219_n797), .B(DP_mult_219_n598), .CI(
        DP_mult_219_n607), .CO(DP_mult_219_n595), .S(DP_mult_219_n596) );
  FA_X1 DP_mult_219_U361 ( .A(DP_mult_219_n820), .B(DP_mult_219_n596), .CI(
        DP_mult_219_n605), .CO(DP_mult_219_n593), .S(DP_mult_219_n594) );
  FA_X1 DP_mult_219_U360 ( .A(DP_mult_219_n843), .B(DP_mult_219_n594), .CI(
        DP_mult_219_n603), .CO(DP_mult_219_n591), .S(DP_mult_219_n592) );
  FA_X1 DP_mult_219_U359 ( .A(DP_mult_219_n866), .B(DP_mult_219_n592), .CI(
        DP_mult_219_n601), .CO(DP_mult_219_n589), .S(DP_mult_219_n590) );
  FA_X1 DP_mult_219_U358 ( .A(DP_mult_219_n889), .B(DP_mult_219_n590), .CI(
        DP_mult_219_n599), .CO(DP_mult_219_n587), .S(DP_mult_219_n588) );
  HA_X1 DP_mult_219_U357 ( .A(DP_mult_219_n597), .B(DP_mult_219_n773), .CO(
        DP_mult_219_n585), .S(DP_mult_219_n586) );
  FA_X1 DP_mult_219_U356 ( .A(DP_mult_219_n796), .B(DP_mult_219_n586), .CI(
        DP_mult_219_n595), .CO(DP_mult_219_n583), .S(DP_mult_219_n584) );
  FA_X1 DP_mult_219_U355 ( .A(DP_mult_219_n819), .B(DP_mult_219_n584), .CI(
        DP_mult_219_n593), .CO(DP_mult_219_n581), .S(DP_mult_219_n582) );
  FA_X1 DP_mult_219_U354 ( .A(DP_mult_219_n842), .B(DP_mult_219_n582), .CI(
        DP_mult_219_n591), .CO(DP_mult_219_n579), .S(DP_mult_219_n580) );
  FA_X1 DP_mult_219_U353 ( .A(DP_mult_219_n865), .B(DP_mult_219_n580), .CI(
        DP_mult_219_n589), .CO(DP_mult_219_n577), .S(DP_mult_219_n578) );
  FA_X1 DP_mult_219_U352 ( .A(DP_mult_219_n888), .B(DP_mult_219_n578), .CI(
        DP_mult_219_n587), .CO(DP_mult_219_n575), .S(DP_mult_219_n576) );
  HA_X1 DP_mult_219_U351 ( .A(DP_mult_219_n585), .B(DP_mult_219_n772), .CO(
        DP_mult_219_n573), .S(DP_mult_219_n574) );
  FA_X1 DP_mult_219_U350 ( .A(DP_mult_219_n795), .B(DP_mult_219_n574), .CI(
        DP_mult_219_n583), .CO(DP_mult_219_n571), .S(DP_mult_219_n572) );
  FA_X1 DP_mult_219_U349 ( .A(DP_mult_219_n818), .B(DP_mult_219_n572), .CI(
        DP_mult_219_n581), .CO(DP_mult_219_n569), .S(DP_mult_219_n570) );
  FA_X1 DP_mult_219_U348 ( .A(DP_mult_219_n841), .B(DP_mult_219_n570), .CI(
        DP_mult_219_n579), .CO(DP_mult_219_n567), .S(DP_mult_219_n568) );
  FA_X1 DP_mult_219_U347 ( .A(DP_mult_219_n864), .B(DP_mult_219_n568), .CI(
        DP_mult_219_n577), .CO(DP_mult_219_n565), .S(DP_mult_219_n566) );
  FA_X1 DP_mult_219_U346 ( .A(DP_mult_219_n887), .B(DP_mult_219_n566), .CI(
        DP_mult_219_n575), .CO(DP_mult_219_n563), .S(DP_mult_219_n564) );
  HA_X1 DP_mult_219_U345 ( .A(DP_mult_219_n748), .B(DP_mult_219_n1610), .CO(
        DP_mult_219_n561), .S(DP_mult_219_n562) );
  FA_X1 DP_mult_219_U344 ( .A(DP_mult_219_n771), .B(DP_mult_219_n562), .CI(
        DP_mult_219_n573), .CO(DP_mult_219_n559), .S(DP_mult_219_n560) );
  FA_X1 DP_mult_219_U343 ( .A(DP_mult_219_n794), .B(DP_mult_219_n560), .CI(
        DP_mult_219_n571), .CO(DP_mult_219_n557), .S(DP_mult_219_n558) );
  FA_X1 DP_mult_219_U342 ( .A(DP_mult_219_n817), .B(DP_mult_219_n558), .CI(
        DP_mult_219_n569), .CO(DP_mult_219_n555), .S(DP_mult_219_n556) );
  FA_X1 DP_mult_219_U341 ( .A(DP_mult_219_n840), .B(DP_mult_219_n556), .CI(
        DP_mult_219_n567), .CO(DP_mult_219_n553), .S(DP_mult_219_n554) );
  FA_X1 DP_mult_219_U340 ( .A(DP_mult_219_n863), .B(DP_mult_219_n554), .CI(
        DP_mult_219_n565), .CO(DP_mult_219_n551), .S(DP_mult_219_n552) );
  FA_X1 DP_mult_219_U339 ( .A(DP_mult_219_n886), .B(DP_mult_219_n552), .CI(
        DP_mult_219_n563), .CO(DP_mult_219_n549), .S(DP_mult_219_n550) );
  HA_X1 DP_mult_219_U338 ( .A(DP_mult_219_n561), .B(DP_mult_219_n747), .CO(
        DP_mult_219_n547), .S(DP_mult_219_n548) );
  FA_X1 DP_mult_219_U337 ( .A(DP_mult_219_n770), .B(DP_mult_219_n548), .CI(
        DP_mult_219_n559), .CO(DP_mult_219_n545), .S(DP_mult_219_n546) );
  FA_X1 DP_mult_219_U336 ( .A(DP_mult_219_n793), .B(DP_mult_219_n546), .CI(
        DP_mult_219_n557), .CO(DP_mult_219_n543), .S(DP_mult_219_n544) );
  FA_X1 DP_mult_219_U335 ( .A(DP_mult_219_n816), .B(DP_mult_219_n544), .CI(
        DP_mult_219_n555), .CO(DP_mult_219_n541), .S(DP_mult_219_n542) );
  FA_X1 DP_mult_219_U334 ( .A(DP_mult_219_n839), .B(DP_mult_219_n542), .CI(
        DP_mult_219_n553), .CO(DP_mult_219_n539), .S(DP_mult_219_n540) );
  FA_X1 DP_mult_219_U333 ( .A(DP_mult_219_n862), .B(DP_mult_219_n540), .CI(
        DP_mult_219_n551), .CO(DP_mult_219_n537), .S(DP_mult_219_n538) );
  FA_X1 DP_mult_219_U332 ( .A(DP_mult_219_n885), .B(DP_mult_219_n538), .CI(
        DP_mult_219_n549), .CO(DP_mult_219_n535), .S(DP_mult_219_n536) );
  HA_X1 DP_mult_219_U331 ( .A(DP_mult_219_n547), .B(DP_mult_219_n746), .CO(
        DP_mult_219_n533), .S(DP_mult_219_n534) );
  FA_X1 DP_mult_219_U330 ( .A(DP_mult_219_n769), .B(DP_mult_219_n534), .CI(
        DP_mult_219_n545), .CO(DP_mult_219_n531), .S(DP_mult_219_n532) );
  FA_X1 DP_mult_219_U329 ( .A(DP_mult_219_n792), .B(DP_mult_219_n532), .CI(
        DP_mult_219_n543), .CO(DP_mult_219_n529), .S(DP_mult_219_n530) );
  FA_X1 DP_mult_219_U328 ( .A(DP_mult_219_n815), .B(DP_mult_219_n530), .CI(
        DP_mult_219_n541), .CO(DP_mult_219_n527), .S(DP_mult_219_n528) );
  FA_X1 DP_mult_219_U327 ( .A(DP_mult_219_n838), .B(DP_mult_219_n528), .CI(
        DP_mult_219_n539), .CO(DP_mult_219_n525), .S(DP_mult_219_n526) );
  FA_X1 DP_mult_219_U326 ( .A(DP_mult_219_n861), .B(DP_mult_219_n526), .CI(
        DP_mult_219_n537), .CO(DP_mult_219_n523), .S(DP_mult_219_n524) );
  FA_X1 DP_mult_219_U325 ( .A(DP_mult_219_n884), .B(DP_mult_219_n524), .CI(
        DP_mult_219_n535), .CO(DP_mult_219_n521), .S(DP_mult_219_n522) );
  HA_X1 DP_mult_219_U324 ( .A(DP_mult_219_n533), .B(DP_mult_219_n745), .CO(
        DP_mult_219_n519), .S(DP_mult_219_n520) );
  FA_X1 DP_mult_219_U323 ( .A(DP_mult_219_n768), .B(DP_mult_219_n520), .CI(
        DP_mult_219_n531), .CO(DP_mult_219_n517), .S(DP_mult_219_n518) );
  FA_X1 DP_mult_219_U322 ( .A(DP_mult_219_n791), .B(DP_mult_219_n518), .CI(
        DP_mult_219_n529), .CO(DP_mult_219_n515), .S(DP_mult_219_n516) );
  FA_X1 DP_mult_219_U321 ( .A(DP_mult_219_n814), .B(DP_mult_219_n516), .CI(
        DP_mult_219_n527), .CO(DP_mult_219_n513), .S(DP_mult_219_n514) );
  FA_X1 DP_mult_219_U320 ( .A(DP_mult_219_n837), .B(DP_mult_219_n514), .CI(
        DP_mult_219_n525), .CO(DP_mult_219_n511), .S(DP_mult_219_n512) );
  FA_X1 DP_mult_219_U319 ( .A(DP_mult_219_n860), .B(DP_mult_219_n512), .CI(
        DP_mult_219_n523), .CO(DP_mult_219_n509), .S(DP_mult_219_n510) );
  FA_X1 DP_mult_219_U318 ( .A(DP_mult_219_n883), .B(DP_mult_219_n510), .CI(
        DP_mult_219_n521), .CO(DP_mult_219_n507), .S(DP_mult_219_n508) );
  FA_X1 DP_mult_219_U315 ( .A(DP_mult_219_n506), .B(DP_mult_219_n744), .CI(
        DP_mult_219_n767), .CO(DP_mult_219_n504), .S(DP_mult_219_n505) );
  FA_X1 DP_mult_219_U314 ( .A(DP_mult_219_n505), .B(DP_mult_219_n517), .CI(
        DP_mult_219_n790), .CO(DP_mult_219_n502), .S(DP_mult_219_n503) );
  FA_X1 DP_mult_219_U313 ( .A(DP_mult_219_n503), .B(DP_mult_219_n515), .CI(
        DP_mult_219_n813), .CO(DP_mult_219_n500), .S(DP_mult_219_n501) );
  FA_X1 DP_mult_219_U312 ( .A(DP_mult_219_n501), .B(DP_mult_219_n513), .CI(
        DP_mult_219_n836), .CO(DP_mult_219_n498), .S(DP_mult_219_n499) );
  FA_X1 DP_mult_219_U311 ( .A(DP_mult_219_n499), .B(DP_mult_219_n511), .CI(
        DP_mult_219_n859), .CO(DP_mult_219_n496), .S(DP_mult_219_n497) );
  FA_X1 DP_mult_219_U310 ( .A(DP_mult_219_n497), .B(DP_mult_219_n509), .CI(
        DP_mult_219_n882), .CO(DP_mult_219_n494), .S(DP_mult_219_n495) );
  FA_X1 DP_mult_219_U308 ( .A(DP_mult_219_n743), .B(DP_mult_219_n493), .CI(
        DP_mult_219_n766), .CO(DP_mult_219_n491), .S(DP_mult_219_n492) );
  FA_X1 DP_mult_219_U307 ( .A(DP_mult_219_n492), .B(DP_mult_219_n504), .CI(
        DP_mult_219_n789), .CO(DP_mult_219_n489), .S(DP_mult_219_n490) );
  FA_X1 DP_mult_219_U306 ( .A(DP_mult_219_n490), .B(DP_mult_219_n502), .CI(
        DP_mult_219_n500), .CO(DP_mult_219_n487), .S(DP_mult_219_n488) );
  FA_X1 DP_mult_219_U305 ( .A(DP_mult_219_n488), .B(DP_mult_219_n812), .CI(
        DP_mult_219_n835), .CO(DP_mult_219_n485), .S(DP_mult_219_n486) );
  FA_X1 DP_mult_219_U304 ( .A(DP_mult_219_n486), .B(DP_mult_219_n498), .CI(
        DP_mult_219_n496), .CO(DP_mult_219_n483), .S(DP_mult_219_n484) );
  FA_X1 DP_mult_219_U303 ( .A(DP_mult_219_n484), .B(DP_mult_219_n858), .CI(
        DP_mult_219_n881), .CO(DP_mult_219_n481), .S(DP_mult_219_n482) );
  FA_X1 DP_mult_219_U301 ( .A(DP_mult_219_n742), .B(DP_mult_219_n493), .CI(
        DP_mult_219_n491), .CO(DP_mult_219_n477), .S(DP_mult_219_n478) );
  FA_X1 DP_mult_219_U300 ( .A(DP_mult_219_n478), .B(DP_mult_219_n765), .CI(
        DP_mult_219_n788), .CO(DP_mult_219_n475), .S(DP_mult_219_n476) );
  FA_X1 DP_mult_219_U299 ( .A(DP_mult_219_n476), .B(DP_mult_219_n489), .CI(
        DP_mult_219_n487), .CO(DP_mult_219_n473), .S(DP_mult_219_n474) );
  FA_X1 DP_mult_219_U298 ( .A(DP_mult_219_n474), .B(DP_mult_219_n811), .CI(
        DP_mult_219_n834), .CO(DP_mult_219_n471), .S(DP_mult_219_n472) );
  FA_X1 DP_mult_219_U297 ( .A(DP_mult_219_n472), .B(DP_mult_219_n485), .CI(
        DP_mult_219_n483), .CO(DP_mult_219_n469), .S(DP_mult_219_n470) );
  FA_X1 DP_mult_219_U296 ( .A(DP_mult_219_n880), .B(DP_mult_219_n857), .CI(
        DP_mult_219_n470), .CO(DP_mult_219_n467), .S(DP_mult_219_n468) );
  FA_X1 DP_mult_219_U295 ( .A(DP_mult_219_n479), .B(DP_mult_219_n879), .CI(
        DP_mult_219_n741), .CO(DP_mult_219_n465), .S(DP_mult_219_n466) );
  FA_X1 DP_mult_219_U294 ( .A(DP_mult_219_n764), .B(DP_mult_219_n466), .CI(
        DP_mult_219_n477), .CO(DP_mult_219_n463), .S(DP_mult_219_n464) );
  FA_X1 DP_mult_219_U293 ( .A(DP_mult_219_n475), .B(DP_mult_219_n464), .CI(
        DP_mult_219_n787), .CO(DP_mult_219_n461), .S(DP_mult_219_n462) );
  FA_X1 DP_mult_219_U292 ( .A(DP_mult_219_n810), .B(DP_mult_219_n462), .CI(
        DP_mult_219_n473), .CO(DP_mult_219_n459), .S(DP_mult_219_n460) );
  FA_X1 DP_mult_219_U291 ( .A(DP_mult_219_n471), .B(DP_mult_219_n460), .CI(
        DP_mult_219_n833), .CO(DP_mult_219_n457), .S(DP_mult_219_n458) );
  FA_X1 DP_mult_219_U290 ( .A(DP_mult_219_n856), .B(DP_mult_219_n458), .CI(
        DP_mult_219_n469), .CO(DP_mult_219_n455), .S(DP_mult_219_n456) );
  FA_X1 DP_mult_219_U288 ( .A(DP_mult_219_n454), .B(DP_mult_219_n465), .CI(
        DP_mult_219_n763), .CO(DP_mult_219_n452), .S(DP_mult_219_n453) );
  FA_X1 DP_mult_219_U287 ( .A(DP_mult_219_n453), .B(DP_mult_219_n463), .CI(
        DP_mult_219_n786), .CO(DP_mult_219_n450), .S(DP_mult_219_n451) );
  FA_X1 DP_mult_219_U286 ( .A(DP_mult_219_n451), .B(DP_mult_219_n461), .CI(
        DP_mult_219_n809), .CO(DP_mult_219_n448), .S(DP_mult_219_n449) );
  FA_X1 DP_mult_219_U285 ( .A(DP_mult_219_n449), .B(DP_mult_219_n459), .CI(
        DP_mult_219_n832), .CO(DP_mult_219_n446), .S(DP_mult_219_n447) );
  FA_X1 DP_mult_219_U284 ( .A(DP_mult_219_n447), .B(DP_mult_219_n457), .CI(
        DP_mult_219_n855), .CO(DP_mult_219_n444), .S(DP_mult_219_n445) );
  FA_X1 DP_mult_219_U282 ( .A(DP_mult_219_n740), .B(DP_mult_219_n454), .CI(
        DP_mult_219_n762), .CO(DP_mult_219_n440), .S(DP_mult_219_n441) );
  FA_X1 DP_mult_219_U281 ( .A(DP_mult_219_n441), .B(DP_mult_219_n452), .CI(
        DP_mult_219_n450), .CO(DP_mult_219_n438), .S(DP_mult_219_n439) );
  FA_X1 DP_mult_219_U280 ( .A(DP_mult_219_n439), .B(DP_mult_219_n785), .CI(
        DP_mult_219_n808), .CO(DP_mult_219_n436), .S(DP_mult_219_n437) );
  FA_X1 DP_mult_219_U279 ( .A(DP_mult_219_n437), .B(DP_mult_219_n448), .CI(
        DP_mult_219_n446), .CO(DP_mult_219_n434), .S(DP_mult_219_n435) );
  FA_X1 DP_mult_219_U278 ( .A(DP_mult_219_n854), .B(DP_mult_219_n831), .CI(
        DP_mult_219_n435), .CO(DP_mult_219_n432), .S(DP_mult_219_n433) );
  FA_X1 DP_mult_219_U277 ( .A(DP_mult_219_n442), .B(DP_mult_219_n853), .CI(
        DP_mult_219_n739), .CO(DP_mult_219_n430), .S(DP_mult_219_n431) );
  FA_X1 DP_mult_219_U276 ( .A(DP_mult_219_n440), .B(DP_mult_219_n431), .CI(
        DP_mult_219_n761), .CO(DP_mult_219_n428), .S(DP_mult_219_n429) );
  FA_X1 DP_mult_219_U275 ( .A(DP_mult_219_n784), .B(DP_mult_219_n429), .CI(
        DP_mult_219_n438), .CO(DP_mult_219_n426), .S(DP_mult_219_n427) );
  FA_X1 DP_mult_219_U274 ( .A(DP_mult_219_n436), .B(DP_mult_219_n427), .CI(
        DP_mult_219_n807), .CO(DP_mult_219_n424), .S(DP_mult_219_n425) );
  FA_X1 DP_mult_219_U273 ( .A(DP_mult_219_n830), .B(DP_mult_219_n425), .CI(
        DP_mult_219_n434), .CO(DP_mult_219_n422), .S(DP_mult_219_n423) );
  FA_X1 DP_mult_219_U271 ( .A(DP_mult_219_n421), .B(DP_mult_219_n430), .CI(
        DP_mult_219_n760), .CO(DP_mult_219_n419), .S(DP_mult_219_n420) );
  FA_X1 DP_mult_219_U270 ( .A(DP_mult_219_n420), .B(DP_mult_219_n428), .CI(
        DP_mult_219_n783), .CO(DP_mult_219_n417), .S(DP_mult_219_n418) );
  FA_X1 DP_mult_219_U269 ( .A(DP_mult_219_n418), .B(DP_mult_219_n426), .CI(
        DP_mult_219_n806), .CO(DP_mult_219_n415), .S(DP_mult_219_n416) );
  FA_X1 DP_mult_219_U268 ( .A(DP_mult_219_n416), .B(DP_mult_219_n424), .CI(
        DP_mult_219_n829), .CO(DP_mult_219_n413), .S(DP_mult_219_n414) );
  FA_X1 DP_mult_219_U266 ( .A(DP_mult_219_n738), .B(DP_mult_219_n421), .CI(
        DP_mult_219_n419), .CO(DP_mult_219_n409), .S(DP_mult_219_n410) );
  FA_X1 DP_mult_219_U265 ( .A(DP_mult_219_n410), .B(DP_mult_219_n759), .CI(
        DP_mult_219_n782), .CO(DP_mult_219_n407), .S(DP_mult_219_n408) );
  FA_X1 DP_mult_219_U264 ( .A(DP_mult_219_n408), .B(DP_mult_219_n417), .CI(
        DP_mult_219_n415), .CO(DP_mult_219_n405), .S(DP_mult_219_n406) );
  FA_X1 DP_mult_219_U263 ( .A(DP_mult_219_n828), .B(DP_mult_219_n805), .CI(
        DP_mult_219_n406), .CO(DP_mult_219_n403), .S(DP_mult_219_n404) );
  FA_X1 DP_mult_219_U262 ( .A(DP_mult_219_n411), .B(DP_mult_219_n827), .CI(
        DP_mult_219_n737), .CO(DP_mult_219_n387), .S(DP_mult_219_n402) );
  FA_X1 DP_mult_219_U261 ( .A(DP_mult_219_n758), .B(DP_mult_219_n402), .CI(
        DP_mult_219_n409), .CO(DP_mult_219_n400), .S(DP_mult_219_n401) );
  FA_X1 DP_mult_219_U260 ( .A(DP_mult_219_n407), .B(DP_mult_219_n401), .CI(
        DP_mult_219_n781), .CO(DP_mult_219_n398), .S(DP_mult_219_n399) );
  FA_X1 DP_mult_219_U259 ( .A(DP_mult_219_n804), .B(DP_mult_219_n399), .CI(
        DP_mult_219_n405), .CO(DP_mult_219_n396), .S(DP_mult_219_n397) );
  FA_X1 DP_mult_219_U257 ( .A(DP_mult_219_n395), .B(DP_mult_219_n736), .CI(
        DP_mult_219_n757), .CO(DP_mult_219_n393), .S(DP_mult_219_n394) );
  FA_X1 DP_mult_219_U256 ( .A(DP_mult_219_n394), .B(DP_mult_219_n400), .CI(
        DP_mult_219_n780), .CO(DP_mult_219_n391), .S(DP_mult_219_n392) );
  FA_X1 DP_mult_219_U255 ( .A(DP_mult_219_n392), .B(DP_mult_219_n398), .CI(
        DP_mult_219_n803), .CO(DP_mult_219_n389), .S(DP_mult_219_n390) );
  FA_X1 DP_mult_219_U253 ( .A(DP_mult_219_n735), .B(DP_mult_219_n395), .CI(
        DP_mult_219_n756), .CO(DP_mult_219_n385), .S(DP_mult_219_n386) );
  FA_X1 DP_mult_219_U252 ( .A(DP_mult_219_n386), .B(DP_mult_219_n393), .CI(
        DP_mult_219_n391), .CO(DP_mult_219_n383), .S(DP_mult_219_n384) );
  FA_X1 DP_mult_219_U251 ( .A(DP_mult_219_n802), .B(DP_mult_219_n779), .CI(
        DP_mult_219_n384), .CO(DP_mult_219_n381), .S(DP_mult_219_n382) );
  FA_X1 DP_mult_219_U250 ( .A(DP_mult_219_n387), .B(DP_mult_219_n801), .CI(
        DP_mult_219_n734), .CO(DP_mult_219_n379), .S(DP_mult_219_n380) );
  FA_X1 DP_mult_219_U249 ( .A(DP_mult_219_n385), .B(DP_mult_219_n380), .CI(
        DP_mult_219_n755), .CO(DP_mult_219_n377), .S(DP_mult_219_n378) );
  FA_X1 DP_mult_219_U248 ( .A(DP_mult_219_n778), .B(DP_mult_219_n378), .CI(
        DP_mult_219_n383), .CO(DP_mult_219_n375), .S(DP_mult_219_n376) );
  FA_X1 DP_mult_219_U246 ( .A(DP_mult_219_n374), .B(DP_mult_219_n379), .CI(
        DP_mult_219_n754), .CO(DP_mult_219_n372), .S(DP_mult_219_n373) );
  FA_X1 DP_mult_219_U245 ( .A(DP_mult_219_n373), .B(DP_mult_219_n377), .CI(
        DP_mult_219_n777), .CO(DP_mult_219_n370), .S(DP_mult_219_n371) );
  FA_X1 DP_mult_219_U243 ( .A(DP_mult_219_n733), .B(DP_mult_219_n374), .CI(
        DP_mult_219_n372), .CO(DP_mult_219_n366), .S(DP_mult_219_n367) );
  FA_X1 DP_mult_219_U242 ( .A(DP_mult_219_n776), .B(DP_mult_219_n753), .CI(
        DP_mult_219_n367), .CO(DP_mult_219_n364), .S(DP_mult_219_n365) );
  FA_X1 DP_mult_219_U241 ( .A(DP_mult_219_n368), .B(DP_mult_219_n775), .CI(
        DP_mult_219_n732), .CO(DP_mult_219_n356), .S(DP_mult_219_n363) );
  FA_X1 DP_mult_219_U240 ( .A(DP_mult_219_n752), .B(DP_mult_219_n363), .CI(
        DP_mult_219_n366), .CO(DP_mult_219_n361), .S(DP_mult_219_n362) );
  FA_X1 DP_mult_219_U238 ( .A(DP_mult_219_n360), .B(DP_mult_219_n731), .CI(
        DP_mult_219_n751), .CO(DP_mult_219_n358), .S(DP_mult_219_n359) );
  FA_X1 DP_mult_219_U236 ( .A(DP_mult_219_n730), .B(DP_mult_219_n360), .CI(
        DP_mult_219_n750), .CO(DP_mult_219_n354), .S(DP_mult_219_n355) );
  FA_X1 DP_mult_219_U235 ( .A(DP_mult_219_n356), .B(DP_mult_219_n749), .CI(
        DP_mult_219_n729), .CO(DP_mult_219_n352), .S(DP_mult_219_n353) );
  FA_X1 DP_mult_219_U204 ( .A(DP_mult_219_n908), .B(DP_mult_219_n536), .CI(
        DP_mult_219_n326), .CO(DP_mult_219_n325), .S(DP_pipe0_coeff_pipe03[0])
         );
  FA_X1 DP_mult_219_U203 ( .A(DP_mult_219_n907), .B(DP_mult_219_n522), .CI(
        DP_mult_219_n325), .CO(DP_mult_219_n324), .S(DP_pipe0_coeff_pipe03[1])
         );
  FA_X1 DP_mult_219_U202 ( .A(DP_mult_219_n508), .B(DP_mult_219_n906), .CI(
        DP_mult_219_n324), .CO(DP_mult_219_n323), .S(DP_pipe0_coeff_pipe03[2])
         );
  FA_X1 DP_mult_219_U201 ( .A(DP_mult_219_n495), .B(DP_mult_219_n507), .CI(
        DP_mult_219_n323), .CO(DP_mult_219_n322), .S(DP_pipe0_coeff_pipe03[3])
         );
  FA_X1 DP_mult_219_U200 ( .A(DP_mult_219_n482), .B(DP_mult_219_n494), .CI(
        DP_mult_219_n322), .CO(DP_mult_219_n321), .S(DP_pipe0_coeff_pipe03[4])
         );
  FA_X1 DP_mult_219_U199 ( .A(DP_mult_219_n468), .B(DP_mult_219_n481), .CI(
        DP_mult_219_n321), .CO(DP_mult_219_n320), .S(DP_pipe0_coeff_pipe03[5])
         );
  FA_X1 DP_mult_219_U198 ( .A(DP_mult_219_n456), .B(DP_mult_219_n467), .CI(
        DP_mult_219_n320), .CO(DP_mult_219_n319), .S(DP_pipe0_coeff_pipe03[6])
         );
  FA_X1 DP_mult_219_U197 ( .A(DP_mult_219_n445), .B(DP_mult_219_n455), .CI(
        DP_mult_219_n319), .CO(DP_mult_219_n318), .S(DP_pipe0_coeff_pipe03[7])
         );
  FA_X1 DP_mult_219_U196 ( .A(DP_mult_219_n433), .B(DP_mult_219_n444), .CI(
        DP_mult_219_n318), .CO(DP_mult_219_n317), .S(DP_pipe0_coeff_pipe03[8])
         );
  FA_X1 DP_mult_219_U195 ( .A(DP_mult_219_n423), .B(DP_mult_219_n432), .CI(
        DP_mult_219_n317), .CO(DP_mult_219_n316), .S(DP_pipe0_coeff_pipe03[9])
         );
  FA_X1 DP_mult_219_U194 ( .A(DP_mult_219_n414), .B(DP_mult_219_n422), .CI(
        DP_mult_219_n316), .CO(DP_mult_219_n315), .S(DP_pipe0_coeff_pipe03[10]) );
  FA_X1 DP_mult_219_U193 ( .A(DP_mult_219_n404), .B(DP_mult_219_n413), .CI(
        DP_mult_219_n315), .CO(DP_mult_219_n314), .S(DP_pipe0_coeff_pipe03[11]) );
  FA_X1 DP_mult_219_U192 ( .A(DP_mult_219_n397), .B(DP_mult_219_n403), .CI(
        DP_mult_219_n314), .CO(DP_mult_219_n313), .S(DP_pipe0_coeff_pipe03[12]) );
  FA_X1 DP_mult_219_U191 ( .A(DP_mult_219_n390), .B(DP_mult_219_n396), .CI(
        DP_mult_219_n313), .CO(DP_mult_219_n312), .S(DP_pipe0_coeff_pipe03[13]) );
  FA_X1 DP_mult_219_U190 ( .A(DP_mult_219_n382), .B(DP_mult_219_n389), .CI(
        DP_mult_219_n312), .CO(DP_mult_219_n311), .S(DP_pipe0_coeff_pipe03[14]) );
  FA_X1 DP_mult_219_U189 ( .A(DP_mult_219_n376), .B(DP_mult_219_n381), .CI(
        DP_mult_219_n311), .CO(DP_mult_219_n310), .S(DP_pipe0_coeff_pipe03[15]) );
  FA_X1 DP_mult_219_U188 ( .A(DP_mult_219_n371), .B(DP_mult_219_n375), .CI(
        DP_mult_219_n310), .CO(DP_mult_219_n309), .S(DP_pipe0_coeff_pipe03[16]) );
  FA_X1 DP_mult_219_U187 ( .A(DP_mult_219_n365), .B(DP_mult_219_n370), .CI(
        DP_mult_219_n309), .CO(DP_mult_219_n308), .S(DP_pipe0_coeff_pipe03[17]) );
  FA_X1 DP_mult_219_U186 ( .A(DP_mult_219_n362), .B(DP_mult_219_n364), .CI(
        DP_mult_219_n308), .CO(DP_mult_219_n307), .S(DP_pipe0_coeff_pipe03[18]) );
  FA_X1 DP_mult_219_U185 ( .A(DP_mult_219_n359), .B(DP_mult_219_n361), .CI(
        DP_mult_219_n307), .CO(DP_mult_219_n306), .S(DP_pipe0_coeff_pipe03[19]) );
  FA_X1 DP_mult_219_U184 ( .A(DP_mult_219_n355), .B(DP_mult_219_n358), .CI(
        DP_mult_219_n306), .CO(DP_mult_219_n305), .S(DP_pipe0_coeff_pipe03[20]) );
  FA_X1 DP_mult_219_U183 ( .A(DP_mult_219_n353), .B(DP_mult_219_n354), .CI(
        DP_mult_219_n305), .CO(DP_mult_219_n304), .S(DP_pipe0_coeff_pipe03[21]) );
  FA_X1 DP_mult_219_U182 ( .A(DP_mult_219_n351), .B(DP_mult_219_n352), .CI(
        DP_mult_219_n304), .CO(DP_mult_219_n303), .S(DP_pipe0_coeff_pipe03[22]) );
  INV_X1 DP_mult_218_U1959 ( .A(DP_coeff_pipe02[1]), .ZN(DP_mult_218_n2159) );
  NOR2_X1 DP_mult_218_U1958 ( .A1(DP_mult_218_n2159), .A2(DP_coeff_pipe02[0]), 
        .ZN(DP_mult_218_n1636) );
  INV_X1 DP_mult_218_U1957 ( .A(DP_coeff_pipe02[2]), .ZN(DP_mult_218_n1742) );
  XNOR2_X1 DP_mult_218_U1956 ( .A(DP_coeff_pipe02[1]), .B(DP_mult_218_n1742), 
        .ZN(DP_mult_218_n2157) );
  AOI221_X1 DP_mult_218_U1955 ( .B1(DP_pipe02[1]), .B2(DP_mult_218_n1563), 
        .C1(DP_mult_218_n1396), .C2(DP_mult_218_n1554), .A(DP_mult_218_n1742), 
        .ZN(DP_mult_218_n2160) );
  INV_X1 DP_mult_218_U1954 ( .A(DP_coeff_pipe02[0]), .ZN(DP_mult_218_n2158) );
  INV_X1 DP_mult_218_U1953 ( .A(DP_pipe02[2]), .ZN(DP_mult_218_n1661) );
  INV_X1 DP_mult_218_U1952 ( .A(DP_mult_218_n1397), .ZN(DP_mult_218_n1650) );
  OAI22_X1 DP_mult_218_U1951 ( .A1(DP_mult_218_n1542), .A2(DP_mult_218_n1661), 
        .B1(DP_mult_218_n1564), .B2(DP_mult_218_n1650), .ZN(DP_mult_218_n2162)
         );
  AOI211_X1 DP_mult_218_U1950 ( .C1(DP_pipe02[1]), .C2(DP_mult_218_n1561), .A(
        DP_mult_218_n2162), .B(DP_pipe02[0]), .ZN(DP_mult_218_n2161) );
  AND2_X1 DP_mult_218_U1949 ( .A1(DP_mult_218_n2160), .A2(DP_mult_218_n2161), 
        .ZN(DP_mult_218_n2153) );
  INV_X1 DP_mult_218_U1948 ( .A(DP_mult_218_n1395), .ZN(DP_mult_218_n1657) );
  INV_X1 DP_mult_218_U1947 ( .A(DP_pipe02[1]), .ZN(DP_mult_218_n1649) );
  OAI22_X1 DP_mult_218_U1946 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1657), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1649), .ZN(DP_mult_218_n2156)
         );
  AOI221_X1 DP_mult_218_U1945 ( .B1(DP_pipe02[3]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[2]), .C2(DP_mult_218_n1563), .A(DP_mult_218_n2156), .ZN(
        DP_mult_218_n2155) );
  XNOR2_X1 DP_mult_218_U1944 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2155), 
        .ZN(DP_mult_218_n2154) );
  AOI222_X1 DP_mult_218_U1943 ( .A1(DP_mult_218_n2153), .A2(DP_mult_218_n2154), 
        .B1(DP_mult_218_n2153), .B2(DP_mult_218_n688), .C1(DP_mult_218_n688), 
        .C2(DP_mult_218_n2154), .ZN(DP_mult_218_n2148) );
  INV_X1 DP_mult_218_U1942 ( .A(DP_mult_218_n1394), .ZN(DP_mult_218_n1660) );
  OAI22_X1 DP_mult_218_U1941 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1660), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1661), .ZN(DP_mult_218_n2152)
         );
  AOI221_X1 DP_mult_218_U1940 ( .B1(DP_pipe02[4]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[3]), .C2(DP_mult_218_n1563), .A(DP_mult_218_n2152), .ZN(
        DP_mult_218_n2151) );
  XNOR2_X1 DP_mult_218_U1939 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2151), 
        .ZN(DP_mult_218_n2149) );
  INV_X1 DP_mult_218_U1938 ( .A(DP_mult_218_n686), .ZN(DP_mult_218_n2150) );
  OAI222_X1 DP_mult_218_U1937 ( .A1(DP_mult_218_n2148), .A2(DP_mult_218_n2149), 
        .B1(DP_mult_218_n2148), .B2(DP_mult_218_n2150), .C1(DP_mult_218_n2150), 
        .C2(DP_mult_218_n2149), .ZN(DP_mult_218_n2144) );
  INV_X1 DP_mult_218_U1936 ( .A(DP_mult_218_n1393), .ZN(DP_mult_218_n1664) );
  INV_X1 DP_mult_218_U1935 ( .A(DP_pipe02[3]), .ZN(DP_mult_218_n1665) );
  OAI22_X1 DP_mult_218_U1934 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1664), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1665), .ZN(DP_mult_218_n2147)
         );
  AOI221_X1 DP_mult_218_U1933 ( .B1(DP_pipe02[5]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[4]), .C2(DP_mult_218_n1563), .A(DP_mult_218_n2147), .ZN(
        DP_mult_218_n2146) );
  XNOR2_X1 DP_mult_218_U1932 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2146), 
        .ZN(DP_mult_218_n2145) );
  AOI222_X1 DP_mult_218_U1931 ( .A1(DP_mult_218_n2144), .A2(DP_mult_218_n2145), 
        .B1(DP_mult_218_n2144), .B2(DP_mult_218_n684), .C1(DP_mult_218_n684), 
        .C2(DP_mult_218_n2145), .ZN(DP_mult_218_n2139) );
  INV_X1 DP_mult_218_U1930 ( .A(DP_mult_218_n1392), .ZN(DP_mult_218_n1668) );
  INV_X1 DP_mult_218_U1929 ( .A(DP_pipe02[4]), .ZN(DP_mult_218_n1669) );
  OAI22_X1 DP_mult_218_U1928 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1668), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1669), .ZN(DP_mult_218_n2143)
         );
  AOI221_X1 DP_mult_218_U1927 ( .B1(DP_pipe02[6]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[5]), .C2(DP_mult_218_n1563), .A(DP_mult_218_n2143), .ZN(
        DP_mult_218_n2142) );
  XNOR2_X1 DP_mult_218_U1926 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2142), 
        .ZN(DP_mult_218_n2140) );
  INV_X1 DP_mult_218_U1925 ( .A(DP_mult_218_n680), .ZN(DP_mult_218_n2141) );
  OAI222_X1 DP_mult_218_U1924 ( .A1(DP_mult_218_n2139), .A2(DP_mult_218_n2140), 
        .B1(DP_mult_218_n2139), .B2(DP_mult_218_n2141), .C1(DP_mult_218_n2141), 
        .C2(DP_mult_218_n2140), .ZN(DP_mult_218_n2135) );
  INV_X1 DP_mult_218_U1923 ( .A(DP_mult_218_n1391), .ZN(DP_mult_218_n1672) );
  INV_X1 DP_mult_218_U1922 ( .A(DP_pipe02[5]), .ZN(DP_mult_218_n1673) );
  OAI22_X1 DP_mult_218_U1921 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1672), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1673), .ZN(DP_mult_218_n2138)
         );
  AOI221_X1 DP_mult_218_U1920 ( .B1(DP_pipe02[7]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[6]), .C2(DP_mult_218_n1563), .A(DP_mult_218_n2138), .ZN(
        DP_mult_218_n2137) );
  XNOR2_X1 DP_mult_218_U1919 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2137), 
        .ZN(DP_mult_218_n2136) );
  AOI222_X1 DP_mult_218_U1918 ( .A1(DP_mult_218_n2135), .A2(DP_mult_218_n2136), 
        .B1(DP_mult_218_n2135), .B2(DP_mult_218_n676), .C1(DP_mult_218_n676), 
        .C2(DP_mult_218_n2136), .ZN(DP_mult_218_n2130) );
  INV_X1 DP_mult_218_U1917 ( .A(DP_mult_218_n1390), .ZN(DP_mult_218_n1676) );
  INV_X1 DP_mult_218_U1916 ( .A(DP_pipe02[6]), .ZN(DP_mult_218_n1677) );
  OAI22_X1 DP_mult_218_U1915 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1676), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1677), .ZN(DP_mult_218_n2134)
         );
  AOI221_X1 DP_mult_218_U1914 ( .B1(DP_pipe02[8]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[7]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2134), .ZN(
        DP_mult_218_n2133) );
  XNOR2_X1 DP_mult_218_U1913 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2133), 
        .ZN(DP_mult_218_n2131) );
  INV_X1 DP_mult_218_U1912 ( .A(DP_mult_218_n672), .ZN(DP_mult_218_n2132) );
  OAI222_X1 DP_mult_218_U1911 ( .A1(DP_mult_218_n2130), .A2(DP_mult_218_n2131), 
        .B1(DP_mult_218_n2130), .B2(DP_mult_218_n2132), .C1(DP_mult_218_n2132), 
        .C2(DP_mult_218_n2131), .ZN(DP_mult_218_n2126) );
  INV_X1 DP_mult_218_U1910 ( .A(DP_mult_218_n1389), .ZN(DP_mult_218_n1680) );
  INV_X1 DP_mult_218_U1909 ( .A(DP_pipe02[7]), .ZN(DP_mult_218_n1681) );
  OAI22_X1 DP_mult_218_U1908 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1680), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1681), .ZN(DP_mult_218_n2129)
         );
  AOI221_X1 DP_mult_218_U1907 ( .B1(DP_pipe02[9]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[8]), .C2(DP_mult_218_n1563), .A(DP_mult_218_n2129), .ZN(
        DP_mult_218_n2128) );
  XNOR2_X1 DP_mult_218_U1906 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2128), 
        .ZN(DP_mult_218_n2127) );
  AOI222_X1 DP_mult_218_U1905 ( .A1(DP_mult_218_n2126), .A2(DP_mult_218_n2127), 
        .B1(DP_mult_218_n2126), .B2(DP_mult_218_n666), .C1(DP_mult_218_n666), 
        .C2(DP_mult_218_n2127), .ZN(DP_mult_218_n2121) );
  INV_X1 DP_mult_218_U1904 ( .A(DP_mult_218_n1388), .ZN(DP_mult_218_n1684) );
  INV_X1 DP_mult_218_U1903 ( .A(DP_pipe02[8]), .ZN(DP_mult_218_n1685) );
  OAI22_X1 DP_mult_218_U1902 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1684), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1685), .ZN(DP_mult_218_n2125)
         );
  AOI221_X1 DP_mult_218_U1901 ( .B1(DP_pipe02[10]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[9]), .C2(DP_mult_218_n1563), .A(DP_mult_218_n2125), .ZN(
        DP_mult_218_n2124) );
  XNOR2_X1 DP_mult_218_U1900 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2124), 
        .ZN(DP_mult_218_n2122) );
  INV_X1 DP_mult_218_U1899 ( .A(DP_mult_218_n660), .ZN(DP_mult_218_n2123) );
  OAI222_X1 DP_mult_218_U1898 ( .A1(DP_mult_218_n2121), .A2(DP_mult_218_n2122), 
        .B1(DP_mult_218_n2121), .B2(DP_mult_218_n2123), .C1(DP_mult_218_n2123), 
        .C2(DP_mult_218_n2122), .ZN(DP_mult_218_n2117) );
  INV_X1 DP_mult_218_U1897 ( .A(DP_mult_218_n1387), .ZN(DP_mult_218_n1688) );
  INV_X1 DP_mult_218_U1896 ( .A(DP_pipe02[9]), .ZN(DP_mult_218_n1689) );
  OAI22_X1 DP_mult_218_U1895 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1688), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1689), .ZN(DP_mult_218_n2120)
         );
  AOI221_X1 DP_mult_218_U1894 ( .B1(DP_pipe02[11]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[10]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2120), 
        .ZN(DP_mult_218_n2119) );
  XNOR2_X1 DP_mult_218_U1893 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2119), 
        .ZN(DP_mult_218_n2118) );
  AOI222_X1 DP_mult_218_U1892 ( .A1(DP_mult_218_n2117), .A2(DP_mult_218_n2118), 
        .B1(DP_mult_218_n2117), .B2(DP_mult_218_n654), .C1(DP_mult_218_n654), 
        .C2(DP_mult_218_n2118), .ZN(DP_mult_218_n2112) );
  INV_X1 DP_mult_218_U1891 ( .A(DP_mult_218_n1386), .ZN(DP_mult_218_n1692) );
  INV_X1 DP_mult_218_U1890 ( .A(DP_pipe02[10]), .ZN(DP_mult_218_n1693) );
  OAI22_X1 DP_mult_218_U1889 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1692), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1693), .ZN(DP_mult_218_n2116)
         );
  AOI221_X1 DP_mult_218_U1888 ( .B1(DP_pipe02[12]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[11]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2116), 
        .ZN(DP_mult_218_n2115) );
  XNOR2_X1 DP_mult_218_U1887 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2115), 
        .ZN(DP_mult_218_n2113) );
  INV_X1 DP_mult_218_U1886 ( .A(DP_mult_218_n646), .ZN(DP_mult_218_n2114) );
  OAI222_X1 DP_mult_218_U1885 ( .A1(DP_mult_218_n2112), .A2(DP_mult_218_n2113), 
        .B1(DP_mult_218_n2112), .B2(DP_mult_218_n2114), .C1(DP_mult_218_n2114), 
        .C2(DP_mult_218_n2113), .ZN(DP_mult_218_n2108) );
  INV_X1 DP_mult_218_U1884 ( .A(DP_mult_218_n1385), .ZN(DP_mult_218_n1696) );
  INV_X1 DP_mult_218_U1883 ( .A(DP_pipe02[11]), .ZN(DP_mult_218_n1697) );
  OAI22_X1 DP_mult_218_U1882 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1696), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1697), .ZN(DP_mult_218_n2111)
         );
  AOI221_X1 DP_mult_218_U1881 ( .B1(DP_pipe02[13]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[12]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2111), 
        .ZN(DP_mult_218_n2110) );
  XNOR2_X1 DP_mult_218_U1880 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2110), 
        .ZN(DP_mult_218_n2109) );
  AOI222_X1 DP_mult_218_U1879 ( .A1(DP_mult_218_n2108), .A2(DP_mult_218_n2109), 
        .B1(DP_mult_218_n2108), .B2(DP_mult_218_n638), .C1(DP_mult_218_n638), 
        .C2(DP_mult_218_n2109), .ZN(DP_mult_218_n2103) );
  INV_X1 DP_mult_218_U1878 ( .A(DP_mult_218_n1384), .ZN(DP_mult_218_n1700) );
  INV_X1 DP_mult_218_U1877 ( .A(DP_pipe02[12]), .ZN(DP_mult_218_n1701) );
  OAI22_X1 DP_mult_218_U1876 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1700), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1701), .ZN(DP_mult_218_n2107)
         );
  AOI221_X1 DP_mult_218_U1875 ( .B1(DP_pipe02[14]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[13]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2107), 
        .ZN(DP_mult_218_n2106) );
  XNOR2_X1 DP_mult_218_U1874 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2106), 
        .ZN(DP_mult_218_n2104) );
  INV_X1 DP_mult_218_U1873 ( .A(DP_mult_218_n630), .ZN(DP_mult_218_n2105) );
  OAI222_X1 DP_mult_218_U1872 ( .A1(DP_mult_218_n2103), .A2(DP_mult_218_n2104), 
        .B1(DP_mult_218_n2103), .B2(DP_mult_218_n2105), .C1(DP_mult_218_n2105), 
        .C2(DP_mult_218_n2104), .ZN(DP_mult_218_n2099) );
  INV_X1 DP_mult_218_U1871 ( .A(DP_mult_218_n1383), .ZN(DP_mult_218_n1704) );
  INV_X1 DP_mult_218_U1870 ( .A(DP_pipe02[13]), .ZN(DP_mult_218_n1705) );
  OAI22_X1 DP_mult_218_U1869 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1704), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1705), .ZN(DP_mult_218_n2102)
         );
  AOI221_X1 DP_mult_218_U1868 ( .B1(DP_pipe02[15]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[14]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2102), 
        .ZN(DP_mult_218_n2101) );
  XNOR2_X1 DP_mult_218_U1867 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2101), 
        .ZN(DP_mult_218_n2100) );
  AOI222_X1 DP_mult_218_U1866 ( .A1(DP_mult_218_n2099), .A2(DP_mult_218_n2100), 
        .B1(DP_mult_218_n2099), .B2(DP_mult_218_n620), .C1(DP_mult_218_n620), 
        .C2(DP_mult_218_n2100), .ZN(DP_mult_218_n2094) );
  INV_X1 DP_mult_218_U1865 ( .A(DP_mult_218_n1382), .ZN(DP_mult_218_n1708) );
  INV_X1 DP_mult_218_U1864 ( .A(DP_pipe02[14]), .ZN(DP_mult_218_n1709) );
  OAI22_X1 DP_mult_218_U1863 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1708), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1709), .ZN(DP_mult_218_n2098)
         );
  AOI221_X1 DP_mult_218_U1862 ( .B1(DP_pipe02[16]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[15]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2098), 
        .ZN(DP_mult_218_n2097) );
  XNOR2_X1 DP_mult_218_U1861 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2097), 
        .ZN(DP_mult_218_n2095) );
  INV_X1 DP_mult_218_U1860 ( .A(DP_mult_218_n610), .ZN(DP_mult_218_n2096) );
  OAI222_X1 DP_mult_218_U1859 ( .A1(DP_mult_218_n2094), .A2(DP_mult_218_n2095), 
        .B1(DP_mult_218_n2094), .B2(DP_mult_218_n2096), .C1(DP_mult_218_n2096), 
        .C2(DP_mult_218_n2095), .ZN(DP_mult_218_n2090) );
  INV_X1 DP_mult_218_U1858 ( .A(DP_mult_218_n1381), .ZN(DP_mult_218_n1712) );
  INV_X1 DP_mult_218_U1857 ( .A(DP_pipe02[15]), .ZN(DP_mult_218_n1713) );
  OAI22_X1 DP_mult_218_U1856 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1712), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1713), .ZN(DP_mult_218_n2093)
         );
  AOI221_X1 DP_mult_218_U1855 ( .B1(DP_pipe02[17]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[16]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2093), 
        .ZN(DP_mult_218_n2092) );
  XNOR2_X1 DP_mult_218_U1854 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2092), 
        .ZN(DP_mult_218_n2091) );
  AOI222_X1 DP_mult_218_U1853 ( .A1(DP_mult_218_n2090), .A2(DP_mult_218_n2091), 
        .B1(DP_mult_218_n2090), .B2(DP_mult_218_n600), .C1(DP_mult_218_n600), 
        .C2(DP_mult_218_n2091), .ZN(DP_mult_218_n2085) );
  INV_X1 DP_mult_218_U1852 ( .A(DP_mult_218_n1380), .ZN(DP_mult_218_n1716) );
  INV_X1 DP_mult_218_U1851 ( .A(DP_pipe02[16]), .ZN(DP_mult_218_n1717) );
  OAI22_X1 DP_mult_218_U1850 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1716), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1717), .ZN(DP_mult_218_n2089)
         );
  AOI221_X1 DP_mult_218_U1849 ( .B1(DP_pipe02[18]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[17]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2089), 
        .ZN(DP_mult_218_n2088) );
  XNOR2_X1 DP_mult_218_U1848 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2088), 
        .ZN(DP_mult_218_n2086) );
  INV_X1 DP_mult_218_U1847 ( .A(DP_mult_218_n588), .ZN(DP_mult_218_n2087) );
  OAI222_X1 DP_mult_218_U1846 ( .A1(DP_mult_218_n2085), .A2(DP_mult_218_n2086), 
        .B1(DP_mult_218_n2085), .B2(DP_mult_218_n2087), .C1(DP_mult_218_n2087), 
        .C2(DP_mult_218_n2086), .ZN(DP_mult_218_n2081) );
  INV_X1 DP_mult_218_U1845 ( .A(DP_mult_218_n1379), .ZN(DP_mult_218_n1720) );
  INV_X1 DP_mult_218_U1844 ( .A(DP_pipe02[17]), .ZN(DP_mult_218_n1721) );
  OAI22_X1 DP_mult_218_U1843 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1720), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1721), .ZN(DP_mult_218_n2084)
         );
  AOI221_X1 DP_mult_218_U1842 ( .B1(DP_pipe02[19]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[18]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2084), 
        .ZN(DP_mult_218_n2083) );
  XNOR2_X1 DP_mult_218_U1841 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2083), 
        .ZN(DP_mult_218_n2082) );
  AOI222_X1 DP_mult_218_U1840 ( .A1(DP_mult_218_n2081), .A2(DP_mult_218_n2082), 
        .B1(DP_mult_218_n2081), .B2(DP_mult_218_n576), .C1(DP_mult_218_n576), 
        .C2(DP_mult_218_n2082), .ZN(DP_mult_218_n2080) );
  INV_X1 DP_mult_218_U1839 ( .A(DP_mult_218_n2080), .ZN(DP_mult_218_n2076) );
  INV_X1 DP_mult_218_U1838 ( .A(DP_mult_218_n1378), .ZN(DP_mult_218_n1724) );
  INV_X1 DP_mult_218_U1837 ( .A(DP_pipe02[18]), .ZN(DP_mult_218_n1725) );
  OAI22_X1 DP_mult_218_U1836 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1724), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1725), .ZN(DP_mult_218_n2079)
         );
  AOI221_X1 DP_mult_218_U1835 ( .B1(DP_pipe02[20]), .B2(DP_mult_218_n1561), 
        .C1(DP_pipe02[19]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2079), 
        .ZN(DP_mult_218_n2078) );
  XNOR2_X1 DP_mult_218_U1834 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n2078), 
        .ZN(DP_mult_218_n2077) );
  AOI222_X1 DP_mult_218_U1833 ( .A1(DP_mult_218_n2076), .A2(DP_mult_218_n2077), 
        .B1(DP_mult_218_n2076), .B2(DP_mult_218_n564), .C1(DP_mult_218_n564), 
        .C2(DP_mult_218_n2077), .ZN(DP_mult_218_n2071) );
  INV_X1 DP_mult_218_U1832 ( .A(DP_mult_218_n1377), .ZN(DP_mult_218_n1728) );
  INV_X1 DP_mult_218_U1831 ( .A(DP_pipe02[19]), .ZN(DP_mult_218_n1729) );
  OAI22_X1 DP_mult_218_U1830 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1728), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1729), .ZN(DP_mult_218_n2075)
         );
  AOI221_X1 DP_mult_218_U1829 ( .B1(DP_mult_218_n1561), .B2(DP_pipe02[21]), 
        .C1(DP_pipe02[20]), .C2(DP_mult_218_n1562), .A(DP_mult_218_n2075), 
        .ZN(DP_mult_218_n2074) );
  XNOR2_X1 DP_mult_218_U1828 ( .A(DP_mult_218_n1742), .B(DP_mult_218_n2074), 
        .ZN(DP_mult_218_n2072) );
  INV_X1 DP_mult_218_U1827 ( .A(DP_mult_218_n550), .ZN(DP_mult_218_n2073) );
  OAI222_X1 DP_mult_218_U1826 ( .A1(DP_mult_218_n2071), .A2(DP_mult_218_n2072), 
        .B1(DP_mult_218_n2071), .B2(DP_mult_218_n2073), .C1(DP_mult_218_n2073), 
        .C2(DP_mult_218_n2072), .ZN(DP_mult_218_n326) );
  XNOR2_X1 DP_mult_218_U1825 ( .A(DP_coeff_pipe02[21]), .B(DP_mult_218_n1608), 
        .ZN(DP_mult_218_n2067) );
  INV_X1 DP_mult_218_U1824 ( .A(DP_mult_218_n2067), .ZN(DP_mult_218_n2070) );
  XNOR2_X1 DP_mult_218_U1823 ( .A(DP_coeff_pipe02[21]), .B(DP_coeff_pipe02[22]), .ZN(DP_mult_218_n2069) );
  XNOR2_X1 DP_mult_218_U1822 ( .A(DP_coeff_pipe02[22]), .B(DP_mult_218_n1611), 
        .ZN(DP_mult_218_n2068) );
  NAND3_X1 DP_mult_218_U1821 ( .A1(DP_mult_218_n2067), .A2(DP_mult_218_n2068), 
        .A3(DP_mult_218_n2069), .ZN(DP_mult_218_n1629) );
  INV_X1 DP_mult_218_U1820 ( .A(DP_pipe02[21]), .ZN(DP_mult_218_n1643) );
  OAI22_X1 DP_mult_218_U1819 ( .A1(DP_mult_218_n1544), .A2(DP_mult_218_n1619), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1643), .ZN(DP_mult_218_n2066)
         );
  AOI221_X1 DP_mult_218_U1818 ( .B1(DP_pipe02[22]), .B2(DP_mult_218_n1560), 
        .C1(DP_mult_218_n1375), .C2(DP_mult_218_n1553), .A(DP_mult_218_n2066), 
        .ZN(DP_mult_218_n2065) );
  XOR2_X1 DP_mult_218_U1817 ( .A(DP_mult_218_n1611), .B(DP_mult_218_n2065), 
        .Z(DP_mult_218_n1627) );
  INV_X1 DP_mult_218_U1816 ( .A(DP_mult_218_n1627), .ZN(DP_mult_218_n351) );
  INV_X1 DP_mult_218_U1815 ( .A(DP_mult_218_n356), .ZN(DP_mult_218_n360) );
  OAI22_X1 DP_mult_218_U1814 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1712), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1713), .ZN(DP_mult_218_n2064)
         );
  AOI221_X1 DP_mult_218_U1813 ( .B1(DP_pipe02[17]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[16]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2064), 
        .ZN(DP_mult_218_n2063) );
  XOR2_X1 DP_mult_218_U1812 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2063), 
        .Z(DP_mult_218_n374) );
  INV_X1 DP_mult_218_U1811 ( .A(DP_mult_218_n374), .ZN(DP_mult_218_n368) );
  INV_X1 DP_mult_218_U1810 ( .A(DP_mult_218_n387), .ZN(DP_mult_218_n395) );
  OAI22_X1 DP_mult_218_U1809 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1688), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1689), .ZN(DP_mult_218_n2062)
         );
  AOI221_X1 DP_mult_218_U1808 ( .B1(DP_pipe02[11]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[10]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2062), 
        .ZN(DP_mult_218_n2061) );
  XOR2_X1 DP_mult_218_U1807 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2061), 
        .Z(DP_mult_218_n421) );
  INV_X1 DP_mult_218_U1806 ( .A(DP_mult_218_n421), .ZN(DP_mult_218_n411) );
  OAI22_X1 DP_mult_218_U1805 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1676), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1677), .ZN(DP_mult_218_n2060)
         );
  AOI221_X1 DP_mult_218_U1804 ( .B1(DP_pipe02[8]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[7]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2060), .ZN(
        DP_mult_218_n2059) );
  XOR2_X1 DP_mult_218_U1803 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2059), 
        .Z(DP_mult_218_n454) );
  INV_X1 DP_mult_218_U1802 ( .A(DP_mult_218_n454), .ZN(DP_mult_218_n442) );
  OAI21_X1 DP_mult_218_U1801 ( .B1(DP_mult_218_n1561), .B2(DP_mult_218_n1563), 
        .A(DP_mult_218_n1615), .ZN(DP_mult_218_n2058) );
  OAI221_X1 DP_mult_218_U1800 ( .B1(DP_mult_218_n1619), .B2(DP_mult_218_n1639), 
        .C1(DP_mult_218_n1620), .C2(DP_mult_218_n1564), .A(DP_mult_218_n2058), 
        .ZN(DP_mult_218_n2057) );
  XOR2_X1 DP_mult_218_U1799 ( .A(DP_mult_218_n2057), .B(DP_mult_218_n1742), 
        .Z(DP_mult_218_n2056) );
  NOR2_X1 DP_mult_218_U1798 ( .A1(DP_mult_218_n2056), .A2(DP_mult_218_n519), 
        .ZN(DP_mult_218_n493) );
  INV_X1 DP_mult_218_U1797 ( .A(DP_mult_218_n493), .ZN(DP_mult_218_n479) );
  XNOR2_X1 DP_mult_218_U1796 ( .A(DP_mult_218_n519), .B(DP_mult_218_n2056), 
        .ZN(DP_mult_218_n506) );
  INV_X1 DP_mult_218_U1795 ( .A(DP_pipe02[20]), .ZN(DP_mult_218_n1640) );
  OAI22_X1 DP_mult_218_U1794 ( .A1(DP_mult_218_n1556), .A2(DP_mult_218_n1640), 
        .B1(DP_mult_218_n1550), .B2(DP_mult_218_n1643), .ZN(DP_mult_218_n2055)
         );
  AOI221_X1 DP_mult_218_U1793 ( .B1(DP_pipe02[22]), .B2(DP_mult_218_n1559), 
        .C1(DP_mult_218_n1376), .C2(DP_mult_218_n1553), .A(DP_mult_218_n2055), 
        .ZN(DP_mult_218_n2054) );
  XNOR2_X1 DP_mult_218_U1792 ( .A(DP_coeff_pipe02[23]), .B(DP_mult_218_n2054), 
        .ZN(DP_mult_218_n729) );
  OAI22_X1 DP_mult_218_U1791 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1728), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1729), .ZN(DP_mult_218_n2053)
         );
  AOI221_X1 DP_mult_218_U1790 ( .B1(DP_pipe02[21]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[20]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2053), 
        .ZN(DP_mult_218_n2052) );
  XNOR2_X1 DP_mult_218_U1789 ( .A(DP_coeff_pipe02[23]), .B(DP_mult_218_n2052), 
        .ZN(DP_mult_218_n730) );
  OAI22_X1 DP_mult_218_U1788 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1724), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1725), .ZN(DP_mult_218_n2051)
         );
  AOI221_X1 DP_mult_218_U1787 ( .B1(DP_pipe02[20]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[19]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2051), 
        .ZN(DP_mult_218_n2050) );
  XNOR2_X1 DP_mult_218_U1786 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2050), 
        .ZN(DP_mult_218_n731) );
  OAI22_X1 DP_mult_218_U1785 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1720), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1721), .ZN(DP_mult_218_n2049)
         );
  AOI221_X1 DP_mult_218_U1784 ( .B1(DP_pipe02[19]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[18]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2049), 
        .ZN(DP_mult_218_n2048) );
  XNOR2_X1 DP_mult_218_U1783 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2048), 
        .ZN(DP_mult_218_n732) );
  OAI22_X1 DP_mult_218_U1782 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1716), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1717), .ZN(DP_mult_218_n2047)
         );
  AOI221_X1 DP_mult_218_U1781 ( .B1(DP_pipe02[18]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[17]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2047), 
        .ZN(DP_mult_218_n2046) );
  XNOR2_X1 DP_mult_218_U1780 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2046), 
        .ZN(DP_mult_218_n733) );
  OAI22_X1 DP_mult_218_U1779 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1708), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1709), .ZN(DP_mult_218_n2045)
         );
  AOI221_X1 DP_mult_218_U1778 ( .B1(DP_pipe02[16]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[15]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2045), 
        .ZN(DP_mult_218_n2044) );
  XNOR2_X1 DP_mult_218_U1777 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2044), 
        .ZN(DP_mult_218_n734) );
  OAI22_X1 DP_mult_218_U1776 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1704), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1705), .ZN(DP_mult_218_n2043)
         );
  AOI221_X1 DP_mult_218_U1775 ( .B1(DP_pipe02[15]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[14]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2043), 
        .ZN(DP_mult_218_n2042) );
  XNOR2_X1 DP_mult_218_U1774 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2042), 
        .ZN(DP_mult_218_n735) );
  OAI22_X1 DP_mult_218_U1773 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1700), 
        .B1(DP_mult_218_n1556), .B2(DP_mult_218_n1701), .ZN(DP_mult_218_n2041)
         );
  AOI221_X1 DP_mult_218_U1772 ( .B1(DP_pipe02[14]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[13]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2041), 
        .ZN(DP_mult_218_n2040) );
  XNOR2_X1 DP_mult_218_U1771 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2040), 
        .ZN(DP_mult_218_n736) );
  OAI22_X1 DP_mult_218_U1770 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1696), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1697), .ZN(DP_mult_218_n2039)
         );
  AOI221_X1 DP_mult_218_U1769 ( .B1(DP_pipe02[13]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[12]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2039), 
        .ZN(DP_mult_218_n2038) );
  XNOR2_X1 DP_mult_218_U1768 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2038), 
        .ZN(DP_mult_218_n737) );
  OAI22_X1 DP_mult_218_U1767 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1692), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1693), .ZN(DP_mult_218_n2037)
         );
  AOI221_X1 DP_mult_218_U1766 ( .B1(DP_pipe02[12]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[11]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2037), 
        .ZN(DP_mult_218_n2036) );
  XNOR2_X1 DP_mult_218_U1765 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2036), 
        .ZN(DP_mult_218_n738) );
  OAI22_X1 DP_mult_218_U1764 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1684), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1685), .ZN(DP_mult_218_n2035)
         );
  AOI221_X1 DP_mult_218_U1763 ( .B1(DP_pipe02[10]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[9]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2035), .ZN(
        DP_mult_218_n2034) );
  XNOR2_X1 DP_mult_218_U1762 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2034), 
        .ZN(DP_mult_218_n739) );
  OAI22_X1 DP_mult_218_U1761 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1680), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1681), .ZN(DP_mult_218_n2033)
         );
  AOI221_X1 DP_mult_218_U1760 ( .B1(DP_pipe02[9]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[8]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2033), .ZN(
        DP_mult_218_n2032) );
  XNOR2_X1 DP_mult_218_U1759 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2032), 
        .ZN(DP_mult_218_n740) );
  OAI22_X1 DP_mult_218_U1758 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1672), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1673), .ZN(DP_mult_218_n2031)
         );
  AOI221_X1 DP_mult_218_U1757 ( .B1(DP_pipe02[7]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[6]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2031), .ZN(
        DP_mult_218_n2030) );
  XNOR2_X1 DP_mult_218_U1756 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2030), 
        .ZN(DP_mult_218_n741) );
  OAI22_X1 DP_mult_218_U1755 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1668), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1669), .ZN(DP_mult_218_n2029)
         );
  AOI221_X1 DP_mult_218_U1754 ( .B1(DP_pipe02[6]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[5]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2029), .ZN(
        DP_mult_218_n2028) );
  XNOR2_X1 DP_mult_218_U1753 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2028), 
        .ZN(DP_mult_218_n742) );
  OAI22_X1 DP_mult_218_U1752 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1664), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1665), .ZN(DP_mult_218_n2027)
         );
  AOI221_X1 DP_mult_218_U1751 ( .B1(DP_pipe02[5]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[4]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2027), .ZN(
        DP_mult_218_n2026) );
  XNOR2_X1 DP_mult_218_U1750 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2026), 
        .ZN(DP_mult_218_n743) );
  OAI22_X1 DP_mult_218_U1749 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1660), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1661), .ZN(DP_mult_218_n2025)
         );
  AOI221_X1 DP_mult_218_U1748 ( .B1(DP_pipe02[4]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[3]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2025), .ZN(
        DP_mult_218_n2024) );
  XNOR2_X1 DP_mult_218_U1747 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2024), 
        .ZN(DP_mult_218_n744) );
  OAI22_X1 DP_mult_218_U1746 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1657), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1649), .ZN(DP_mult_218_n2023)
         );
  AOI221_X1 DP_mult_218_U1745 ( .B1(DP_pipe02[3]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[2]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2023), .ZN(
        DP_mult_218_n2022) );
  XNOR2_X1 DP_mult_218_U1744 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2022), 
        .ZN(DP_mult_218_n745) );
  INV_X1 DP_mult_218_U1743 ( .A(DP_mult_218_n1396), .ZN(DP_mult_218_n1653) );
  INV_X1 DP_mult_218_U1742 ( .A(DP_pipe02[0]), .ZN(DP_mult_218_n1647) );
  OAI22_X1 DP_mult_218_U1741 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1653), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1567), .ZN(DP_mult_218_n2021)
         );
  AOI221_X1 DP_mult_218_U1740 ( .B1(DP_pipe02[2]), .B2(DP_mult_218_n1559), 
        .C1(DP_pipe02[1]), .C2(DP_mult_218_n1560), .A(DP_mult_218_n2021), .ZN(
        DP_mult_218_n2020) );
  XNOR2_X1 DP_mult_218_U1739 ( .A(DP_mult_218_n1610), .B(DP_mult_218_n2020), 
        .ZN(DP_mult_218_n746) );
  OAI222_X1 DP_mult_218_U1738 ( .A1(DP_mult_218_n1544), .A2(DP_mult_218_n1649), 
        .B1(DP_mult_218_n1550), .B2(DP_mult_218_n1566), .C1(DP_mult_218_n1558), 
        .C2(DP_mult_218_n1650), .ZN(DP_mult_218_n2019) );
  XNOR2_X1 DP_mult_218_U1737 ( .A(DP_mult_218_n2019), .B(DP_mult_218_n1611), 
        .ZN(DP_mult_218_n747) );
  OAI22_X1 DP_mult_218_U1736 ( .A1(DP_mult_218_n1544), .A2(DP_mult_218_n1567), 
        .B1(DP_mult_218_n1558), .B2(DP_mult_218_n1567), .ZN(DP_mult_218_n2018)
         );
  XNOR2_X1 DP_mult_218_U1735 ( .A(DP_mult_218_n2018), .B(DP_mult_218_n1611), 
        .ZN(DP_mult_218_n748) );
  XOR2_X1 DP_mult_218_U1734 ( .A(DP_coeff_pipe02[18]), .B(DP_mult_218_n1607), 
        .Z(DP_mult_218_n2017) );
  XOR2_X1 DP_mult_218_U1733 ( .A(DP_coeff_pipe02[19]), .B(DP_mult_218_n1608), 
        .Z(DP_mult_218_n2016) );
  XNOR2_X1 DP_mult_218_U1732 ( .A(DP_coeff_pipe02[18]), .B(DP_coeff_pipe02[19]), .ZN(DP_mult_218_n2015) );
  NAND3_X1 DP_mult_218_U1731 ( .A1(DP_mult_218_n2017), .A2(DP_mult_218_n2016), 
        .A3(DP_mult_218_n2015), .ZN(DP_mult_218_n1967) );
  INV_X1 DP_mult_218_U1730 ( .A(DP_mult_218_n2017), .ZN(DP_mult_218_n2014) );
  OAI21_X1 DP_mult_218_U1729 ( .B1(DP_mult_218_n1594), .B2(DP_mult_218_n1595), 
        .A(DP_mult_218_n1615), .ZN(DP_mult_218_n2013) );
  OAI221_X1 DP_mult_218_U1728 ( .B1(DP_mult_218_n1617), .B2(DP_mult_218_n1597), 
        .C1(DP_mult_218_n1620), .C2(DP_mult_218_n1593), .A(DP_mult_218_n2013), 
        .ZN(DP_mult_218_n2012) );
  XNOR2_X1 DP_mult_218_U1727 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n2012), 
        .ZN(DP_mult_218_n749) );
  INV_X1 DP_mult_218_U1726 ( .A(DP_mult_218_n1374), .ZN(DP_mult_218_n1633) );
  INV_X1 DP_mult_218_U1725 ( .A(DP_pipe02[22]), .ZN(DP_mult_218_n1634) );
  OAI22_X1 DP_mult_218_U1724 ( .A1(DP_mult_218_n1633), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1634), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n2011)
         );
  AOI221_X1 DP_mult_218_U1723 ( .B1(DP_mult_218_n1594), .B2(DP_mult_218_n1614), 
        .C1(DP_mult_218_n1595), .C2(DP_mult_218_n1615), .A(DP_mult_218_n2011), 
        .ZN(DP_mult_218_n2010) );
  XNOR2_X1 DP_mult_218_U1722 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n2010), 
        .ZN(DP_mult_218_n750) );
  OAI22_X1 DP_mult_218_U1721 ( .A1(DP_mult_218_n1617), .A2(DP_mult_218_n1543), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n2009)
         );
  AOI221_X1 DP_mult_218_U1720 ( .B1(DP_mult_218_n1595), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1547), .C2(DP_mult_218_n1375), .A(DP_mult_218_n2009), 
        .ZN(DP_mult_218_n2008) );
  XNOR2_X1 DP_mult_218_U1719 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n2008), 
        .ZN(DP_mult_218_n751) );
  OAI22_X1 DP_mult_218_U1718 ( .A1(DP_mult_218_n1640), .A2(DP_mult_218_n1597), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1552), .ZN(DP_mult_218_n2007)
         );
  AOI221_X1 DP_mult_218_U1717 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1547), .C2(DP_mult_218_n1376), .A(DP_mult_218_n2007), 
        .ZN(DP_mult_218_n2006) );
  XNOR2_X1 DP_mult_218_U1716 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n2006), 
        .ZN(DP_mult_218_n752) );
  OAI22_X1 DP_mult_218_U1715 ( .A1(DP_mult_218_n1728), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1729), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n2005)
         );
  AOI221_X1 DP_mult_218_U1714 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[21]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[20]), .A(DP_mult_218_n2005), 
        .ZN(DP_mult_218_n2004) );
  XNOR2_X1 DP_mult_218_U1713 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n2004), 
        .ZN(DP_mult_218_n753) );
  OAI22_X1 DP_mult_218_U1712 ( .A1(DP_mult_218_n1724), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1725), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n2003)
         );
  AOI221_X1 DP_mult_218_U1711 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[20]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[19]), .A(DP_mult_218_n2003), 
        .ZN(DP_mult_218_n2002) );
  XNOR2_X1 DP_mult_218_U1710 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n2002), 
        .ZN(DP_mult_218_n754) );
  OAI22_X1 DP_mult_218_U1709 ( .A1(DP_mult_218_n1720), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1721), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n2001)
         );
  AOI221_X1 DP_mult_218_U1708 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[19]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[18]), .A(DP_mult_218_n2001), 
        .ZN(DP_mult_218_n2000) );
  XNOR2_X1 DP_mult_218_U1707 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n2000), 
        .ZN(DP_mult_218_n755) );
  OAI22_X1 DP_mult_218_U1706 ( .A1(DP_mult_218_n1716), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1717), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n1999)
         );
  AOI221_X1 DP_mult_218_U1705 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[18]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[17]), .A(DP_mult_218_n1999), 
        .ZN(DP_mult_218_n1998) );
  XNOR2_X1 DP_mult_218_U1704 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n1998), 
        .ZN(DP_mult_218_n756) );
  OAI22_X1 DP_mult_218_U1703 ( .A1(DP_mult_218_n1712), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1713), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n1997)
         );
  AOI221_X1 DP_mult_218_U1702 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[17]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[16]), .A(DP_mult_218_n1997), 
        .ZN(DP_mult_218_n1996) );
  XNOR2_X1 DP_mult_218_U1701 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n1996), 
        .ZN(DP_mult_218_n757) );
  OAI22_X1 DP_mult_218_U1700 ( .A1(DP_mult_218_n1708), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1709), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n1995)
         );
  AOI221_X1 DP_mult_218_U1699 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[16]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[15]), .A(DP_mult_218_n1995), 
        .ZN(DP_mult_218_n1994) );
  XNOR2_X1 DP_mult_218_U1698 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n1994), 
        .ZN(DP_mult_218_n758) );
  OAI22_X1 DP_mult_218_U1697 ( .A1(DP_mult_218_n1704), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1705), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n1993)
         );
  AOI221_X1 DP_mult_218_U1696 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[15]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[14]), .A(DP_mult_218_n1993), 
        .ZN(DP_mult_218_n1992) );
  XNOR2_X1 DP_mult_218_U1695 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n1992), 
        .ZN(DP_mult_218_n759) );
  OAI22_X1 DP_mult_218_U1694 ( .A1(DP_mult_218_n1700), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1701), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n1991)
         );
  AOI221_X1 DP_mult_218_U1693 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[14]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[13]), .A(DP_mult_218_n1991), 
        .ZN(DP_mult_218_n1990) );
  XNOR2_X1 DP_mult_218_U1692 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n1990), 
        .ZN(DP_mult_218_n760) );
  OAI22_X1 DP_mult_218_U1691 ( .A1(DP_mult_218_n1696), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1697), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n1989)
         );
  AOI221_X1 DP_mult_218_U1690 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[13]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[12]), .A(DP_mult_218_n1989), 
        .ZN(DP_mult_218_n1988) );
  XNOR2_X1 DP_mult_218_U1689 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n1988), 
        .ZN(DP_mult_218_n761) );
  OAI22_X1 DP_mult_218_U1688 ( .A1(DP_mult_218_n1692), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1693), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1987)
         );
  AOI221_X1 DP_mult_218_U1687 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[12]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[11]), .A(DP_mult_218_n1987), 
        .ZN(DP_mult_218_n1986) );
  XNOR2_X1 DP_mult_218_U1686 ( .A(DP_mult_218_n1609), .B(DP_mult_218_n1986), 
        .ZN(DP_mult_218_n762) );
  OAI22_X1 DP_mult_218_U1685 ( .A1(DP_mult_218_n1688), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1689), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1985)
         );
  AOI221_X1 DP_mult_218_U1684 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[11]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[10]), .A(DP_mult_218_n1985), 
        .ZN(DP_mult_218_n1984) );
  XNOR2_X1 DP_mult_218_U1683 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1984), 
        .ZN(DP_mult_218_n763) );
  OAI22_X1 DP_mult_218_U1682 ( .A1(DP_mult_218_n1684), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1685), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1983)
         );
  AOI221_X1 DP_mult_218_U1681 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[10]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[9]), .A(DP_mult_218_n1983), .ZN(
        DP_mult_218_n1982) );
  XNOR2_X1 DP_mult_218_U1680 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1982), 
        .ZN(DP_mult_218_n764) );
  OAI22_X1 DP_mult_218_U1679 ( .A1(DP_mult_218_n1680), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1681), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1981)
         );
  AOI221_X1 DP_mult_218_U1678 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[9]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[8]), .A(DP_mult_218_n1981), .ZN(
        DP_mult_218_n1980) );
  XNOR2_X1 DP_mult_218_U1677 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1980), 
        .ZN(DP_mult_218_n765) );
  OAI22_X1 DP_mult_218_U1676 ( .A1(DP_mult_218_n1676), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1677), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1979)
         );
  AOI221_X1 DP_mult_218_U1675 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[8]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[7]), .A(DP_mult_218_n1979), .ZN(
        DP_mult_218_n1978) );
  XNOR2_X1 DP_mult_218_U1674 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1978), 
        .ZN(DP_mult_218_n766) );
  OAI22_X1 DP_mult_218_U1673 ( .A1(DP_mult_218_n1672), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1673), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1977)
         );
  AOI221_X1 DP_mult_218_U1672 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[7]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[6]), .A(DP_mult_218_n1977), .ZN(
        DP_mult_218_n1976) );
  XNOR2_X1 DP_mult_218_U1671 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1976), 
        .ZN(DP_mult_218_n767) );
  OAI22_X1 DP_mult_218_U1670 ( .A1(DP_mult_218_n1668), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1669), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1975)
         );
  AOI221_X1 DP_mult_218_U1669 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[6]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[5]), .A(DP_mult_218_n1975), .ZN(
        DP_mult_218_n1974) );
  XNOR2_X1 DP_mult_218_U1668 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1974), 
        .ZN(DP_mult_218_n768) );
  OAI22_X1 DP_mult_218_U1667 ( .A1(DP_mult_218_n1664), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1665), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1973)
         );
  AOI221_X1 DP_mult_218_U1666 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[5]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[4]), .A(DP_mult_218_n1973), .ZN(
        DP_mult_218_n1972) );
  XNOR2_X1 DP_mult_218_U1665 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1972), 
        .ZN(DP_mult_218_n769) );
  OAI22_X1 DP_mult_218_U1664 ( .A1(DP_mult_218_n1660), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1661), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1971)
         );
  AOI221_X1 DP_mult_218_U1663 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[4]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[3]), .A(DP_mult_218_n1971), .ZN(
        DP_mult_218_n1970) );
  XNOR2_X1 DP_mult_218_U1662 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1970), 
        .ZN(DP_mult_218_n770) );
  OAI22_X1 DP_mult_218_U1661 ( .A1(DP_mult_218_n1657), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1649), .B2(DP_mult_218_n1597), .ZN(DP_mult_218_n1969)
         );
  AOI221_X1 DP_mult_218_U1660 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[3]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[2]), .A(DP_mult_218_n1969), .ZN(
        DP_mult_218_n1968) );
  XNOR2_X1 DP_mult_218_U1659 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1968), 
        .ZN(DP_mult_218_n771) );
  OAI22_X1 DP_mult_218_U1658 ( .A1(DP_mult_218_n1653), .A2(DP_mult_218_n1593), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1596), .ZN(DP_mult_218_n1966)
         );
  AOI221_X1 DP_mult_218_U1657 ( .B1(DP_mult_218_n1594), .B2(DP_pipe02[2]), 
        .C1(DP_mult_218_n1595), .C2(DP_pipe02[1]), .A(DP_mult_218_n1966), .ZN(
        DP_mult_218_n1965) );
  XNOR2_X1 DP_mult_218_U1656 ( .A(DP_mult_218_n1608), .B(DP_mult_218_n1965), 
        .ZN(DP_mult_218_n772) );
  OAI222_X1 DP_mult_218_U1655 ( .A1(DP_mult_218_n1649), .A2(DP_mult_218_n1543), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1552), .C1(DP_mult_218_n1650), 
        .C2(DP_mult_218_n1593), .ZN(DP_mult_218_n1964) );
  XOR2_X1 DP_mult_218_U1654 ( .A(DP_mult_218_n1964), .B(DP_mult_218_n1608), 
        .Z(DP_mult_218_n773) );
  OAI22_X1 DP_mult_218_U1653 ( .A1(DP_mult_218_n1565), .A2(DP_mult_218_n1543), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1593), .ZN(DP_mult_218_n1963)
         );
  XOR2_X1 DP_mult_218_U1652 ( .A(DP_mult_218_n1963), .B(DP_mult_218_n1608), 
        .Z(DP_mult_218_n774) );
  XOR2_X1 DP_mult_218_U1651 ( .A(DP_coeff_pipe02[15]), .B(DP_mult_218_n1605), 
        .Z(DP_mult_218_n1962) );
  XNOR2_X1 DP_mult_218_U1650 ( .A(DP_coeff_pipe02[16]), .B(DP_mult_218_n1607), 
        .ZN(DP_mult_218_n1961) );
  XNOR2_X1 DP_mult_218_U1649 ( .A(DP_coeff_pipe02[15]), .B(DP_coeff_pipe02[16]), .ZN(DP_mult_218_n1960) );
  NAND3_X1 DP_mult_218_U1648 ( .A1(DP_mult_218_n1962), .A2(DP_mult_218_n1961), 
        .A3(DP_mult_218_n1960), .ZN(DP_mult_218_n1912) );
  INV_X1 DP_mult_218_U1647 ( .A(DP_mult_218_n1962), .ZN(DP_mult_218_n1959) );
  OAI21_X1 DP_mult_218_U1646 ( .B1(DP_mult_218_n1589), .B2(DP_mult_218_n1590), 
        .A(DP_mult_218_n1615), .ZN(DP_mult_218_n1958) );
  OAI221_X1 DP_mult_218_U1645 ( .B1(DP_mult_218_n1619), .B2(DP_mult_218_n1592), 
        .C1(DP_mult_218_n1617), .C2(DP_mult_218_n1588), .A(DP_mult_218_n1958), 
        .ZN(DP_mult_218_n1957) );
  XNOR2_X1 DP_mult_218_U1644 ( .A(DP_coeff_pipe02[17]), .B(DP_mult_218_n1957), 
        .ZN(DP_mult_218_n775) );
  OAI22_X1 DP_mult_218_U1643 ( .A1(DP_mult_218_n1633), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1634), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1956)
         );
  AOI221_X1 DP_mult_218_U1642 ( .B1(DP_mult_218_n1589), .B2(DP_mult_218_n1614), 
        .C1(DP_mult_218_n1590), .C2(DP_mult_218_n1615), .A(DP_mult_218_n1956), 
        .ZN(DP_mult_218_n1955) );
  XNOR2_X1 DP_mult_218_U1641 ( .A(DP_coeff_pipe02[17]), .B(DP_mult_218_n1955), 
        .ZN(DP_mult_218_n776) );
  OAI22_X1 DP_mult_218_U1640 ( .A1(DP_mult_218_n1617), .A2(DP_mult_218_n1546), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1954)
         );
  AOI221_X1 DP_mult_218_U1639 ( .B1(DP_mult_218_n1590), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1549), .C2(DP_mult_218_n1375), .A(DP_mult_218_n1954), 
        .ZN(DP_mult_218_n1953) );
  XNOR2_X1 DP_mult_218_U1638 ( .A(DP_coeff_pipe02[17]), .B(DP_mult_218_n1953), 
        .ZN(DP_mult_218_n777) );
  OAI22_X1 DP_mult_218_U1637 ( .A1(DP_mult_218_n1640), .A2(DP_mult_218_n1592), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1551), .ZN(DP_mult_218_n1952)
         );
  AOI221_X1 DP_mult_218_U1636 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1549), .C2(DP_mult_218_n1376), .A(DP_mult_218_n1952), 
        .ZN(DP_mult_218_n1951) );
  XNOR2_X1 DP_mult_218_U1635 ( .A(DP_coeff_pipe02[17]), .B(DP_mult_218_n1951), 
        .ZN(DP_mult_218_n778) );
  OAI22_X1 DP_mult_218_U1634 ( .A1(DP_mult_218_n1728), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1729), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1950)
         );
  AOI221_X1 DP_mult_218_U1633 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[21]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[20]), .A(DP_mult_218_n1950), 
        .ZN(DP_mult_218_n1949) );
  XNOR2_X1 DP_mult_218_U1632 ( .A(DP_coeff_pipe02[17]), .B(DP_mult_218_n1949), 
        .ZN(DP_mult_218_n779) );
  OAI22_X1 DP_mult_218_U1631 ( .A1(DP_mult_218_n1724), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1725), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1948)
         );
  AOI221_X1 DP_mult_218_U1630 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[20]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[19]), .A(DP_mult_218_n1948), 
        .ZN(DP_mult_218_n1947) );
  XNOR2_X1 DP_mult_218_U1629 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1947), 
        .ZN(DP_mult_218_n780) );
  OAI22_X1 DP_mult_218_U1628 ( .A1(DP_mult_218_n1720), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1721), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1946)
         );
  AOI221_X1 DP_mult_218_U1627 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[19]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[18]), .A(DP_mult_218_n1946), 
        .ZN(DP_mult_218_n1945) );
  XNOR2_X1 DP_mult_218_U1626 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1945), 
        .ZN(DP_mult_218_n781) );
  OAI22_X1 DP_mult_218_U1625 ( .A1(DP_mult_218_n1716), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1717), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1944)
         );
  AOI221_X1 DP_mult_218_U1624 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[18]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[17]), .A(DP_mult_218_n1944), 
        .ZN(DP_mult_218_n1943) );
  XNOR2_X1 DP_mult_218_U1623 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1943), 
        .ZN(DP_mult_218_n782) );
  OAI22_X1 DP_mult_218_U1622 ( .A1(DP_mult_218_n1712), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1713), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1942)
         );
  AOI221_X1 DP_mult_218_U1621 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[17]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[16]), .A(DP_mult_218_n1942), 
        .ZN(DP_mult_218_n1941) );
  XNOR2_X1 DP_mult_218_U1620 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1941), 
        .ZN(DP_mult_218_n783) );
  OAI22_X1 DP_mult_218_U1619 ( .A1(DP_mult_218_n1708), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1709), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1940)
         );
  AOI221_X1 DP_mult_218_U1618 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[16]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[15]), .A(DP_mult_218_n1940), 
        .ZN(DP_mult_218_n1939) );
  XNOR2_X1 DP_mult_218_U1617 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1939), 
        .ZN(DP_mult_218_n784) );
  OAI22_X1 DP_mult_218_U1616 ( .A1(DP_mult_218_n1704), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1705), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1938)
         );
  AOI221_X1 DP_mult_218_U1615 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[15]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[14]), .A(DP_mult_218_n1938), 
        .ZN(DP_mult_218_n1937) );
  XNOR2_X1 DP_mult_218_U1614 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1937), 
        .ZN(DP_mult_218_n785) );
  OAI22_X1 DP_mult_218_U1613 ( .A1(DP_mult_218_n1700), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1701), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1936)
         );
  AOI221_X1 DP_mult_218_U1612 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[14]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[13]), .A(DP_mult_218_n1936), 
        .ZN(DP_mult_218_n1935) );
  XNOR2_X1 DP_mult_218_U1611 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1935), 
        .ZN(DP_mult_218_n786) );
  OAI22_X1 DP_mult_218_U1610 ( .A1(DP_mult_218_n1696), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1697), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1934)
         );
  AOI221_X1 DP_mult_218_U1609 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[13]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[12]), .A(DP_mult_218_n1934), 
        .ZN(DP_mult_218_n1933) );
  XNOR2_X1 DP_mult_218_U1608 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1933), 
        .ZN(DP_mult_218_n787) );
  OAI22_X1 DP_mult_218_U1607 ( .A1(DP_mult_218_n1692), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1693), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1932)
         );
  AOI221_X1 DP_mult_218_U1606 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[12]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[11]), .A(DP_mult_218_n1932), 
        .ZN(DP_mult_218_n1931) );
  XNOR2_X1 DP_mult_218_U1605 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1931), 
        .ZN(DP_mult_218_n788) );
  OAI22_X1 DP_mult_218_U1604 ( .A1(DP_mult_218_n1688), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1689), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1930)
         );
  AOI221_X1 DP_mult_218_U1603 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[11]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[10]), .A(DP_mult_218_n1930), 
        .ZN(DP_mult_218_n1929) );
  XNOR2_X1 DP_mult_218_U1602 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1929), 
        .ZN(DP_mult_218_n789) );
  OAI22_X1 DP_mult_218_U1601 ( .A1(DP_mult_218_n1684), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1685), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1928)
         );
  AOI221_X1 DP_mult_218_U1600 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[10]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[9]), .A(DP_mult_218_n1928), .ZN(
        DP_mult_218_n1927) );
  XNOR2_X1 DP_mult_218_U1599 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1927), 
        .ZN(DP_mult_218_n790) );
  OAI22_X1 DP_mult_218_U1598 ( .A1(DP_mult_218_n1680), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1681), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1926)
         );
  AOI221_X1 DP_mult_218_U1597 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[9]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[8]), .A(DP_mult_218_n1926), .ZN(
        DP_mult_218_n1925) );
  XNOR2_X1 DP_mult_218_U1596 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1925), 
        .ZN(DP_mult_218_n791) );
  OAI22_X1 DP_mult_218_U1595 ( .A1(DP_mult_218_n1676), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1677), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1924)
         );
  AOI221_X1 DP_mult_218_U1594 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[8]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[7]), .A(DP_mult_218_n1924), .ZN(
        DP_mult_218_n1923) );
  XNOR2_X1 DP_mult_218_U1593 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1923), 
        .ZN(DP_mult_218_n792) );
  OAI22_X1 DP_mult_218_U1592 ( .A1(DP_mult_218_n1672), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1673), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1922)
         );
  AOI221_X1 DP_mult_218_U1591 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[7]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[6]), .A(DP_mult_218_n1922), .ZN(
        DP_mult_218_n1921) );
  XNOR2_X1 DP_mult_218_U1590 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1921), 
        .ZN(DP_mult_218_n793) );
  OAI22_X1 DP_mult_218_U1589 ( .A1(DP_mult_218_n1668), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1669), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1920)
         );
  AOI221_X1 DP_mult_218_U1588 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[6]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[5]), .A(DP_mult_218_n1920), .ZN(
        DP_mult_218_n1919) );
  XNOR2_X1 DP_mult_218_U1587 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1919), 
        .ZN(DP_mult_218_n794) );
  OAI22_X1 DP_mult_218_U1586 ( .A1(DP_mult_218_n1664), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1665), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1918)
         );
  AOI221_X1 DP_mult_218_U1585 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[5]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[4]), .A(DP_mult_218_n1918), .ZN(
        DP_mult_218_n1917) );
  XNOR2_X1 DP_mult_218_U1584 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1917), 
        .ZN(DP_mult_218_n795) );
  OAI22_X1 DP_mult_218_U1583 ( .A1(DP_mult_218_n1660), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1661), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1916)
         );
  AOI221_X1 DP_mult_218_U1582 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[4]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[3]), .A(DP_mult_218_n1916), .ZN(
        DP_mult_218_n1915) );
  XNOR2_X1 DP_mult_218_U1581 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1915), 
        .ZN(DP_mult_218_n796) );
  OAI22_X1 DP_mult_218_U1580 ( .A1(DP_mult_218_n1657), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1649), .B2(DP_mult_218_n1592), .ZN(DP_mult_218_n1914)
         );
  AOI221_X1 DP_mult_218_U1579 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[3]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[2]), .A(DP_mult_218_n1914), .ZN(
        DP_mult_218_n1913) );
  XNOR2_X1 DP_mult_218_U1578 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1913), 
        .ZN(DP_mult_218_n797) );
  OAI22_X1 DP_mult_218_U1577 ( .A1(DP_mult_218_n1653), .A2(DP_mult_218_n1588), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1591), .ZN(DP_mult_218_n1911)
         );
  AOI221_X1 DP_mult_218_U1576 ( .B1(DP_mult_218_n1589), .B2(DP_pipe02[2]), 
        .C1(DP_mult_218_n1590), .C2(DP_pipe02[1]), .A(DP_mult_218_n1911), .ZN(
        DP_mult_218_n1910) );
  XNOR2_X1 DP_mult_218_U1575 ( .A(DP_mult_218_n1606), .B(DP_mult_218_n1910), 
        .ZN(DP_mult_218_n798) );
  OAI222_X1 DP_mult_218_U1574 ( .A1(DP_mult_218_n1649), .A2(DP_mult_218_n1546), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1551), .C1(DP_mult_218_n1650), 
        .C2(DP_mult_218_n1588), .ZN(DP_mult_218_n1909) );
  XNOR2_X1 DP_mult_218_U1573 ( .A(DP_mult_218_n1909), .B(DP_mult_218_n1607), 
        .ZN(DP_mult_218_n799) );
  OAI22_X1 DP_mult_218_U1572 ( .A1(DP_mult_218_n1565), .A2(DP_mult_218_n1546), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1588), .ZN(DP_mult_218_n1908)
         );
  XNOR2_X1 DP_mult_218_U1571 ( .A(DP_mult_218_n1908), .B(DP_mult_218_n1607), 
        .ZN(DP_mult_218_n800) );
  XOR2_X1 DP_mult_218_U1570 ( .A(DP_coeff_pipe02[12]), .B(DP_mult_218_n1603), 
        .Z(DP_mult_218_n1907) );
  XNOR2_X1 DP_mult_218_U1569 ( .A(DP_coeff_pipe02[13]), .B(DP_mult_218_n1605), 
        .ZN(DP_mult_218_n1906) );
  XNOR2_X1 DP_mult_218_U1568 ( .A(DP_coeff_pipe02[12]), .B(DP_coeff_pipe02[13]), .ZN(DP_mult_218_n1905) );
  NAND3_X1 DP_mult_218_U1567 ( .A1(DP_mult_218_n1907), .A2(DP_mult_218_n1906), 
        .A3(DP_mult_218_n1905), .ZN(DP_mult_218_n1857) );
  INV_X1 DP_mult_218_U1566 ( .A(DP_mult_218_n1907), .ZN(DP_mult_218_n1904) );
  OAI21_X1 DP_mult_218_U1565 ( .B1(DP_mult_218_n1584), .B2(DP_mult_218_n1585), 
        .A(DP_mult_218_n1615), .ZN(DP_mult_218_n1903) );
  OAI221_X1 DP_mult_218_U1564 ( .B1(DP_mult_218_n1617), .B2(DP_mult_218_n1587), 
        .C1(DP_mult_218_n1620), .C2(DP_mult_218_n1583), .A(DP_mult_218_n1903), 
        .ZN(DP_mult_218_n1902) );
  XNOR2_X1 DP_mult_218_U1563 ( .A(DP_coeff_pipe02[14]), .B(DP_mult_218_n1902), 
        .ZN(DP_mult_218_n801) );
  OAI22_X1 DP_mult_218_U1562 ( .A1(DP_mult_218_n1633), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1634), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1901)
         );
  AOI221_X1 DP_mult_218_U1561 ( .B1(DP_mult_218_n1584), .B2(DP_mult_218_n1615), 
        .C1(DP_mult_218_n1585), .C2(DP_mult_218_n1615), .A(DP_mult_218_n1901), 
        .ZN(DP_mult_218_n1900) );
  XNOR2_X1 DP_mult_218_U1560 ( .A(DP_coeff_pipe02[14]), .B(DP_mult_218_n1900), 
        .ZN(DP_mult_218_n802) );
  OAI22_X1 DP_mult_218_U1559 ( .A1(DP_mult_218_n1617), .A2(DP_mult_218_n1545), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1899)
         );
  AOI221_X1 DP_mult_218_U1558 ( .B1(DP_mult_218_n1585), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1548), .C2(DP_mult_218_n1375), .A(DP_mult_218_n1899), 
        .ZN(DP_mult_218_n1898) );
  XNOR2_X1 DP_mult_218_U1557 ( .A(DP_coeff_pipe02[14]), .B(DP_mult_218_n1898), 
        .ZN(DP_mult_218_n803) );
  OAI22_X1 DP_mult_218_U1556 ( .A1(DP_mult_218_n1640), .A2(DP_mult_218_n1587), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1555), .ZN(DP_mult_218_n1897)
         );
  AOI221_X1 DP_mult_218_U1555 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1548), .C2(DP_mult_218_n1376), .A(DP_mult_218_n1897), 
        .ZN(DP_mult_218_n1896) );
  XNOR2_X1 DP_mult_218_U1554 ( .A(DP_coeff_pipe02[14]), .B(DP_mult_218_n1896), 
        .ZN(DP_mult_218_n804) );
  OAI22_X1 DP_mult_218_U1553 ( .A1(DP_mult_218_n1728), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1729), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1895)
         );
  AOI221_X1 DP_mult_218_U1552 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[21]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[20]), .A(DP_mult_218_n1895), 
        .ZN(DP_mult_218_n1894) );
  XNOR2_X1 DP_mult_218_U1551 ( .A(DP_coeff_pipe02[14]), .B(DP_mult_218_n1894), 
        .ZN(DP_mult_218_n805) );
  OAI22_X1 DP_mult_218_U1550 ( .A1(DP_mult_218_n1724), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1725), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1893)
         );
  AOI221_X1 DP_mult_218_U1549 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[20]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[19]), .A(DP_mult_218_n1893), 
        .ZN(DP_mult_218_n1892) );
  XNOR2_X1 DP_mult_218_U1548 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1892), 
        .ZN(DP_mult_218_n806) );
  OAI22_X1 DP_mult_218_U1547 ( .A1(DP_mult_218_n1720), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1721), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1891)
         );
  AOI221_X1 DP_mult_218_U1546 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[19]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[18]), .A(DP_mult_218_n1891), 
        .ZN(DP_mult_218_n1890) );
  XNOR2_X1 DP_mult_218_U1545 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1890), 
        .ZN(DP_mult_218_n807) );
  OAI22_X1 DP_mult_218_U1544 ( .A1(DP_mult_218_n1716), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1717), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1889)
         );
  AOI221_X1 DP_mult_218_U1543 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[18]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[17]), .A(DP_mult_218_n1889), 
        .ZN(DP_mult_218_n1888) );
  XNOR2_X1 DP_mult_218_U1542 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1888), 
        .ZN(DP_mult_218_n808) );
  OAI22_X1 DP_mult_218_U1541 ( .A1(DP_mult_218_n1712), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1713), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1887)
         );
  AOI221_X1 DP_mult_218_U1540 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[17]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[16]), .A(DP_mult_218_n1887), 
        .ZN(DP_mult_218_n1886) );
  XNOR2_X1 DP_mult_218_U1539 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1886), 
        .ZN(DP_mult_218_n809) );
  OAI22_X1 DP_mult_218_U1538 ( .A1(DP_mult_218_n1708), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1709), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1885)
         );
  AOI221_X1 DP_mult_218_U1537 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[16]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[15]), .A(DP_mult_218_n1885), 
        .ZN(DP_mult_218_n1884) );
  XNOR2_X1 DP_mult_218_U1536 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1884), 
        .ZN(DP_mult_218_n810) );
  OAI22_X1 DP_mult_218_U1535 ( .A1(DP_mult_218_n1704), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1705), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1883)
         );
  AOI221_X1 DP_mult_218_U1534 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[15]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[14]), .A(DP_mult_218_n1883), 
        .ZN(DP_mult_218_n1882) );
  XNOR2_X1 DP_mult_218_U1533 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1882), 
        .ZN(DP_mult_218_n811) );
  OAI22_X1 DP_mult_218_U1532 ( .A1(DP_mult_218_n1700), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1701), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1881)
         );
  AOI221_X1 DP_mult_218_U1531 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[14]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[13]), .A(DP_mult_218_n1881), 
        .ZN(DP_mult_218_n1880) );
  XNOR2_X1 DP_mult_218_U1530 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1880), 
        .ZN(DP_mult_218_n812) );
  OAI22_X1 DP_mult_218_U1529 ( .A1(DP_mult_218_n1696), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1697), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1879)
         );
  AOI221_X1 DP_mult_218_U1528 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[13]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[12]), .A(DP_mult_218_n1879), 
        .ZN(DP_mult_218_n1878) );
  XNOR2_X1 DP_mult_218_U1527 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1878), 
        .ZN(DP_mult_218_n813) );
  OAI22_X1 DP_mult_218_U1526 ( .A1(DP_mult_218_n1692), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1693), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1877)
         );
  AOI221_X1 DP_mult_218_U1525 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[12]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[11]), .A(DP_mult_218_n1877), 
        .ZN(DP_mult_218_n1876) );
  XNOR2_X1 DP_mult_218_U1524 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1876), 
        .ZN(DP_mult_218_n814) );
  OAI22_X1 DP_mult_218_U1523 ( .A1(DP_mult_218_n1688), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1689), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1875)
         );
  AOI221_X1 DP_mult_218_U1522 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[11]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[10]), .A(DP_mult_218_n1875), 
        .ZN(DP_mult_218_n1874) );
  XNOR2_X1 DP_mult_218_U1521 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1874), 
        .ZN(DP_mult_218_n815) );
  OAI22_X1 DP_mult_218_U1520 ( .A1(DP_mult_218_n1684), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1685), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1873)
         );
  AOI221_X1 DP_mult_218_U1519 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[10]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[9]), .A(DP_mult_218_n1873), .ZN(
        DP_mult_218_n1872) );
  XNOR2_X1 DP_mult_218_U1518 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1872), 
        .ZN(DP_mult_218_n816) );
  OAI22_X1 DP_mult_218_U1517 ( .A1(DP_mult_218_n1680), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1681), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1871)
         );
  AOI221_X1 DP_mult_218_U1516 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[9]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[8]), .A(DP_mult_218_n1871), .ZN(
        DP_mult_218_n1870) );
  XNOR2_X1 DP_mult_218_U1515 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1870), 
        .ZN(DP_mult_218_n817) );
  OAI22_X1 DP_mult_218_U1514 ( .A1(DP_mult_218_n1676), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1677), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1869)
         );
  AOI221_X1 DP_mult_218_U1513 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[8]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[7]), .A(DP_mult_218_n1869), .ZN(
        DP_mult_218_n1868) );
  XNOR2_X1 DP_mult_218_U1512 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1868), 
        .ZN(DP_mult_218_n818) );
  OAI22_X1 DP_mult_218_U1511 ( .A1(DP_mult_218_n1672), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1673), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1867)
         );
  AOI221_X1 DP_mult_218_U1510 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[7]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[6]), .A(DP_mult_218_n1867), .ZN(
        DP_mult_218_n1866) );
  XNOR2_X1 DP_mult_218_U1509 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1866), 
        .ZN(DP_mult_218_n819) );
  OAI22_X1 DP_mult_218_U1508 ( .A1(DP_mult_218_n1668), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1669), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1865)
         );
  AOI221_X1 DP_mult_218_U1507 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[6]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[5]), .A(DP_mult_218_n1865), .ZN(
        DP_mult_218_n1864) );
  XNOR2_X1 DP_mult_218_U1506 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1864), 
        .ZN(DP_mult_218_n820) );
  OAI22_X1 DP_mult_218_U1505 ( .A1(DP_mult_218_n1664), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1665), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1863)
         );
  AOI221_X1 DP_mult_218_U1504 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[5]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[4]), .A(DP_mult_218_n1863), .ZN(
        DP_mult_218_n1862) );
  XNOR2_X1 DP_mult_218_U1503 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1862), 
        .ZN(DP_mult_218_n821) );
  OAI22_X1 DP_mult_218_U1502 ( .A1(DP_mult_218_n1660), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1661), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1861)
         );
  AOI221_X1 DP_mult_218_U1501 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[4]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[3]), .A(DP_mult_218_n1861), .ZN(
        DP_mult_218_n1860) );
  XNOR2_X1 DP_mult_218_U1500 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1860), 
        .ZN(DP_mult_218_n822) );
  OAI22_X1 DP_mult_218_U1499 ( .A1(DP_mult_218_n1657), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1649), .B2(DP_mult_218_n1587), .ZN(DP_mult_218_n1859)
         );
  AOI221_X1 DP_mult_218_U1498 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[3]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[2]), .A(DP_mult_218_n1859), .ZN(
        DP_mult_218_n1858) );
  XNOR2_X1 DP_mult_218_U1497 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1858), 
        .ZN(DP_mult_218_n823) );
  OAI22_X1 DP_mult_218_U1496 ( .A1(DP_mult_218_n1653), .A2(DP_mult_218_n1583), 
        .B1(DP_mult_218_n1565), .B2(DP_mult_218_n1586), .ZN(DP_mult_218_n1856)
         );
  AOI221_X1 DP_mult_218_U1495 ( .B1(DP_mult_218_n1584), .B2(DP_pipe02[2]), 
        .C1(DP_mult_218_n1585), .C2(DP_pipe02[1]), .A(DP_mult_218_n1856), .ZN(
        DP_mult_218_n1855) );
  XNOR2_X1 DP_mult_218_U1494 ( .A(DP_mult_218_n1604), .B(DP_mult_218_n1855), 
        .ZN(DP_mult_218_n824) );
  OAI222_X1 DP_mult_218_U1493 ( .A1(DP_mult_218_n1649), .A2(DP_mult_218_n1545), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1555), .C1(DP_mult_218_n1650), 
        .C2(DP_mult_218_n1583), .ZN(DP_mult_218_n1854) );
  XNOR2_X1 DP_mult_218_U1492 ( .A(DP_mult_218_n1854), .B(DP_mult_218_n1605), 
        .ZN(DP_mult_218_n825) );
  OAI22_X1 DP_mult_218_U1491 ( .A1(DP_mult_218_n1565), .A2(DP_mult_218_n1545), 
        .B1(DP_mult_218_n1565), .B2(DP_mult_218_n1583), .ZN(DP_mult_218_n1853)
         );
  XNOR2_X1 DP_mult_218_U1490 ( .A(DP_mult_218_n1853), .B(DP_mult_218_n1605), 
        .ZN(DP_mult_218_n826) );
  XOR2_X1 DP_mult_218_U1489 ( .A(DP_coeff_pipe02[9]), .B(DP_mult_218_n1601), 
        .Z(DP_mult_218_n1852) );
  XNOR2_X1 DP_mult_218_U1488 ( .A(DP_coeff_pipe02[10]), .B(DP_mult_218_n1603), 
        .ZN(DP_mult_218_n1851) );
  XNOR2_X1 DP_mult_218_U1487 ( .A(DP_coeff_pipe02[10]), .B(DP_coeff_pipe02[9]), 
        .ZN(DP_mult_218_n1850) );
  NAND3_X1 DP_mult_218_U1486 ( .A1(DP_mult_218_n1852), .A2(DP_mult_218_n1851), 
        .A3(DP_mult_218_n1850), .ZN(DP_mult_218_n1802) );
  INV_X1 DP_mult_218_U1485 ( .A(DP_mult_218_n1852), .ZN(DP_mult_218_n1849) );
  OAI21_X1 DP_mult_218_U1484 ( .B1(DP_mult_218_n1579), .B2(DP_mult_218_n1580), 
        .A(DP_mult_218_n1615), .ZN(DP_mult_218_n1848) );
  OAI221_X1 DP_mult_218_U1483 ( .B1(DP_mult_218_n1618), .B2(DP_mult_218_n1582), 
        .C1(DP_mult_218_n1617), .C2(DP_mult_218_n1578), .A(DP_mult_218_n1848), 
        .ZN(DP_mult_218_n1847) );
  XNOR2_X1 DP_mult_218_U1482 ( .A(DP_coeff_pipe02[11]), .B(DP_mult_218_n1847), 
        .ZN(DP_mult_218_n827) );
  OAI22_X1 DP_mult_218_U1481 ( .A1(DP_mult_218_n1633), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1634), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1846)
         );
  AOI221_X1 DP_mult_218_U1480 ( .B1(DP_mult_218_n1579), .B2(DP_mult_218_n1615), 
        .C1(DP_mult_218_n1580), .C2(DP_mult_218_n1615), .A(DP_mult_218_n1846), 
        .ZN(DP_mult_218_n1845) );
  XNOR2_X1 DP_mult_218_U1479 ( .A(DP_coeff_pipe02[11]), .B(DP_mult_218_n1845), 
        .ZN(DP_mult_218_n828) );
  OAI22_X1 DP_mult_218_U1478 ( .A1(DP_mult_218_n1617), .A2(DP_mult_218_n1540), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1844)
         );
  AOI221_X1 DP_mult_218_U1477 ( .B1(DP_mult_218_n1580), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1541), .C2(DP_mult_218_n1375), .A(DP_mult_218_n1844), 
        .ZN(DP_mult_218_n1843) );
  XNOR2_X1 DP_mult_218_U1476 ( .A(DP_coeff_pipe02[11]), .B(DP_mult_218_n1843), 
        .ZN(DP_mult_218_n829) );
  OAI22_X1 DP_mult_218_U1475 ( .A1(DP_mult_218_n1640), .A2(DP_mult_218_n1582), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1533), .ZN(DP_mult_218_n1842)
         );
  AOI221_X1 DP_mult_218_U1474 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1541), .C2(DP_mult_218_n1376), .A(DP_mult_218_n1842), 
        .ZN(DP_mult_218_n1841) );
  XNOR2_X1 DP_mult_218_U1473 ( .A(DP_coeff_pipe02[11]), .B(DP_mult_218_n1841), 
        .ZN(DP_mult_218_n830) );
  OAI22_X1 DP_mult_218_U1472 ( .A1(DP_mult_218_n1728), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1729), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1840)
         );
  AOI221_X1 DP_mult_218_U1471 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[21]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[20]), .A(DP_mult_218_n1840), 
        .ZN(DP_mult_218_n1839) );
  XNOR2_X1 DP_mult_218_U1470 ( .A(DP_coeff_pipe02[11]), .B(DP_mult_218_n1839), 
        .ZN(DP_mult_218_n831) );
  OAI22_X1 DP_mult_218_U1469 ( .A1(DP_mult_218_n1724), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1725), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1838)
         );
  AOI221_X1 DP_mult_218_U1468 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[20]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[19]), .A(DP_mult_218_n1838), 
        .ZN(DP_mult_218_n1837) );
  XNOR2_X1 DP_mult_218_U1467 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1837), 
        .ZN(DP_mult_218_n832) );
  OAI22_X1 DP_mult_218_U1466 ( .A1(DP_mult_218_n1720), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1721), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1836)
         );
  AOI221_X1 DP_mult_218_U1465 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[19]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[18]), .A(DP_mult_218_n1836), 
        .ZN(DP_mult_218_n1835) );
  XNOR2_X1 DP_mult_218_U1464 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1835), 
        .ZN(DP_mult_218_n833) );
  OAI22_X1 DP_mult_218_U1463 ( .A1(DP_mult_218_n1716), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1717), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1834)
         );
  AOI221_X1 DP_mult_218_U1462 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[18]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[17]), .A(DP_mult_218_n1834), 
        .ZN(DP_mult_218_n1833) );
  XNOR2_X1 DP_mult_218_U1461 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1833), 
        .ZN(DP_mult_218_n834) );
  OAI22_X1 DP_mult_218_U1460 ( .A1(DP_mult_218_n1712), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1713), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1832)
         );
  AOI221_X1 DP_mult_218_U1459 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[17]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[16]), .A(DP_mult_218_n1832), 
        .ZN(DP_mult_218_n1831) );
  XNOR2_X1 DP_mult_218_U1458 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1831), 
        .ZN(DP_mult_218_n835) );
  OAI22_X1 DP_mult_218_U1457 ( .A1(DP_mult_218_n1708), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1709), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1830)
         );
  AOI221_X1 DP_mult_218_U1456 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[16]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[15]), .A(DP_mult_218_n1830), 
        .ZN(DP_mult_218_n1829) );
  XNOR2_X1 DP_mult_218_U1455 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1829), 
        .ZN(DP_mult_218_n836) );
  OAI22_X1 DP_mult_218_U1454 ( .A1(DP_mult_218_n1704), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1705), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1828)
         );
  AOI221_X1 DP_mult_218_U1453 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[15]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[14]), .A(DP_mult_218_n1828), 
        .ZN(DP_mult_218_n1827) );
  XNOR2_X1 DP_mult_218_U1452 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1827), 
        .ZN(DP_mult_218_n837) );
  OAI22_X1 DP_mult_218_U1451 ( .A1(DP_mult_218_n1700), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1701), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1826)
         );
  AOI221_X1 DP_mult_218_U1450 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[14]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[13]), .A(DP_mult_218_n1826), 
        .ZN(DP_mult_218_n1825) );
  XNOR2_X1 DP_mult_218_U1449 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1825), 
        .ZN(DP_mult_218_n838) );
  OAI22_X1 DP_mult_218_U1448 ( .A1(DP_mult_218_n1696), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1697), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1824)
         );
  AOI221_X1 DP_mult_218_U1447 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[13]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[12]), .A(DP_mult_218_n1824), 
        .ZN(DP_mult_218_n1823) );
  XNOR2_X1 DP_mult_218_U1446 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1823), 
        .ZN(DP_mult_218_n839) );
  OAI22_X1 DP_mult_218_U1445 ( .A1(DP_mult_218_n1692), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1693), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1822)
         );
  AOI221_X1 DP_mult_218_U1444 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[12]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[11]), .A(DP_mult_218_n1822), 
        .ZN(DP_mult_218_n1821) );
  XNOR2_X1 DP_mult_218_U1443 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1821), 
        .ZN(DP_mult_218_n840) );
  OAI22_X1 DP_mult_218_U1442 ( .A1(DP_mult_218_n1688), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1689), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1820)
         );
  AOI221_X1 DP_mult_218_U1441 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[11]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[10]), .A(DP_mult_218_n1820), 
        .ZN(DP_mult_218_n1819) );
  XNOR2_X1 DP_mult_218_U1440 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1819), 
        .ZN(DP_mult_218_n841) );
  OAI22_X1 DP_mult_218_U1439 ( .A1(DP_mult_218_n1684), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1685), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1818)
         );
  AOI221_X1 DP_mult_218_U1438 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[10]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[9]), .A(DP_mult_218_n1818), .ZN(
        DP_mult_218_n1817) );
  XNOR2_X1 DP_mult_218_U1437 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1817), 
        .ZN(DP_mult_218_n842) );
  OAI22_X1 DP_mult_218_U1436 ( .A1(DP_mult_218_n1680), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1681), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1816)
         );
  AOI221_X1 DP_mult_218_U1435 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[9]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[8]), .A(DP_mult_218_n1816), .ZN(
        DP_mult_218_n1815) );
  XNOR2_X1 DP_mult_218_U1434 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1815), 
        .ZN(DP_mult_218_n843) );
  OAI22_X1 DP_mult_218_U1433 ( .A1(DP_mult_218_n1676), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1677), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1814)
         );
  AOI221_X1 DP_mult_218_U1432 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[8]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[7]), .A(DP_mult_218_n1814), .ZN(
        DP_mult_218_n1813) );
  XNOR2_X1 DP_mult_218_U1431 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1813), 
        .ZN(DP_mult_218_n844) );
  OAI22_X1 DP_mult_218_U1430 ( .A1(DP_mult_218_n1672), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1673), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1812)
         );
  AOI221_X1 DP_mult_218_U1429 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[7]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[6]), .A(DP_mult_218_n1812), .ZN(
        DP_mult_218_n1811) );
  XNOR2_X1 DP_mult_218_U1428 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1811), 
        .ZN(DP_mult_218_n845) );
  OAI22_X1 DP_mult_218_U1427 ( .A1(DP_mult_218_n1668), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1669), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1810)
         );
  AOI221_X1 DP_mult_218_U1426 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[6]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[5]), .A(DP_mult_218_n1810), .ZN(
        DP_mult_218_n1809) );
  XNOR2_X1 DP_mult_218_U1425 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1809), 
        .ZN(DP_mult_218_n846) );
  OAI22_X1 DP_mult_218_U1424 ( .A1(DP_mult_218_n1664), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1665), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1808)
         );
  AOI221_X1 DP_mult_218_U1423 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[5]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[4]), .A(DP_mult_218_n1808), .ZN(
        DP_mult_218_n1807) );
  XNOR2_X1 DP_mult_218_U1422 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1807), 
        .ZN(DP_mult_218_n847) );
  OAI22_X1 DP_mult_218_U1421 ( .A1(DP_mult_218_n1660), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1661), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1806)
         );
  AOI221_X1 DP_mult_218_U1420 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[4]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[3]), .A(DP_mult_218_n1806), .ZN(
        DP_mult_218_n1805) );
  XNOR2_X1 DP_mult_218_U1419 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1805), 
        .ZN(DP_mult_218_n848) );
  OAI22_X1 DP_mult_218_U1418 ( .A1(DP_mult_218_n1657), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1649), .B2(DP_mult_218_n1582), .ZN(DP_mult_218_n1804)
         );
  AOI221_X1 DP_mult_218_U1417 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[3]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[2]), .A(DP_mult_218_n1804), .ZN(
        DP_mult_218_n1803) );
  XNOR2_X1 DP_mult_218_U1416 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1803), 
        .ZN(DP_mult_218_n849) );
  OAI22_X1 DP_mult_218_U1415 ( .A1(DP_mult_218_n1653), .A2(DP_mult_218_n1578), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1581), .ZN(DP_mult_218_n1801)
         );
  AOI221_X1 DP_mult_218_U1414 ( .B1(DP_mult_218_n1579), .B2(DP_pipe02[2]), 
        .C1(DP_mult_218_n1580), .C2(DP_pipe02[1]), .A(DP_mult_218_n1801), .ZN(
        DP_mult_218_n1800) );
  XNOR2_X1 DP_mult_218_U1413 ( .A(DP_mult_218_n1602), .B(DP_mult_218_n1800), 
        .ZN(DP_mult_218_n850) );
  OAI222_X1 DP_mult_218_U1412 ( .A1(DP_mult_218_n1649), .A2(DP_mult_218_n1540), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1533), .C1(DP_mult_218_n1650), 
        .C2(DP_mult_218_n1578), .ZN(DP_mult_218_n1799) );
  XNOR2_X1 DP_mult_218_U1411 ( .A(DP_mult_218_n1799), .B(DP_mult_218_n1603), 
        .ZN(DP_mult_218_n851) );
  OAI22_X1 DP_mult_218_U1410 ( .A1(DP_mult_218_n1565), .A2(DP_mult_218_n1540), 
        .B1(DP_mult_218_n1565), .B2(DP_mult_218_n1578), .ZN(DP_mult_218_n1798)
         );
  XNOR2_X1 DP_mult_218_U1409 ( .A(DP_mult_218_n1798), .B(DP_mult_218_n1603), 
        .ZN(DP_mult_218_n852) );
  XOR2_X1 DP_mult_218_U1408 ( .A(DP_coeff_pipe02[6]), .B(DP_mult_218_n1599), 
        .Z(DP_mult_218_n1797) );
  XNOR2_X1 DP_mult_218_U1407 ( .A(DP_coeff_pipe02[7]), .B(DP_mult_218_n1601), 
        .ZN(DP_mult_218_n1796) );
  XNOR2_X1 DP_mult_218_U1406 ( .A(DP_coeff_pipe02[6]), .B(DP_coeff_pipe02[7]), 
        .ZN(DP_mult_218_n1795) );
  NAND3_X1 DP_mult_218_U1405 ( .A1(DP_mult_218_n1797), .A2(DP_mult_218_n1796), 
        .A3(DP_mult_218_n1795), .ZN(DP_mult_218_n1747) );
  INV_X1 DP_mult_218_U1404 ( .A(DP_mult_218_n1797), .ZN(DP_mult_218_n1794) );
  OAI21_X1 DP_mult_218_U1403 ( .B1(DP_mult_218_n1574), .B2(DP_mult_218_n1575), 
        .A(DP_mult_218_n1615), .ZN(DP_mult_218_n1793) );
  OAI221_X1 DP_mult_218_U1402 ( .B1(DP_mult_218_n1618), .B2(DP_mult_218_n1577), 
        .C1(DP_mult_218_n1617), .C2(DP_mult_218_n1573), .A(DP_mult_218_n1793), 
        .ZN(DP_mult_218_n1792) );
  XNOR2_X1 DP_mult_218_U1401 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1792), 
        .ZN(DP_mult_218_n853) );
  OAI22_X1 DP_mult_218_U1400 ( .A1(DP_mult_218_n1633), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1634), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1791)
         );
  AOI221_X1 DP_mult_218_U1399 ( .B1(DP_mult_218_n1574), .B2(DP_mult_218_n1614), 
        .C1(DP_mult_218_n1575), .C2(DP_mult_218_n1615), .A(DP_mult_218_n1791), 
        .ZN(DP_mult_218_n1790) );
  XNOR2_X1 DP_mult_218_U1398 ( .A(DP_coeff_pipe02[8]), .B(DP_mult_218_n1790), 
        .ZN(DP_mult_218_n854) );
  OAI22_X1 DP_mult_218_U1397 ( .A1(DP_mult_218_n1617), .A2(DP_mult_218_n1534), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1789)
         );
  AOI221_X1 DP_mult_218_U1396 ( .B1(DP_mult_218_n1575), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1535), .C2(DP_mult_218_n1375), .A(DP_mult_218_n1789), 
        .ZN(DP_mult_218_n1788) );
  XNOR2_X1 DP_mult_218_U1395 ( .A(DP_coeff_pipe02[8]), .B(DP_mult_218_n1788), 
        .ZN(DP_mult_218_n855) );
  OAI22_X1 DP_mult_218_U1394 ( .A1(DP_mult_218_n1640), .A2(DP_mult_218_n1577), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1536), .ZN(DP_mult_218_n1787)
         );
  AOI221_X1 DP_mult_218_U1393 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1535), .C2(DP_mult_218_n1376), .A(DP_mult_218_n1787), 
        .ZN(DP_mult_218_n1786) );
  XNOR2_X1 DP_mult_218_U1392 ( .A(DP_coeff_pipe02[8]), .B(DP_mult_218_n1786), 
        .ZN(DP_mult_218_n856) );
  OAI22_X1 DP_mult_218_U1391 ( .A1(DP_mult_218_n1728), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1729), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1785)
         );
  AOI221_X1 DP_mult_218_U1390 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[21]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[20]), .A(DP_mult_218_n1785), 
        .ZN(DP_mult_218_n1784) );
  XNOR2_X1 DP_mult_218_U1389 ( .A(DP_coeff_pipe02[8]), .B(DP_mult_218_n1784), 
        .ZN(DP_mult_218_n857) );
  OAI22_X1 DP_mult_218_U1388 ( .A1(DP_mult_218_n1724), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1725), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1783)
         );
  AOI221_X1 DP_mult_218_U1387 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[20]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[19]), .A(DP_mult_218_n1783), 
        .ZN(DP_mult_218_n1782) );
  XNOR2_X1 DP_mult_218_U1386 ( .A(DP_coeff_pipe02[8]), .B(DP_mult_218_n1782), 
        .ZN(DP_mult_218_n858) );
  OAI22_X1 DP_mult_218_U1385 ( .A1(DP_mult_218_n1720), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1721), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1781)
         );
  AOI221_X1 DP_mult_218_U1384 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[19]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[18]), .A(DP_mult_218_n1781), 
        .ZN(DP_mult_218_n1780) );
  XNOR2_X1 DP_mult_218_U1383 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1780), 
        .ZN(DP_mult_218_n859) );
  OAI22_X1 DP_mult_218_U1382 ( .A1(DP_mult_218_n1716), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1717), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1779)
         );
  AOI221_X1 DP_mult_218_U1381 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[18]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[17]), .A(DP_mult_218_n1779), 
        .ZN(DP_mult_218_n1778) );
  XNOR2_X1 DP_mult_218_U1380 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1778), 
        .ZN(DP_mult_218_n860) );
  OAI22_X1 DP_mult_218_U1379 ( .A1(DP_mult_218_n1712), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1713), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1777)
         );
  AOI221_X1 DP_mult_218_U1378 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[17]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[16]), .A(DP_mult_218_n1777), 
        .ZN(DP_mult_218_n1776) );
  XNOR2_X1 DP_mult_218_U1377 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1776), 
        .ZN(DP_mult_218_n861) );
  OAI22_X1 DP_mult_218_U1376 ( .A1(DP_mult_218_n1708), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1709), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1775)
         );
  AOI221_X1 DP_mult_218_U1375 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[16]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[15]), .A(DP_mult_218_n1775), 
        .ZN(DP_mult_218_n1774) );
  XNOR2_X1 DP_mult_218_U1374 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1774), 
        .ZN(DP_mult_218_n862) );
  OAI22_X1 DP_mult_218_U1373 ( .A1(DP_mult_218_n1704), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1705), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1773)
         );
  AOI221_X1 DP_mult_218_U1372 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[15]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[14]), .A(DP_mult_218_n1773), 
        .ZN(DP_mult_218_n1772) );
  XNOR2_X1 DP_mult_218_U1371 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1772), 
        .ZN(DP_mult_218_n863) );
  OAI22_X1 DP_mult_218_U1370 ( .A1(DP_mult_218_n1700), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1701), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1771)
         );
  AOI221_X1 DP_mult_218_U1369 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[14]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[13]), .A(DP_mult_218_n1771), 
        .ZN(DP_mult_218_n1770) );
  XNOR2_X1 DP_mult_218_U1368 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1770), 
        .ZN(DP_mult_218_n864) );
  OAI22_X1 DP_mult_218_U1367 ( .A1(DP_mult_218_n1696), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1697), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1769)
         );
  AOI221_X1 DP_mult_218_U1366 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[13]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[12]), .A(DP_mult_218_n1769), 
        .ZN(DP_mult_218_n1768) );
  XNOR2_X1 DP_mult_218_U1365 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1768), 
        .ZN(DP_mult_218_n865) );
  OAI22_X1 DP_mult_218_U1364 ( .A1(DP_mult_218_n1692), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1693), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1767)
         );
  AOI221_X1 DP_mult_218_U1363 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[12]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[11]), .A(DP_mult_218_n1767), 
        .ZN(DP_mult_218_n1766) );
  XNOR2_X1 DP_mult_218_U1362 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1766), 
        .ZN(DP_mult_218_n866) );
  OAI22_X1 DP_mult_218_U1361 ( .A1(DP_mult_218_n1688), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1689), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1765)
         );
  AOI221_X1 DP_mult_218_U1360 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[11]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[10]), .A(DP_mult_218_n1765), 
        .ZN(DP_mult_218_n1764) );
  XNOR2_X1 DP_mult_218_U1359 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1764), 
        .ZN(DP_mult_218_n867) );
  OAI22_X1 DP_mult_218_U1358 ( .A1(DP_mult_218_n1684), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1685), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1763)
         );
  AOI221_X1 DP_mult_218_U1357 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[10]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[9]), .A(DP_mult_218_n1763), .ZN(
        DP_mult_218_n1762) );
  XNOR2_X1 DP_mult_218_U1356 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1762), 
        .ZN(DP_mult_218_n868) );
  OAI22_X1 DP_mult_218_U1355 ( .A1(DP_mult_218_n1680), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1681), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1761)
         );
  AOI221_X1 DP_mult_218_U1354 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[9]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[8]), .A(DP_mult_218_n1761), .ZN(
        DP_mult_218_n1760) );
  XNOR2_X1 DP_mult_218_U1353 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1760), 
        .ZN(DP_mult_218_n869) );
  OAI22_X1 DP_mult_218_U1352 ( .A1(DP_mult_218_n1676), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1677), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1759)
         );
  AOI221_X1 DP_mult_218_U1351 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[8]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[7]), .A(DP_mult_218_n1759), .ZN(
        DP_mult_218_n1758) );
  XNOR2_X1 DP_mult_218_U1350 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1758), 
        .ZN(DP_mult_218_n870) );
  OAI22_X1 DP_mult_218_U1349 ( .A1(DP_mult_218_n1672), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1673), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1757)
         );
  AOI221_X1 DP_mult_218_U1348 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[7]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[6]), .A(DP_mult_218_n1757), .ZN(
        DP_mult_218_n1756) );
  XNOR2_X1 DP_mult_218_U1347 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1756), 
        .ZN(DP_mult_218_n871) );
  OAI22_X1 DP_mult_218_U1346 ( .A1(DP_mult_218_n1668), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1669), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1755)
         );
  AOI221_X1 DP_mult_218_U1345 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[6]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[5]), .A(DP_mult_218_n1755), .ZN(
        DP_mult_218_n1754) );
  XNOR2_X1 DP_mult_218_U1344 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1754), 
        .ZN(DP_mult_218_n872) );
  OAI22_X1 DP_mult_218_U1343 ( .A1(DP_mult_218_n1664), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1665), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1753)
         );
  AOI221_X1 DP_mult_218_U1342 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[5]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[4]), .A(DP_mult_218_n1753), .ZN(
        DP_mult_218_n1752) );
  XNOR2_X1 DP_mult_218_U1341 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1752), 
        .ZN(DP_mult_218_n873) );
  OAI22_X1 DP_mult_218_U1340 ( .A1(DP_mult_218_n1660), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1661), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1751)
         );
  AOI221_X1 DP_mult_218_U1339 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[4]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[3]), .A(DP_mult_218_n1751), .ZN(
        DP_mult_218_n1750) );
  XNOR2_X1 DP_mult_218_U1338 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1750), 
        .ZN(DP_mult_218_n874) );
  OAI22_X1 DP_mult_218_U1337 ( .A1(DP_mult_218_n1657), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1649), .B2(DP_mult_218_n1577), .ZN(DP_mult_218_n1749)
         );
  AOI221_X1 DP_mult_218_U1336 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[3]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[2]), .A(DP_mult_218_n1749), .ZN(
        DP_mult_218_n1748) );
  XNOR2_X1 DP_mult_218_U1335 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1748), 
        .ZN(DP_mult_218_n875) );
  OAI22_X1 DP_mult_218_U1334 ( .A1(DP_mult_218_n1653), .A2(DP_mult_218_n1573), 
        .B1(DP_mult_218_n1565), .B2(DP_mult_218_n1576), .ZN(DP_mult_218_n1746)
         );
  AOI221_X1 DP_mult_218_U1333 ( .B1(DP_mult_218_n1574), .B2(DP_pipe02[2]), 
        .C1(DP_mult_218_n1575), .C2(DP_pipe02[1]), .A(DP_mult_218_n1746), .ZN(
        DP_mult_218_n1745) );
  XNOR2_X1 DP_mult_218_U1332 ( .A(DP_mult_218_n1600), .B(DP_mult_218_n1745), 
        .ZN(DP_mult_218_n876) );
  OAI222_X1 DP_mult_218_U1331 ( .A1(DP_mult_218_n1649), .A2(DP_mult_218_n1534), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1536), .C1(DP_mult_218_n1650), 
        .C2(DP_mult_218_n1573), .ZN(DP_mult_218_n1744) );
  XNOR2_X1 DP_mult_218_U1330 ( .A(DP_mult_218_n1744), .B(DP_mult_218_n1601), 
        .ZN(DP_mult_218_n877) );
  OAI22_X1 DP_mult_218_U1329 ( .A1(DP_mult_218_n1565), .A2(DP_mult_218_n1534), 
        .B1(DP_mult_218_n1565), .B2(DP_mult_218_n1573), .ZN(DP_mult_218_n1743)
         );
  XNOR2_X1 DP_mult_218_U1328 ( .A(DP_mult_218_n1743), .B(DP_mult_218_n1601), 
        .ZN(DP_mult_218_n878) );
  XOR2_X1 DP_mult_218_U1327 ( .A(DP_coeff_pipe02[3]), .B(DP_mult_218_n1742), 
        .Z(DP_mult_218_n1741) );
  XNOR2_X1 DP_mult_218_U1326 ( .A(DP_coeff_pipe02[4]), .B(DP_mult_218_n1599), 
        .ZN(DP_mult_218_n1740) );
  XNOR2_X1 DP_mult_218_U1325 ( .A(DP_coeff_pipe02[3]), .B(DP_coeff_pipe02[4]), 
        .ZN(DP_mult_218_n1739) );
  NAND3_X1 DP_mult_218_U1324 ( .A1(DP_mult_218_n1741), .A2(DP_mult_218_n1740), 
        .A3(DP_mult_218_n1739), .ZN(DP_mult_218_n1654) );
  INV_X1 DP_mult_218_U1323 ( .A(DP_mult_218_n1741), .ZN(DP_mult_218_n1738) );
  OAI21_X1 DP_mult_218_U1322 ( .B1(DP_mult_218_n1569), .B2(DP_mult_218_n1570), 
        .A(DP_mult_218_n1615), .ZN(DP_mult_218_n1737) );
  OAI221_X1 DP_mult_218_U1321 ( .B1(DP_mult_218_n1618), .B2(DP_mult_218_n1572), 
        .C1(DP_mult_218_n1618), .C2(DP_mult_218_n1568), .A(DP_mult_218_n1737), 
        .ZN(DP_mult_218_n1736) );
  XNOR2_X1 DP_mult_218_U1320 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1736), 
        .ZN(DP_mult_218_n879) );
  OAI22_X1 DP_mult_218_U1319 ( .A1(DP_mult_218_n1633), .A2(DP_mult_218_n1568), 
        .B1(DP_mult_218_n1634), .B2(DP_mult_218_n1572), .ZN(DP_mult_218_n1735)
         );
  AOI221_X1 DP_mult_218_U1318 ( .B1(DP_mult_218_n1569), .B2(DP_mult_218_n1614), 
        .C1(DP_mult_218_n1570), .C2(DP_mult_218_n1615), .A(DP_mult_218_n1735), 
        .ZN(DP_mult_218_n1734) );
  XNOR2_X1 DP_mult_218_U1317 ( .A(DP_coeff_pipe02[5]), .B(DP_mult_218_n1734), 
        .ZN(DP_mult_218_n880) );
  OAI22_X1 DP_mult_218_U1316 ( .A1(DP_mult_218_n1616), .A2(DP_mult_218_n1538), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1572), .ZN(DP_mult_218_n1733)
         );
  AOI221_X1 DP_mult_218_U1315 ( .B1(DP_mult_218_n1570), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1537), .C2(DP_mult_218_n1375), .A(DP_mult_218_n1733), 
        .ZN(DP_mult_218_n1732) );
  XNOR2_X1 DP_mult_218_U1314 ( .A(DP_coeff_pipe02[5]), .B(DP_mult_218_n1732), 
        .ZN(DP_mult_218_n881) );
  OAI22_X1 DP_mult_218_U1313 ( .A1(DP_mult_218_n1640), .A2(DP_mult_218_n1572), 
        .B1(DP_mult_218_n1643), .B2(DP_mult_218_n1539), .ZN(DP_mult_218_n1731)
         );
  AOI221_X1 DP_mult_218_U1312 ( .B1(DP_mult_218_n1569), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1537), .C2(DP_mult_218_n1376), .A(DP_mult_218_n1731), 
        .ZN(DP_mult_218_n1730) );
  XNOR2_X1 DP_mult_218_U1311 ( .A(DP_coeff_pipe02[5]), .B(DP_mult_218_n1730), 
        .ZN(DP_mult_218_n882) );
  OAI22_X1 DP_mult_218_U1310 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1728), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1729), .ZN(DP_mult_218_n1727)
         );
  AOI221_X1 DP_mult_218_U1309 ( .B1(DP_mult_218_n1569), .B2(DP_pipe02[21]), 
        .C1(DP_mult_218_n1570), .C2(DP_pipe02[20]), .A(DP_mult_218_n1727), 
        .ZN(DP_mult_218_n1726) );
  XNOR2_X1 DP_mult_218_U1308 ( .A(DP_coeff_pipe02[5]), .B(DP_mult_218_n1726), 
        .ZN(DP_mult_218_n883) );
  OAI22_X1 DP_mult_218_U1307 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1724), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1725), .ZN(DP_mult_218_n1723)
         );
  AOI221_X1 DP_mult_218_U1306 ( .B1(DP_mult_218_n1569), .B2(DP_pipe02[20]), 
        .C1(DP_pipe02[19]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1723), 
        .ZN(DP_mult_218_n1722) );
  XNOR2_X1 DP_mult_218_U1305 ( .A(DP_coeff_pipe02[5]), .B(DP_mult_218_n1722), 
        .ZN(DP_mult_218_n884) );
  OAI22_X1 DP_mult_218_U1304 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1720), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1721), .ZN(DP_mult_218_n1719)
         );
  AOI221_X1 DP_mult_218_U1303 ( .B1(DP_pipe02[19]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[18]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1719), 
        .ZN(DP_mult_218_n1718) );
  XNOR2_X1 DP_mult_218_U1302 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1718), 
        .ZN(DP_mult_218_n885) );
  OAI22_X1 DP_mult_218_U1301 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1716), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1717), .ZN(DP_mult_218_n1715)
         );
  AOI221_X1 DP_mult_218_U1300 ( .B1(DP_pipe02[18]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[17]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1715), 
        .ZN(DP_mult_218_n1714) );
  XNOR2_X1 DP_mult_218_U1299 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1714), 
        .ZN(DP_mult_218_n886) );
  OAI22_X1 DP_mult_218_U1298 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1712), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1713), .ZN(DP_mult_218_n1711)
         );
  AOI221_X1 DP_mult_218_U1297 ( .B1(DP_pipe02[17]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[16]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1711), 
        .ZN(DP_mult_218_n1710) );
  XNOR2_X1 DP_mult_218_U1296 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1710), 
        .ZN(DP_mult_218_n887) );
  OAI22_X1 DP_mult_218_U1295 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1708), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1709), .ZN(DP_mult_218_n1707)
         );
  AOI221_X1 DP_mult_218_U1294 ( .B1(DP_pipe02[16]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[15]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1707), 
        .ZN(DP_mult_218_n1706) );
  XNOR2_X1 DP_mult_218_U1293 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1706), 
        .ZN(DP_mult_218_n888) );
  OAI22_X1 DP_mult_218_U1292 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1704), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1705), .ZN(DP_mult_218_n1703)
         );
  AOI221_X1 DP_mult_218_U1291 ( .B1(DP_pipe02[15]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[14]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1703), 
        .ZN(DP_mult_218_n1702) );
  XNOR2_X1 DP_mult_218_U1290 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1702), 
        .ZN(DP_mult_218_n889) );
  OAI22_X1 DP_mult_218_U1289 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1700), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1701), .ZN(DP_mult_218_n1699)
         );
  AOI221_X1 DP_mult_218_U1288 ( .B1(DP_pipe02[14]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[13]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1699), 
        .ZN(DP_mult_218_n1698) );
  XNOR2_X1 DP_mult_218_U1287 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1698), 
        .ZN(DP_mult_218_n890) );
  OAI22_X1 DP_mult_218_U1286 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1696), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1697), .ZN(DP_mult_218_n1695)
         );
  AOI221_X1 DP_mult_218_U1285 ( .B1(DP_pipe02[13]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[12]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1695), 
        .ZN(DP_mult_218_n1694) );
  XNOR2_X1 DP_mult_218_U1284 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1694), 
        .ZN(DP_mult_218_n891) );
  OAI22_X1 DP_mult_218_U1283 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1692), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1693), .ZN(DP_mult_218_n1691)
         );
  AOI221_X1 DP_mult_218_U1282 ( .B1(DP_pipe02[12]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[11]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1691), 
        .ZN(DP_mult_218_n1690) );
  XNOR2_X1 DP_mult_218_U1281 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1690), 
        .ZN(DP_mult_218_n892) );
  OAI22_X1 DP_mult_218_U1280 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1688), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1689), .ZN(DP_mult_218_n1687)
         );
  AOI221_X1 DP_mult_218_U1279 ( .B1(DP_pipe02[11]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[10]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1687), 
        .ZN(DP_mult_218_n1686) );
  XNOR2_X1 DP_mult_218_U1278 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1686), 
        .ZN(DP_mult_218_n893) );
  OAI22_X1 DP_mult_218_U1277 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1684), 
        .B1(DP_mult_218_n1572), .B2(DP_mult_218_n1685), .ZN(DP_mult_218_n1683)
         );
  AOI221_X1 DP_mult_218_U1276 ( .B1(DP_pipe02[10]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[9]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1683), .ZN(
        DP_mult_218_n1682) );
  XNOR2_X1 DP_mult_218_U1275 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1682), 
        .ZN(DP_mult_218_n894) );
  OAI22_X1 DP_mult_218_U1274 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1680), 
        .B1(DP_mult_218_n1572), .B2(DP_mult_218_n1681), .ZN(DP_mult_218_n1679)
         );
  AOI221_X1 DP_mult_218_U1273 ( .B1(DP_pipe02[9]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[8]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1679), .ZN(
        DP_mult_218_n1678) );
  XNOR2_X1 DP_mult_218_U1272 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1678), 
        .ZN(DP_mult_218_n895) );
  OAI22_X1 DP_mult_218_U1271 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1676), 
        .B1(DP_mult_218_n1571), .B2(DP_mult_218_n1677), .ZN(DP_mult_218_n1675)
         );
  AOI221_X1 DP_mult_218_U1270 ( .B1(DP_pipe02[8]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[7]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1675), .ZN(
        DP_mult_218_n1674) );
  XNOR2_X1 DP_mult_218_U1269 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1674), 
        .ZN(DP_mult_218_n896) );
  OAI22_X1 DP_mult_218_U1268 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1672), 
        .B1(DP_mult_218_n1572), .B2(DP_mult_218_n1673), .ZN(DP_mult_218_n1671)
         );
  AOI221_X1 DP_mult_218_U1267 ( .B1(DP_pipe02[7]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[6]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1671), .ZN(
        DP_mult_218_n1670) );
  XNOR2_X1 DP_mult_218_U1266 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1670), 
        .ZN(DP_mult_218_n897) );
  OAI22_X1 DP_mult_218_U1265 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1668), 
        .B1(DP_mult_218_n1572), .B2(DP_mult_218_n1669), .ZN(DP_mult_218_n1667)
         );
  AOI221_X1 DP_mult_218_U1264 ( .B1(DP_pipe02[6]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[5]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1667), .ZN(
        DP_mult_218_n1666) );
  XNOR2_X1 DP_mult_218_U1263 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1666), 
        .ZN(DP_mult_218_n898) );
  OAI22_X1 DP_mult_218_U1262 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1664), 
        .B1(DP_mult_218_n1572), .B2(DP_mult_218_n1665), .ZN(DP_mult_218_n1663)
         );
  AOI221_X1 DP_mult_218_U1261 ( .B1(DP_pipe02[5]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[4]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1663), .ZN(
        DP_mult_218_n1662) );
  XNOR2_X1 DP_mult_218_U1260 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1662), 
        .ZN(DP_mult_218_n899) );
  OAI22_X1 DP_mult_218_U1259 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1660), 
        .B1(DP_mult_218_n1661), .B2(DP_mult_218_n1572), .ZN(DP_mult_218_n1659)
         );
  AOI221_X1 DP_mult_218_U1258 ( .B1(DP_pipe02[4]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[3]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1659), .ZN(
        DP_mult_218_n1658) );
  XNOR2_X1 DP_mult_218_U1257 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1658), 
        .ZN(DP_mult_218_n900) );
  OAI22_X1 DP_mult_218_U1256 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1657), 
        .B1(DP_mult_218_n1649), .B2(DP_mult_218_n1572), .ZN(DP_mult_218_n1656)
         );
  AOI221_X1 DP_mult_218_U1255 ( .B1(DP_pipe02[3]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[2]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1656), .ZN(
        DP_mult_218_n1655) );
  XNOR2_X1 DP_mult_218_U1254 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1655), 
        .ZN(DP_mult_218_n901) );
  OAI22_X1 DP_mult_218_U1253 ( .A1(DP_mult_218_n1568), .A2(DP_mult_218_n1653), 
        .B1(DP_mult_218_n1565), .B2(DP_mult_218_n1572), .ZN(DP_mult_218_n1652)
         );
  AOI221_X1 DP_mult_218_U1252 ( .B1(DP_pipe02[2]), .B2(DP_mult_218_n1569), 
        .C1(DP_pipe02[1]), .C2(DP_mult_218_n1570), .A(DP_mult_218_n1652), .ZN(
        DP_mult_218_n1651) );
  XNOR2_X1 DP_mult_218_U1251 ( .A(DP_mult_218_n1598), .B(DP_mult_218_n1651), 
        .ZN(DP_mult_218_n902) );
  OAI222_X1 DP_mult_218_U1250 ( .A1(DP_mult_218_n1538), .A2(DP_mult_218_n1649), 
        .B1(DP_mult_218_n1566), .B2(DP_mult_218_n1539), .C1(DP_mult_218_n1568), 
        .C2(DP_mult_218_n1650), .ZN(DP_mult_218_n1648) );
  XNOR2_X1 DP_mult_218_U1249 ( .A(DP_mult_218_n1648), .B(DP_mult_218_n1599), 
        .ZN(DP_mult_218_n903) );
  OAI22_X1 DP_mult_218_U1248 ( .A1(DP_mult_218_n1565), .A2(DP_mult_218_n1538), 
        .B1(DP_mult_218_n1568), .B2(DP_mult_218_n1567), .ZN(DP_mult_218_n1646)
         );
  XNOR2_X1 DP_mult_218_U1247 ( .A(DP_mult_218_n1646), .B(DP_mult_218_n1599), 
        .ZN(DP_mult_218_n904) );
  OAI22_X1 DP_mult_218_U1246 ( .A1(DP_mult_218_n1633), .A2(DP_mult_218_n1564), 
        .B1(DP_mult_218_n1634), .B2(DP_mult_218_n1639), .ZN(DP_mult_218_n1645)
         );
  AOI221_X1 DP_mult_218_U1245 ( .B1(DP_mult_218_n1561), .B2(DP_mult_218_n1614), 
        .C1(DP_mult_218_n1563), .C2(DP_mult_218_n1615), .A(DP_mult_218_n1645), 
        .ZN(DP_mult_218_n1644) );
  XNOR2_X1 DP_mult_218_U1244 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n1644), 
        .ZN(DP_mult_218_n906) );
  OAI22_X1 DP_mult_218_U1243 ( .A1(DP_mult_218_n1643), .A2(DP_mult_218_n1639), 
        .B1(DP_mult_218_n1617), .B2(DP_mult_218_n1542), .ZN(DP_mult_218_n1642)
         );
  AOI221_X1 DP_mult_218_U1242 ( .B1(DP_mult_218_n1563), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1554), .C2(DP_mult_218_n1375), .A(DP_mult_218_n1642), 
        .ZN(DP_mult_218_n1641) );
  XNOR2_X1 DP_mult_218_U1241 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n1641), 
        .ZN(DP_mult_218_n907) );
  INV_X1 DP_mult_218_U1240 ( .A(DP_mult_218_n1376), .ZN(DP_mult_218_n1638) );
  OAI22_X1 DP_mult_218_U1239 ( .A1(DP_mult_218_n1564), .A2(DP_mult_218_n1638), 
        .B1(DP_mult_218_n1639), .B2(DP_mult_218_n1640), .ZN(DP_mult_218_n1637)
         );
  AOI221_X1 DP_mult_218_U1238 ( .B1(DP_mult_218_n1561), .B2(DP_pipe02[22]), 
        .C1(DP_mult_218_n1563), .C2(DP_pipe02[21]), .A(DP_mult_218_n1637), 
        .ZN(DP_mult_218_n1635) );
  XNOR2_X1 DP_mult_218_U1237 ( .A(DP_coeff_pipe02[2]), .B(DP_mult_218_n1635), 
        .ZN(DP_mult_218_n908) );
  OAI22_X1 DP_mult_218_U1236 ( .A1(DP_mult_218_n1558), .A2(DP_mult_218_n1633), 
        .B1(DP_mult_218_n1557), .B2(DP_mult_218_n1634), .ZN(DP_mult_218_n1632)
         );
  AOI221_X1 DP_mult_218_U1235 ( .B1(DP_mult_218_n1613), .B2(DP_mult_218_n1559), 
        .C1(DP_mult_218_n1560), .C2(DP_mult_218_n1615), .A(DP_mult_218_n1632), 
        .ZN(DP_mult_218_n1631) );
  XOR2_X1 DP_mult_218_U1234 ( .A(DP_coeff_pipe02[23]), .B(DP_mult_218_n1631), 
        .Z(DP_mult_218_n1625) );
  INV_X1 DP_mult_218_U1233 ( .A(DP_mult_218_n1625), .ZN(DP_mult_218_n1621) );
  OAI21_X1 DP_mult_218_U1232 ( .B1(DP_mult_218_n1559), .B2(DP_mult_218_n1560), 
        .A(DP_mult_218_n1615), .ZN(DP_mult_218_n1630) );
  OAI221_X1 DP_mult_218_U1231 ( .B1(DP_mult_218_n1617), .B2(DP_mult_218_n1557), 
        .C1(DP_mult_218_n1617), .C2(DP_mult_218_n1558), .A(DP_mult_218_n1630), 
        .ZN(DP_mult_218_n1628) );
  XOR2_X1 DP_mult_218_U1230 ( .A(DP_mult_218_n1628), .B(DP_mult_218_n1611), 
        .Z(DP_mult_218_n1622) );
  AOI222_X1 DP_mult_218_U1229 ( .A1(DP_mult_218_n1627), .A2(DP_mult_218_n303), 
        .B1(DP_mult_218_n1625), .B2(DP_mult_218_n303), .C1(DP_mult_218_n1627), 
        .C2(DP_mult_218_n1625), .ZN(DP_mult_218_n1624) );
  INV_X1 DP_mult_218_U1228 ( .A(DP_mult_218_n1622), .ZN(DP_mult_218_n1626) );
  OAI22_X1 DP_mult_218_U1227 ( .A1(DP_mult_218_n1624), .A2(DP_mult_218_n1625), 
        .B1(DP_mult_218_n1624), .B2(DP_mult_218_n1626), .ZN(DP_mult_218_n1623)
         );
  AOI21_X1 DP_mult_218_U1226 ( .B1(DP_mult_218_n1621), .B2(DP_mult_218_n1622), 
        .A(DP_mult_218_n1623), .ZN(DP_pipe0_coeff_pipe02[23]) );
  INV_X1 DP_mult_218_U1225 ( .A(DP_mult_218_n1614), .ZN(DP_mult_218_n1620) );
  INV_X1 DP_mult_218_U1224 ( .A(DP_mult_218_n1613), .ZN(DP_mult_218_n1619) );
  INV_X1 DP_mult_218_U1223 ( .A(DP_mult_218_n1613), .ZN(DP_mult_218_n1618) );
  INV_X1 DP_mult_218_U1222 ( .A(DP_mult_218_n1612), .ZN(DP_mult_218_n1617) );
  INV_X1 DP_mult_218_U1221 ( .A(DP_mult_218_n1612), .ZN(DP_mult_218_n1616) );
  CLKBUF_X1 DP_mult_218_U1220 ( .A(DP_pipe02[23]), .Z(DP_mult_218_n1614) );
  CLKBUF_X1 DP_mult_218_U1219 ( .A(DP_pipe02[23]), .Z(DP_mult_218_n1613) );
  CLKBUF_X1 DP_mult_218_U1218 ( .A(DP_pipe02[23]), .Z(DP_mult_218_n1612) );
  INV_X1 DP_mult_218_U1217 ( .A(DP_coeff_pipe02[23]), .ZN(DP_mult_218_n1611)
         );
  BUF_X1 DP_mult_218_U1216 ( .A(DP_mult_218_n1647), .Z(DP_mult_218_n1567) );
  BUF_X1 DP_mult_218_U1215 ( .A(DP_mult_218_n1647), .Z(DP_mult_218_n1566) );
  BUF_X1 DP_mult_218_U1214 ( .A(DP_mult_218_n1647), .Z(DP_mult_218_n1565) );
  BUF_X1 DP_mult_218_U1213 ( .A(DP_coeff_pipe02[20]), .Z(DP_mult_218_n1609) );
  INV_X1 DP_mult_218_U1212 ( .A(DP_coeff_pipe02[17]), .ZN(DP_mult_218_n1607)
         );
  INV_X1 DP_mult_218_U1211 ( .A(DP_coeff_pipe02[14]), .ZN(DP_mult_218_n1605)
         );
  INV_X1 DP_mult_218_U1210 ( .A(DP_coeff_pipe02[11]), .ZN(DP_mult_218_n1603)
         );
  BUF_X1 DP_mult_218_U1209 ( .A(DP_coeff_pipe02[20]), .Z(DP_mult_218_n1608) );
  INV_X1 DP_mult_218_U1208 ( .A(DP_mult_218_n1611), .ZN(DP_mult_218_n1610) );
  INV_X1 DP_mult_218_U1207 ( .A(DP_mult_218_n1616), .ZN(DP_mult_218_n1615) );
  OR2_X1 DP_mult_218_U1206 ( .A1(DP_mult_218_n1904), .A2(DP_mult_218_n1905), 
        .ZN(DP_mult_218_n1555) );
  AND2_X1 DP_mult_218_U1205 ( .A1(DP_coeff_pipe02[0]), .A2(DP_mult_218_n2157), 
        .ZN(DP_mult_218_n1554) );
  INV_X1 DP_mult_218_U1204 ( .A(DP_mult_218_n1603), .ZN(DP_mult_218_n1602) );
  AND2_X1 DP_mult_218_U1203 ( .A1(DP_mult_218_n2070), .A2(DP_mult_218_n2068), 
        .ZN(DP_mult_218_n1553) );
  OR2_X1 DP_mult_218_U1202 ( .A1(DP_mult_218_n2014), .A2(DP_mult_218_n2015), 
        .ZN(DP_mult_218_n1552) );
  OR2_X1 DP_mult_218_U1201 ( .A1(DP_mult_218_n1959), .A2(DP_mult_218_n1960), 
        .ZN(DP_mult_218_n1551) );
  OR2_X1 DP_mult_218_U1200 ( .A1(DP_mult_218_n2070), .A2(DP_mult_218_n2069), 
        .ZN(DP_mult_218_n1550) );
  AND2_X1 DP_mult_218_U1199 ( .A1(DP_mult_218_n1959), .A2(DP_mult_218_n1961), 
        .ZN(DP_mult_218_n1549) );
  AND2_X1 DP_mult_218_U1198 ( .A1(DP_mult_218_n1904), .A2(DP_mult_218_n1906), 
        .ZN(DP_mult_218_n1548) );
  AND2_X1 DP_mult_218_U1197 ( .A1(DP_mult_218_n2014), .A2(DP_mult_218_n2016), 
        .ZN(DP_mult_218_n1547) );
  OR2_X1 DP_mult_218_U1196 ( .A1(DP_mult_218_n1961), .A2(DP_mult_218_n1962), 
        .ZN(DP_mult_218_n1546) );
  OR2_X1 DP_mult_218_U1195 ( .A1(DP_mult_218_n1906), .A2(DP_mult_218_n1907), 
        .ZN(DP_mult_218_n1545) );
  OR2_X1 DP_mult_218_U1194 ( .A1(DP_mult_218_n2068), .A2(DP_mult_218_n2067), 
        .ZN(DP_mult_218_n1544) );
  OR2_X1 DP_mult_218_U1193 ( .A1(DP_mult_218_n2016), .A2(DP_mult_218_n2017), 
        .ZN(DP_mult_218_n1543) );
  INV_X1 DP_mult_218_U1192 ( .A(DP_mult_218_n1607), .ZN(DP_mult_218_n1606) );
  INV_X1 DP_mult_218_U1191 ( .A(DP_mult_218_n1605), .ZN(DP_mult_218_n1604) );
  BUF_X1 DP_mult_218_U1190 ( .A(DP_mult_218_n1636), .Z(DP_mult_218_n1562) );
  OR2_X1 DP_mult_218_U1189 ( .A1(DP_mult_218_n2158), .A2(DP_mult_218_n2157), 
        .ZN(DP_mult_218_n1542) );
  BUF_X1 DP_mult_218_U1188 ( .A(DP_mult_218_n1629), .Z(DP_mult_218_n1556) );
  BUF_X1 DP_mult_218_U1187 ( .A(DP_mult_218_n1636), .Z(DP_mult_218_n1563) );
  INV_X1 DP_mult_218_U1186 ( .A(DP_mult_218_n1554), .ZN(DP_mult_218_n1564) );
  INV_X1 DP_mult_218_U1185 ( .A(DP_mult_218_n1543), .ZN(DP_mult_218_n1594) );
  INV_X1 DP_mult_218_U1184 ( .A(DP_mult_218_n1546), .ZN(DP_mult_218_n1589) );
  INV_X1 DP_mult_218_U1183 ( .A(DP_mult_218_n1545), .ZN(DP_mult_218_n1584) );
  INV_X1 DP_mult_218_U1182 ( .A(DP_mult_218_n1555), .ZN(DP_mult_218_n1585) );
  NAND3_X1 DP_mult_218_U1181 ( .A1(DP_mult_218_n2157), .A2(DP_mult_218_n2158), 
        .A3(DP_mult_218_n2159), .ZN(DP_mult_218_n1639) );
  AND2_X1 DP_mult_218_U1180 ( .A1(DP_mult_218_n1849), .A2(DP_mult_218_n1851), 
        .ZN(DP_mult_218_n1541) );
  OR2_X1 DP_mult_218_U1179 ( .A1(DP_mult_218_n1851), .A2(DP_mult_218_n1852), 
        .ZN(DP_mult_218_n1540) );
  BUF_X1 DP_mult_218_U1178 ( .A(DP_mult_218_n1967), .Z(DP_mult_218_n1597) );
  BUF_X1 DP_mult_218_U1177 ( .A(DP_mult_218_n1912), .Z(DP_mult_218_n1592) );
  BUF_X1 DP_mult_218_U1176 ( .A(DP_mult_218_n1857), .Z(DP_mult_218_n1587) );
  BUF_X1 DP_mult_218_U1175 ( .A(DP_mult_218_n1912), .Z(DP_mult_218_n1591) );
  BUF_X1 DP_mult_218_U1174 ( .A(DP_mult_218_n1967), .Z(DP_mult_218_n1596) );
  BUF_X1 DP_mult_218_U1173 ( .A(DP_mult_218_n1857), .Z(DP_mult_218_n1586) );
  BUF_X1 DP_mult_218_U1172 ( .A(DP_mult_218_n1629), .Z(DP_mult_218_n1557) );
  INV_X1 DP_mult_218_U1171 ( .A(DP_mult_218_n1547), .ZN(DP_mult_218_n1593) );
  INV_X1 DP_mult_218_U1170 ( .A(DP_mult_218_n1548), .ZN(DP_mult_218_n1583) );
  INV_X1 DP_mult_218_U1169 ( .A(DP_mult_218_n1549), .ZN(DP_mult_218_n1588) );
  INV_X1 DP_mult_218_U1168 ( .A(DP_mult_218_n1544), .ZN(DP_mult_218_n1559) );
  INV_X1 DP_mult_218_U1167 ( .A(DP_mult_218_n1552), .ZN(DP_mult_218_n1595) );
  INV_X1 DP_mult_218_U1166 ( .A(DP_mult_218_n1551), .ZN(DP_mult_218_n1590) );
  INV_X1 DP_mult_218_U1165 ( .A(DP_mult_218_n1553), .ZN(DP_mult_218_n1558) );
  INV_X1 DP_mult_218_U1164 ( .A(DP_mult_218_n1550), .ZN(DP_mult_218_n1560) );
  INV_X1 DP_mult_218_U1163 ( .A(DP_mult_218_n1540), .ZN(DP_mult_218_n1579) );
  INV_X1 DP_mult_218_U1162 ( .A(DP_coeff_pipe02[8]), .ZN(DP_mult_218_n1601) );
  INV_X1 DP_mult_218_U1161 ( .A(DP_coeff_pipe02[5]), .ZN(DP_mult_218_n1599) );
  BUF_X1 DP_mult_218_U1160 ( .A(DP_mult_218_n1802), .Z(DP_mult_218_n1582) );
  BUF_X1 DP_mult_218_U1159 ( .A(DP_mult_218_n1802), .Z(DP_mult_218_n1581) );
  OR2_X1 DP_mult_218_U1158 ( .A1(DP_mult_218_n1738), .A2(DP_mult_218_n1739), 
        .ZN(DP_mult_218_n1539) );
  OR2_X1 DP_mult_218_U1157 ( .A1(DP_mult_218_n1740), .A2(DP_mult_218_n1741), 
        .ZN(DP_mult_218_n1538) );
  INV_X1 DP_mult_218_U1156 ( .A(DP_mult_218_n1542), .ZN(DP_mult_218_n1561) );
  INV_X1 DP_mult_218_U1155 ( .A(DP_mult_218_n1541), .ZN(DP_mult_218_n1578) );
  AND2_X1 DP_mult_218_U1154 ( .A1(DP_mult_218_n1738), .A2(DP_mult_218_n1740), 
        .ZN(DP_mult_218_n1537) );
  BUF_X1 DP_mult_218_U1153 ( .A(DP_mult_218_n1654), .Z(DP_mult_218_n1572) );
  BUF_X1 DP_mult_218_U1152 ( .A(DP_mult_218_n1654), .Z(DP_mult_218_n1571) );
  INV_X1 DP_mult_218_U1151 ( .A(DP_mult_218_n1538), .ZN(DP_mult_218_n1569) );
  INV_X1 DP_mult_218_U1150 ( .A(DP_mult_218_n1539), .ZN(DP_mult_218_n1570) );
  INV_X1 DP_mult_218_U1149 ( .A(DP_mult_218_n1601), .ZN(DP_mult_218_n1600) );
  INV_X1 DP_mult_218_U1148 ( .A(DP_mult_218_n1599), .ZN(DP_mult_218_n1598) );
  OR2_X1 DP_mult_218_U1147 ( .A1(DP_mult_218_n1794), .A2(DP_mult_218_n1795), 
        .ZN(DP_mult_218_n1536) );
  AND2_X1 DP_mult_218_U1146 ( .A1(DP_mult_218_n1794), .A2(DP_mult_218_n1796), 
        .ZN(DP_mult_218_n1535) );
  OR2_X1 DP_mult_218_U1145 ( .A1(DP_mult_218_n1796), .A2(DP_mult_218_n1797), 
        .ZN(DP_mult_218_n1534) );
  INV_X1 DP_mult_218_U1144 ( .A(DP_mult_218_n1537), .ZN(DP_mult_218_n1568) );
  INV_X1 DP_mult_218_U1143 ( .A(DP_mult_218_n1534), .ZN(DP_mult_218_n1574) );
  OR2_X1 DP_mult_218_U1142 ( .A1(DP_mult_218_n1849), .A2(DP_mult_218_n1850), 
        .ZN(DP_mult_218_n1533) );
  BUF_X1 DP_mult_218_U1141 ( .A(DP_mult_218_n1747), .Z(DP_mult_218_n1577) );
  BUF_X1 DP_mult_218_U1140 ( .A(DP_mult_218_n1747), .Z(DP_mult_218_n1576) );
  INV_X1 DP_mult_218_U1139 ( .A(DP_mult_218_n1535), .ZN(DP_mult_218_n1573) );
  INV_X1 DP_mult_218_U1138 ( .A(DP_mult_218_n1536), .ZN(DP_mult_218_n1575) );
  INV_X1 DP_mult_218_U1137 ( .A(DP_mult_218_n1533), .ZN(DP_mult_218_n1580) );
  HA_X1 DP_mult_218_U1134 ( .A(DP_pipe02[0]), .B(DP_pipe02[1]), .CO(
        DP_mult_218_n727), .S(DP_mult_218_n1397) );
  FA_X1 DP_mult_218_U1133 ( .A(DP_pipe02[1]), .B(DP_pipe02[2]), .CI(
        DP_mult_218_n727), .CO(DP_mult_218_n726), .S(DP_mult_218_n1396) );
  FA_X1 DP_mult_218_U1132 ( .A(DP_pipe02[2]), .B(DP_pipe02[3]), .CI(
        DP_mult_218_n726), .CO(DP_mult_218_n725), .S(DP_mult_218_n1395) );
  FA_X1 DP_mult_218_U1131 ( .A(DP_pipe02[3]), .B(DP_pipe02[4]), .CI(
        DP_mult_218_n725), .CO(DP_mult_218_n724), .S(DP_mult_218_n1394) );
  FA_X1 DP_mult_218_U1130 ( .A(DP_pipe02[4]), .B(DP_pipe02[5]), .CI(
        DP_mult_218_n724), .CO(DP_mult_218_n723), .S(DP_mult_218_n1393) );
  FA_X1 DP_mult_218_U1129 ( .A(DP_pipe02[5]), .B(DP_pipe02[6]), .CI(
        DP_mult_218_n723), .CO(DP_mult_218_n722), .S(DP_mult_218_n1392) );
  FA_X1 DP_mult_218_U1128 ( .A(DP_pipe02[6]), .B(DP_pipe02[7]), .CI(
        DP_mult_218_n722), .CO(DP_mult_218_n721), .S(DP_mult_218_n1391) );
  FA_X1 DP_mult_218_U1127 ( .A(DP_pipe02[7]), .B(DP_pipe02[8]), .CI(
        DP_mult_218_n721), .CO(DP_mult_218_n720), .S(DP_mult_218_n1390) );
  FA_X1 DP_mult_218_U1126 ( .A(DP_pipe02[8]), .B(DP_pipe02[9]), .CI(
        DP_mult_218_n720), .CO(DP_mult_218_n719), .S(DP_mult_218_n1389) );
  FA_X1 DP_mult_218_U1125 ( .A(DP_pipe02[9]), .B(DP_pipe02[10]), .CI(
        DP_mult_218_n719), .CO(DP_mult_218_n718), .S(DP_mult_218_n1388) );
  FA_X1 DP_mult_218_U1124 ( .A(DP_pipe02[10]), .B(DP_pipe02[11]), .CI(
        DP_mult_218_n718), .CO(DP_mult_218_n717), .S(DP_mult_218_n1387) );
  FA_X1 DP_mult_218_U1123 ( .A(DP_pipe02[11]), .B(DP_pipe02[12]), .CI(
        DP_mult_218_n717), .CO(DP_mult_218_n716), .S(DP_mult_218_n1386) );
  FA_X1 DP_mult_218_U1122 ( .A(DP_pipe02[12]), .B(DP_pipe02[13]), .CI(
        DP_mult_218_n716), .CO(DP_mult_218_n715), .S(DP_mult_218_n1385) );
  FA_X1 DP_mult_218_U1121 ( .A(DP_pipe02[13]), .B(DP_pipe02[14]), .CI(
        DP_mult_218_n715), .CO(DP_mult_218_n714), .S(DP_mult_218_n1384) );
  FA_X1 DP_mult_218_U1120 ( .A(DP_pipe02[14]), .B(DP_pipe02[15]), .CI(
        DP_mult_218_n714), .CO(DP_mult_218_n713), .S(DP_mult_218_n1383) );
  FA_X1 DP_mult_218_U1119 ( .A(DP_pipe02[15]), .B(DP_pipe02[16]), .CI(
        DP_mult_218_n713), .CO(DP_mult_218_n712), .S(DP_mult_218_n1382) );
  FA_X1 DP_mult_218_U1118 ( .A(DP_pipe02[16]), .B(DP_pipe02[17]), .CI(
        DP_mult_218_n712), .CO(DP_mult_218_n711), .S(DP_mult_218_n1381) );
  FA_X1 DP_mult_218_U1117 ( .A(DP_pipe02[17]), .B(DP_pipe02[18]), .CI(
        DP_mult_218_n711), .CO(DP_mult_218_n710), .S(DP_mult_218_n1380) );
  FA_X1 DP_mult_218_U1116 ( .A(DP_pipe02[18]), .B(DP_pipe02[19]), .CI(
        DP_mult_218_n710), .CO(DP_mult_218_n709), .S(DP_mult_218_n1379) );
  FA_X1 DP_mult_218_U1115 ( .A(DP_pipe02[19]), .B(DP_pipe02[20]), .CI(
        DP_mult_218_n709), .CO(DP_mult_218_n708), .S(DP_mult_218_n1378) );
  FA_X1 DP_mult_218_U1114 ( .A(DP_pipe02[20]), .B(DP_pipe02[21]), .CI(
        DP_mult_218_n708), .CO(DP_mult_218_n707), .S(DP_mult_218_n1377) );
  FA_X1 DP_mult_218_U1113 ( .A(DP_pipe02[21]), .B(DP_pipe02[22]), .CI(
        DP_mult_218_n707), .CO(DP_mult_218_n706), .S(DP_mult_218_n1376) );
  FA_X1 DP_mult_218_U1112 ( .A(DP_pipe02[22]), .B(DP_mult_218_n1615), .CI(
        DP_mult_218_n706), .CO(DP_mult_218_n1374), .S(DP_mult_218_n1375) );
  HA_X1 DP_mult_218_U408 ( .A(DP_mult_218_n904), .B(DP_mult_218_n1598), .CO(
        DP_mult_218_n687), .S(DP_mult_218_n688) );
  HA_X1 DP_mult_218_U407 ( .A(DP_mult_218_n687), .B(DP_mult_218_n903), .CO(
        DP_mult_218_n685), .S(DP_mult_218_n686) );
  HA_X1 DP_mult_218_U406 ( .A(DP_mult_218_n685), .B(DP_mult_218_n902), .CO(
        DP_mult_218_n683), .S(DP_mult_218_n684) );
  HA_X1 DP_mult_218_U405 ( .A(DP_mult_218_n878), .B(DP_mult_218_n1600), .CO(
        DP_mult_218_n681), .S(DP_mult_218_n682) );
  FA_X1 DP_mult_218_U404 ( .A(DP_mult_218_n901), .B(DP_mult_218_n682), .CI(
        DP_mult_218_n683), .CO(DP_mult_218_n679), .S(DP_mult_218_n680) );
  HA_X1 DP_mult_218_U403 ( .A(DP_mult_218_n681), .B(DP_mult_218_n877), .CO(
        DP_mult_218_n677), .S(DP_mult_218_n678) );
  FA_X1 DP_mult_218_U402 ( .A(DP_mult_218_n900), .B(DP_mult_218_n678), .CI(
        DP_mult_218_n679), .CO(DP_mult_218_n675), .S(DP_mult_218_n676) );
  HA_X1 DP_mult_218_U401 ( .A(DP_mult_218_n677), .B(DP_mult_218_n876), .CO(
        DP_mult_218_n673), .S(DP_mult_218_n674) );
  FA_X1 DP_mult_218_U400 ( .A(DP_mult_218_n899), .B(DP_mult_218_n674), .CI(
        DP_mult_218_n675), .CO(DP_mult_218_n671), .S(DP_mult_218_n672) );
  HA_X1 DP_mult_218_U399 ( .A(DP_mult_218_n852), .B(DP_mult_218_n1602), .CO(
        DP_mult_218_n669), .S(DP_mult_218_n670) );
  FA_X1 DP_mult_218_U398 ( .A(DP_mult_218_n875), .B(DP_mult_218_n670), .CI(
        DP_mult_218_n673), .CO(DP_mult_218_n667), .S(DP_mult_218_n668) );
  FA_X1 DP_mult_218_U397 ( .A(DP_mult_218_n898), .B(DP_mult_218_n668), .CI(
        DP_mult_218_n671), .CO(DP_mult_218_n665), .S(DP_mult_218_n666) );
  HA_X1 DP_mult_218_U396 ( .A(DP_mult_218_n669), .B(DP_mult_218_n851), .CO(
        DP_mult_218_n663), .S(DP_mult_218_n664) );
  FA_X1 DP_mult_218_U395 ( .A(DP_mult_218_n874), .B(DP_mult_218_n664), .CI(
        DP_mult_218_n667), .CO(DP_mult_218_n661), .S(DP_mult_218_n662) );
  FA_X1 DP_mult_218_U394 ( .A(DP_mult_218_n897), .B(DP_mult_218_n662), .CI(
        DP_mult_218_n665), .CO(DP_mult_218_n659), .S(DP_mult_218_n660) );
  HA_X1 DP_mult_218_U393 ( .A(DP_mult_218_n663), .B(DP_mult_218_n850), .CO(
        DP_mult_218_n657), .S(DP_mult_218_n658) );
  FA_X1 DP_mult_218_U392 ( .A(DP_mult_218_n873), .B(DP_mult_218_n658), .CI(
        DP_mult_218_n661), .CO(DP_mult_218_n655), .S(DP_mult_218_n656) );
  FA_X1 DP_mult_218_U391 ( .A(DP_mult_218_n896), .B(DP_mult_218_n656), .CI(
        DP_mult_218_n659), .CO(DP_mult_218_n653), .S(DP_mult_218_n654) );
  HA_X1 DP_mult_218_U390 ( .A(DP_mult_218_n826), .B(DP_mult_218_n1604), .CO(
        DP_mult_218_n651), .S(DP_mult_218_n652) );
  FA_X1 DP_mult_218_U389 ( .A(DP_mult_218_n849), .B(DP_mult_218_n652), .CI(
        DP_mult_218_n657), .CO(DP_mult_218_n649), .S(DP_mult_218_n650) );
  FA_X1 DP_mult_218_U388 ( .A(DP_mult_218_n872), .B(DP_mult_218_n650), .CI(
        DP_mult_218_n655), .CO(DP_mult_218_n647), .S(DP_mult_218_n648) );
  FA_X1 DP_mult_218_U387 ( .A(DP_mult_218_n895), .B(DP_mult_218_n648), .CI(
        DP_mult_218_n653), .CO(DP_mult_218_n645), .S(DP_mult_218_n646) );
  HA_X1 DP_mult_218_U386 ( .A(DP_mult_218_n651), .B(DP_mult_218_n825), .CO(
        DP_mult_218_n643), .S(DP_mult_218_n644) );
  FA_X1 DP_mult_218_U385 ( .A(DP_mult_218_n848), .B(DP_mult_218_n644), .CI(
        DP_mult_218_n649), .CO(DP_mult_218_n641), .S(DP_mult_218_n642) );
  FA_X1 DP_mult_218_U384 ( .A(DP_mult_218_n871), .B(DP_mult_218_n642), .CI(
        DP_mult_218_n647), .CO(DP_mult_218_n639), .S(DP_mult_218_n640) );
  FA_X1 DP_mult_218_U383 ( .A(DP_mult_218_n894), .B(DP_mult_218_n640), .CI(
        DP_mult_218_n645), .CO(DP_mult_218_n637), .S(DP_mult_218_n638) );
  HA_X1 DP_mult_218_U382 ( .A(DP_mult_218_n643), .B(DP_mult_218_n824), .CO(
        DP_mult_218_n635), .S(DP_mult_218_n636) );
  FA_X1 DP_mult_218_U381 ( .A(DP_mult_218_n847), .B(DP_mult_218_n636), .CI(
        DP_mult_218_n641), .CO(DP_mult_218_n633), .S(DP_mult_218_n634) );
  FA_X1 DP_mult_218_U380 ( .A(DP_mult_218_n870), .B(DP_mult_218_n634), .CI(
        DP_mult_218_n639), .CO(DP_mult_218_n631), .S(DP_mult_218_n632) );
  FA_X1 DP_mult_218_U379 ( .A(DP_mult_218_n893), .B(DP_mult_218_n632), .CI(
        DP_mult_218_n637), .CO(DP_mult_218_n629), .S(DP_mult_218_n630) );
  HA_X1 DP_mult_218_U378 ( .A(DP_mult_218_n800), .B(DP_mult_218_n1606), .CO(
        DP_mult_218_n627), .S(DP_mult_218_n628) );
  FA_X1 DP_mult_218_U377 ( .A(DP_mult_218_n823), .B(DP_mult_218_n628), .CI(
        DP_mult_218_n635), .CO(DP_mult_218_n625), .S(DP_mult_218_n626) );
  FA_X1 DP_mult_218_U376 ( .A(DP_mult_218_n846), .B(DP_mult_218_n626), .CI(
        DP_mult_218_n633), .CO(DP_mult_218_n623), .S(DP_mult_218_n624) );
  FA_X1 DP_mult_218_U375 ( .A(DP_mult_218_n869), .B(DP_mult_218_n624), .CI(
        DP_mult_218_n631), .CO(DP_mult_218_n621), .S(DP_mult_218_n622) );
  FA_X1 DP_mult_218_U374 ( .A(DP_mult_218_n892), .B(DP_mult_218_n622), .CI(
        DP_mult_218_n629), .CO(DP_mult_218_n619), .S(DP_mult_218_n620) );
  HA_X1 DP_mult_218_U373 ( .A(DP_mult_218_n627), .B(DP_mult_218_n799), .CO(
        DP_mult_218_n617), .S(DP_mult_218_n618) );
  FA_X1 DP_mult_218_U372 ( .A(DP_mult_218_n822), .B(DP_mult_218_n618), .CI(
        DP_mult_218_n625), .CO(DP_mult_218_n615), .S(DP_mult_218_n616) );
  FA_X1 DP_mult_218_U371 ( .A(DP_mult_218_n845), .B(DP_mult_218_n616), .CI(
        DP_mult_218_n623), .CO(DP_mult_218_n613), .S(DP_mult_218_n614) );
  FA_X1 DP_mult_218_U370 ( .A(DP_mult_218_n868), .B(DP_mult_218_n614), .CI(
        DP_mult_218_n621), .CO(DP_mult_218_n611), .S(DP_mult_218_n612) );
  FA_X1 DP_mult_218_U369 ( .A(DP_mult_218_n891), .B(DP_mult_218_n612), .CI(
        DP_mult_218_n619), .CO(DP_mult_218_n609), .S(DP_mult_218_n610) );
  HA_X1 DP_mult_218_U368 ( .A(DP_mult_218_n617), .B(DP_mult_218_n798), .CO(
        DP_mult_218_n607), .S(DP_mult_218_n608) );
  FA_X1 DP_mult_218_U367 ( .A(DP_mult_218_n821), .B(DP_mult_218_n608), .CI(
        DP_mult_218_n615), .CO(DP_mult_218_n605), .S(DP_mult_218_n606) );
  FA_X1 DP_mult_218_U366 ( .A(DP_mult_218_n844), .B(DP_mult_218_n606), .CI(
        DP_mult_218_n613), .CO(DP_mult_218_n603), .S(DP_mult_218_n604) );
  FA_X1 DP_mult_218_U365 ( .A(DP_mult_218_n867), .B(DP_mult_218_n604), .CI(
        DP_mult_218_n611), .CO(DP_mult_218_n601), .S(DP_mult_218_n602) );
  FA_X1 DP_mult_218_U364 ( .A(DP_mult_218_n890), .B(DP_mult_218_n602), .CI(
        DP_mult_218_n609), .CO(DP_mult_218_n599), .S(DP_mult_218_n600) );
  HA_X1 DP_mult_218_U363 ( .A(DP_mult_218_n774), .B(DP_mult_218_n1608), .CO(
        DP_mult_218_n597), .S(DP_mult_218_n598) );
  FA_X1 DP_mult_218_U362 ( .A(DP_mult_218_n797), .B(DP_mult_218_n598), .CI(
        DP_mult_218_n607), .CO(DP_mult_218_n595), .S(DP_mult_218_n596) );
  FA_X1 DP_mult_218_U361 ( .A(DP_mult_218_n820), .B(DP_mult_218_n596), .CI(
        DP_mult_218_n605), .CO(DP_mult_218_n593), .S(DP_mult_218_n594) );
  FA_X1 DP_mult_218_U360 ( .A(DP_mult_218_n843), .B(DP_mult_218_n594), .CI(
        DP_mult_218_n603), .CO(DP_mult_218_n591), .S(DP_mult_218_n592) );
  FA_X1 DP_mult_218_U359 ( .A(DP_mult_218_n866), .B(DP_mult_218_n592), .CI(
        DP_mult_218_n601), .CO(DP_mult_218_n589), .S(DP_mult_218_n590) );
  FA_X1 DP_mult_218_U358 ( .A(DP_mult_218_n889), .B(DP_mult_218_n590), .CI(
        DP_mult_218_n599), .CO(DP_mult_218_n587), .S(DP_mult_218_n588) );
  HA_X1 DP_mult_218_U357 ( .A(DP_mult_218_n597), .B(DP_mult_218_n773), .CO(
        DP_mult_218_n585), .S(DP_mult_218_n586) );
  FA_X1 DP_mult_218_U356 ( .A(DP_mult_218_n796), .B(DP_mult_218_n586), .CI(
        DP_mult_218_n595), .CO(DP_mult_218_n583), .S(DP_mult_218_n584) );
  FA_X1 DP_mult_218_U355 ( .A(DP_mult_218_n819), .B(DP_mult_218_n584), .CI(
        DP_mult_218_n593), .CO(DP_mult_218_n581), .S(DP_mult_218_n582) );
  FA_X1 DP_mult_218_U354 ( .A(DP_mult_218_n842), .B(DP_mult_218_n582), .CI(
        DP_mult_218_n591), .CO(DP_mult_218_n579), .S(DP_mult_218_n580) );
  FA_X1 DP_mult_218_U353 ( .A(DP_mult_218_n865), .B(DP_mult_218_n580), .CI(
        DP_mult_218_n589), .CO(DP_mult_218_n577), .S(DP_mult_218_n578) );
  FA_X1 DP_mult_218_U352 ( .A(DP_mult_218_n888), .B(DP_mult_218_n578), .CI(
        DP_mult_218_n587), .CO(DP_mult_218_n575), .S(DP_mult_218_n576) );
  HA_X1 DP_mult_218_U351 ( .A(DP_mult_218_n585), .B(DP_mult_218_n772), .CO(
        DP_mult_218_n573), .S(DP_mult_218_n574) );
  FA_X1 DP_mult_218_U350 ( .A(DP_mult_218_n795), .B(DP_mult_218_n574), .CI(
        DP_mult_218_n583), .CO(DP_mult_218_n571), .S(DP_mult_218_n572) );
  FA_X1 DP_mult_218_U349 ( .A(DP_mult_218_n818), .B(DP_mult_218_n572), .CI(
        DP_mult_218_n581), .CO(DP_mult_218_n569), .S(DP_mult_218_n570) );
  FA_X1 DP_mult_218_U348 ( .A(DP_mult_218_n841), .B(DP_mult_218_n570), .CI(
        DP_mult_218_n579), .CO(DP_mult_218_n567), .S(DP_mult_218_n568) );
  FA_X1 DP_mult_218_U347 ( .A(DP_mult_218_n864), .B(DP_mult_218_n568), .CI(
        DP_mult_218_n577), .CO(DP_mult_218_n565), .S(DP_mult_218_n566) );
  FA_X1 DP_mult_218_U346 ( .A(DP_mult_218_n887), .B(DP_mult_218_n566), .CI(
        DP_mult_218_n575), .CO(DP_mult_218_n563), .S(DP_mult_218_n564) );
  HA_X1 DP_mult_218_U345 ( .A(DP_mult_218_n748), .B(DP_mult_218_n1610), .CO(
        DP_mult_218_n561), .S(DP_mult_218_n562) );
  FA_X1 DP_mult_218_U344 ( .A(DP_mult_218_n771), .B(DP_mult_218_n562), .CI(
        DP_mult_218_n573), .CO(DP_mult_218_n559), .S(DP_mult_218_n560) );
  FA_X1 DP_mult_218_U343 ( .A(DP_mult_218_n794), .B(DP_mult_218_n560), .CI(
        DP_mult_218_n571), .CO(DP_mult_218_n557), .S(DP_mult_218_n558) );
  FA_X1 DP_mult_218_U342 ( .A(DP_mult_218_n817), .B(DP_mult_218_n558), .CI(
        DP_mult_218_n569), .CO(DP_mult_218_n555), .S(DP_mult_218_n556) );
  FA_X1 DP_mult_218_U341 ( .A(DP_mult_218_n840), .B(DP_mult_218_n556), .CI(
        DP_mult_218_n567), .CO(DP_mult_218_n553), .S(DP_mult_218_n554) );
  FA_X1 DP_mult_218_U340 ( .A(DP_mult_218_n863), .B(DP_mult_218_n554), .CI(
        DP_mult_218_n565), .CO(DP_mult_218_n551), .S(DP_mult_218_n552) );
  FA_X1 DP_mult_218_U339 ( .A(DP_mult_218_n886), .B(DP_mult_218_n552), .CI(
        DP_mult_218_n563), .CO(DP_mult_218_n549), .S(DP_mult_218_n550) );
  HA_X1 DP_mult_218_U338 ( .A(DP_mult_218_n561), .B(DP_mult_218_n747), .CO(
        DP_mult_218_n547), .S(DP_mult_218_n548) );
  FA_X1 DP_mult_218_U337 ( .A(DP_mult_218_n770), .B(DP_mult_218_n548), .CI(
        DP_mult_218_n559), .CO(DP_mult_218_n545), .S(DP_mult_218_n546) );
  FA_X1 DP_mult_218_U336 ( .A(DP_mult_218_n793), .B(DP_mult_218_n546), .CI(
        DP_mult_218_n557), .CO(DP_mult_218_n543), .S(DP_mult_218_n544) );
  FA_X1 DP_mult_218_U335 ( .A(DP_mult_218_n816), .B(DP_mult_218_n544), .CI(
        DP_mult_218_n555), .CO(DP_mult_218_n541), .S(DP_mult_218_n542) );
  FA_X1 DP_mult_218_U334 ( .A(DP_mult_218_n839), .B(DP_mult_218_n542), .CI(
        DP_mult_218_n553), .CO(DP_mult_218_n539), .S(DP_mult_218_n540) );
  FA_X1 DP_mult_218_U333 ( .A(DP_mult_218_n862), .B(DP_mult_218_n540), .CI(
        DP_mult_218_n551), .CO(DP_mult_218_n537), .S(DP_mult_218_n538) );
  FA_X1 DP_mult_218_U332 ( .A(DP_mult_218_n885), .B(DP_mult_218_n538), .CI(
        DP_mult_218_n549), .CO(DP_mult_218_n535), .S(DP_mult_218_n536) );
  HA_X1 DP_mult_218_U331 ( .A(DP_mult_218_n547), .B(DP_mult_218_n746), .CO(
        DP_mult_218_n533), .S(DP_mult_218_n534) );
  FA_X1 DP_mult_218_U330 ( .A(DP_mult_218_n769), .B(DP_mult_218_n534), .CI(
        DP_mult_218_n545), .CO(DP_mult_218_n531), .S(DP_mult_218_n532) );
  FA_X1 DP_mult_218_U329 ( .A(DP_mult_218_n792), .B(DP_mult_218_n532), .CI(
        DP_mult_218_n543), .CO(DP_mult_218_n529), .S(DP_mult_218_n530) );
  FA_X1 DP_mult_218_U328 ( .A(DP_mult_218_n815), .B(DP_mult_218_n530), .CI(
        DP_mult_218_n541), .CO(DP_mult_218_n527), .S(DP_mult_218_n528) );
  FA_X1 DP_mult_218_U327 ( .A(DP_mult_218_n838), .B(DP_mult_218_n528), .CI(
        DP_mult_218_n539), .CO(DP_mult_218_n525), .S(DP_mult_218_n526) );
  FA_X1 DP_mult_218_U326 ( .A(DP_mult_218_n861), .B(DP_mult_218_n526), .CI(
        DP_mult_218_n537), .CO(DP_mult_218_n523), .S(DP_mult_218_n524) );
  FA_X1 DP_mult_218_U325 ( .A(DP_mult_218_n884), .B(DP_mult_218_n524), .CI(
        DP_mult_218_n535), .CO(DP_mult_218_n521), .S(DP_mult_218_n522) );
  HA_X1 DP_mult_218_U324 ( .A(DP_mult_218_n533), .B(DP_mult_218_n745), .CO(
        DP_mult_218_n519), .S(DP_mult_218_n520) );
  FA_X1 DP_mult_218_U323 ( .A(DP_mult_218_n768), .B(DP_mult_218_n520), .CI(
        DP_mult_218_n531), .CO(DP_mult_218_n517), .S(DP_mult_218_n518) );
  FA_X1 DP_mult_218_U322 ( .A(DP_mult_218_n791), .B(DP_mult_218_n518), .CI(
        DP_mult_218_n529), .CO(DP_mult_218_n515), .S(DP_mult_218_n516) );
  FA_X1 DP_mult_218_U321 ( .A(DP_mult_218_n814), .B(DP_mult_218_n516), .CI(
        DP_mult_218_n527), .CO(DP_mult_218_n513), .S(DP_mult_218_n514) );
  FA_X1 DP_mult_218_U320 ( .A(DP_mult_218_n837), .B(DP_mult_218_n514), .CI(
        DP_mult_218_n525), .CO(DP_mult_218_n511), .S(DP_mult_218_n512) );
  FA_X1 DP_mult_218_U319 ( .A(DP_mult_218_n860), .B(DP_mult_218_n512), .CI(
        DP_mult_218_n523), .CO(DP_mult_218_n509), .S(DP_mult_218_n510) );
  FA_X1 DP_mult_218_U318 ( .A(DP_mult_218_n883), .B(DP_mult_218_n510), .CI(
        DP_mult_218_n521), .CO(DP_mult_218_n507), .S(DP_mult_218_n508) );
  FA_X1 DP_mult_218_U315 ( .A(DP_mult_218_n506), .B(DP_mult_218_n744), .CI(
        DP_mult_218_n767), .CO(DP_mult_218_n504), .S(DP_mult_218_n505) );
  FA_X1 DP_mult_218_U314 ( .A(DP_mult_218_n505), .B(DP_mult_218_n517), .CI(
        DP_mult_218_n790), .CO(DP_mult_218_n502), .S(DP_mult_218_n503) );
  FA_X1 DP_mult_218_U313 ( .A(DP_mult_218_n503), .B(DP_mult_218_n515), .CI(
        DP_mult_218_n813), .CO(DP_mult_218_n500), .S(DP_mult_218_n501) );
  FA_X1 DP_mult_218_U312 ( .A(DP_mult_218_n501), .B(DP_mult_218_n513), .CI(
        DP_mult_218_n836), .CO(DP_mult_218_n498), .S(DP_mult_218_n499) );
  FA_X1 DP_mult_218_U311 ( .A(DP_mult_218_n499), .B(DP_mult_218_n511), .CI(
        DP_mult_218_n859), .CO(DP_mult_218_n496), .S(DP_mult_218_n497) );
  FA_X1 DP_mult_218_U310 ( .A(DP_mult_218_n497), .B(DP_mult_218_n509), .CI(
        DP_mult_218_n882), .CO(DP_mult_218_n494), .S(DP_mult_218_n495) );
  FA_X1 DP_mult_218_U308 ( .A(DP_mult_218_n743), .B(DP_mult_218_n493), .CI(
        DP_mult_218_n766), .CO(DP_mult_218_n491), .S(DP_mult_218_n492) );
  FA_X1 DP_mult_218_U307 ( .A(DP_mult_218_n492), .B(DP_mult_218_n504), .CI(
        DP_mult_218_n789), .CO(DP_mult_218_n489), .S(DP_mult_218_n490) );
  FA_X1 DP_mult_218_U306 ( .A(DP_mult_218_n490), .B(DP_mult_218_n502), .CI(
        DP_mult_218_n500), .CO(DP_mult_218_n487), .S(DP_mult_218_n488) );
  FA_X1 DP_mult_218_U305 ( .A(DP_mult_218_n488), .B(DP_mult_218_n812), .CI(
        DP_mult_218_n835), .CO(DP_mult_218_n485), .S(DP_mult_218_n486) );
  FA_X1 DP_mult_218_U304 ( .A(DP_mult_218_n486), .B(DP_mult_218_n498), .CI(
        DP_mult_218_n496), .CO(DP_mult_218_n483), .S(DP_mult_218_n484) );
  FA_X1 DP_mult_218_U303 ( .A(DP_mult_218_n484), .B(DP_mult_218_n858), .CI(
        DP_mult_218_n881), .CO(DP_mult_218_n481), .S(DP_mult_218_n482) );
  FA_X1 DP_mult_218_U301 ( .A(DP_mult_218_n742), .B(DP_mult_218_n493), .CI(
        DP_mult_218_n491), .CO(DP_mult_218_n477), .S(DP_mult_218_n478) );
  FA_X1 DP_mult_218_U300 ( .A(DP_mult_218_n478), .B(DP_mult_218_n765), .CI(
        DP_mult_218_n788), .CO(DP_mult_218_n475), .S(DP_mult_218_n476) );
  FA_X1 DP_mult_218_U299 ( .A(DP_mult_218_n476), .B(DP_mult_218_n489), .CI(
        DP_mult_218_n487), .CO(DP_mult_218_n473), .S(DP_mult_218_n474) );
  FA_X1 DP_mult_218_U298 ( .A(DP_mult_218_n474), .B(DP_mult_218_n811), .CI(
        DP_mult_218_n834), .CO(DP_mult_218_n471), .S(DP_mult_218_n472) );
  FA_X1 DP_mult_218_U297 ( .A(DP_mult_218_n472), .B(DP_mult_218_n485), .CI(
        DP_mult_218_n483), .CO(DP_mult_218_n469), .S(DP_mult_218_n470) );
  FA_X1 DP_mult_218_U296 ( .A(DP_mult_218_n880), .B(DP_mult_218_n857), .CI(
        DP_mult_218_n470), .CO(DP_mult_218_n467), .S(DP_mult_218_n468) );
  FA_X1 DP_mult_218_U295 ( .A(DP_mult_218_n479), .B(DP_mult_218_n879), .CI(
        DP_mult_218_n741), .CO(DP_mult_218_n465), .S(DP_mult_218_n466) );
  FA_X1 DP_mult_218_U294 ( .A(DP_mult_218_n764), .B(DP_mult_218_n466), .CI(
        DP_mult_218_n477), .CO(DP_mult_218_n463), .S(DP_mult_218_n464) );
  FA_X1 DP_mult_218_U293 ( .A(DP_mult_218_n475), .B(DP_mult_218_n464), .CI(
        DP_mult_218_n787), .CO(DP_mult_218_n461), .S(DP_mult_218_n462) );
  FA_X1 DP_mult_218_U292 ( .A(DP_mult_218_n810), .B(DP_mult_218_n462), .CI(
        DP_mult_218_n473), .CO(DP_mult_218_n459), .S(DP_mult_218_n460) );
  FA_X1 DP_mult_218_U291 ( .A(DP_mult_218_n471), .B(DP_mult_218_n460), .CI(
        DP_mult_218_n833), .CO(DP_mult_218_n457), .S(DP_mult_218_n458) );
  FA_X1 DP_mult_218_U290 ( .A(DP_mult_218_n856), .B(DP_mult_218_n458), .CI(
        DP_mult_218_n469), .CO(DP_mult_218_n455), .S(DP_mult_218_n456) );
  FA_X1 DP_mult_218_U288 ( .A(DP_mult_218_n454), .B(DP_mult_218_n465), .CI(
        DP_mult_218_n763), .CO(DP_mult_218_n452), .S(DP_mult_218_n453) );
  FA_X1 DP_mult_218_U287 ( .A(DP_mult_218_n453), .B(DP_mult_218_n463), .CI(
        DP_mult_218_n786), .CO(DP_mult_218_n450), .S(DP_mult_218_n451) );
  FA_X1 DP_mult_218_U286 ( .A(DP_mult_218_n451), .B(DP_mult_218_n461), .CI(
        DP_mult_218_n809), .CO(DP_mult_218_n448), .S(DP_mult_218_n449) );
  FA_X1 DP_mult_218_U285 ( .A(DP_mult_218_n449), .B(DP_mult_218_n459), .CI(
        DP_mult_218_n832), .CO(DP_mult_218_n446), .S(DP_mult_218_n447) );
  FA_X1 DP_mult_218_U284 ( .A(DP_mult_218_n447), .B(DP_mult_218_n457), .CI(
        DP_mult_218_n855), .CO(DP_mult_218_n444), .S(DP_mult_218_n445) );
  FA_X1 DP_mult_218_U282 ( .A(DP_mult_218_n740), .B(DP_mult_218_n454), .CI(
        DP_mult_218_n762), .CO(DP_mult_218_n440), .S(DP_mult_218_n441) );
  FA_X1 DP_mult_218_U281 ( .A(DP_mult_218_n441), .B(DP_mult_218_n452), .CI(
        DP_mult_218_n450), .CO(DP_mult_218_n438), .S(DP_mult_218_n439) );
  FA_X1 DP_mult_218_U280 ( .A(DP_mult_218_n439), .B(DP_mult_218_n785), .CI(
        DP_mult_218_n808), .CO(DP_mult_218_n436), .S(DP_mult_218_n437) );
  FA_X1 DP_mult_218_U279 ( .A(DP_mult_218_n437), .B(DP_mult_218_n448), .CI(
        DP_mult_218_n446), .CO(DP_mult_218_n434), .S(DP_mult_218_n435) );
  FA_X1 DP_mult_218_U278 ( .A(DP_mult_218_n854), .B(DP_mult_218_n831), .CI(
        DP_mult_218_n435), .CO(DP_mult_218_n432), .S(DP_mult_218_n433) );
  FA_X1 DP_mult_218_U277 ( .A(DP_mult_218_n442), .B(DP_mult_218_n853), .CI(
        DP_mult_218_n739), .CO(DP_mult_218_n430), .S(DP_mult_218_n431) );
  FA_X1 DP_mult_218_U276 ( .A(DP_mult_218_n440), .B(DP_mult_218_n431), .CI(
        DP_mult_218_n761), .CO(DP_mult_218_n428), .S(DP_mult_218_n429) );
  FA_X1 DP_mult_218_U275 ( .A(DP_mult_218_n784), .B(DP_mult_218_n429), .CI(
        DP_mult_218_n438), .CO(DP_mult_218_n426), .S(DP_mult_218_n427) );
  FA_X1 DP_mult_218_U274 ( .A(DP_mult_218_n436), .B(DP_mult_218_n427), .CI(
        DP_mult_218_n807), .CO(DP_mult_218_n424), .S(DP_mult_218_n425) );
  FA_X1 DP_mult_218_U273 ( .A(DP_mult_218_n830), .B(DP_mult_218_n425), .CI(
        DP_mult_218_n434), .CO(DP_mult_218_n422), .S(DP_mult_218_n423) );
  FA_X1 DP_mult_218_U271 ( .A(DP_mult_218_n421), .B(DP_mult_218_n430), .CI(
        DP_mult_218_n760), .CO(DP_mult_218_n419), .S(DP_mult_218_n420) );
  FA_X1 DP_mult_218_U270 ( .A(DP_mult_218_n420), .B(DP_mult_218_n428), .CI(
        DP_mult_218_n783), .CO(DP_mult_218_n417), .S(DP_mult_218_n418) );
  FA_X1 DP_mult_218_U269 ( .A(DP_mult_218_n418), .B(DP_mult_218_n426), .CI(
        DP_mult_218_n806), .CO(DP_mult_218_n415), .S(DP_mult_218_n416) );
  FA_X1 DP_mult_218_U268 ( .A(DP_mult_218_n416), .B(DP_mult_218_n424), .CI(
        DP_mult_218_n829), .CO(DP_mult_218_n413), .S(DP_mult_218_n414) );
  FA_X1 DP_mult_218_U266 ( .A(DP_mult_218_n738), .B(DP_mult_218_n421), .CI(
        DP_mult_218_n419), .CO(DP_mult_218_n409), .S(DP_mult_218_n410) );
  FA_X1 DP_mult_218_U265 ( .A(DP_mult_218_n410), .B(DP_mult_218_n759), .CI(
        DP_mult_218_n782), .CO(DP_mult_218_n407), .S(DP_mult_218_n408) );
  FA_X1 DP_mult_218_U264 ( .A(DP_mult_218_n408), .B(DP_mult_218_n417), .CI(
        DP_mult_218_n415), .CO(DP_mult_218_n405), .S(DP_mult_218_n406) );
  FA_X1 DP_mult_218_U263 ( .A(DP_mult_218_n828), .B(DP_mult_218_n805), .CI(
        DP_mult_218_n406), .CO(DP_mult_218_n403), .S(DP_mult_218_n404) );
  FA_X1 DP_mult_218_U262 ( .A(DP_mult_218_n411), .B(DP_mult_218_n827), .CI(
        DP_mult_218_n737), .CO(DP_mult_218_n387), .S(DP_mult_218_n402) );
  FA_X1 DP_mult_218_U261 ( .A(DP_mult_218_n758), .B(DP_mult_218_n402), .CI(
        DP_mult_218_n409), .CO(DP_mult_218_n400), .S(DP_mult_218_n401) );
  FA_X1 DP_mult_218_U260 ( .A(DP_mult_218_n407), .B(DP_mult_218_n401), .CI(
        DP_mult_218_n781), .CO(DP_mult_218_n398), .S(DP_mult_218_n399) );
  FA_X1 DP_mult_218_U259 ( .A(DP_mult_218_n804), .B(DP_mult_218_n399), .CI(
        DP_mult_218_n405), .CO(DP_mult_218_n396), .S(DP_mult_218_n397) );
  FA_X1 DP_mult_218_U257 ( .A(DP_mult_218_n395), .B(DP_mult_218_n736), .CI(
        DP_mult_218_n757), .CO(DP_mult_218_n393), .S(DP_mult_218_n394) );
  FA_X1 DP_mult_218_U256 ( .A(DP_mult_218_n394), .B(DP_mult_218_n400), .CI(
        DP_mult_218_n780), .CO(DP_mult_218_n391), .S(DP_mult_218_n392) );
  FA_X1 DP_mult_218_U255 ( .A(DP_mult_218_n392), .B(DP_mult_218_n398), .CI(
        DP_mult_218_n803), .CO(DP_mult_218_n389), .S(DP_mult_218_n390) );
  FA_X1 DP_mult_218_U253 ( .A(DP_mult_218_n735), .B(DP_mult_218_n395), .CI(
        DP_mult_218_n756), .CO(DP_mult_218_n385), .S(DP_mult_218_n386) );
  FA_X1 DP_mult_218_U252 ( .A(DP_mult_218_n386), .B(DP_mult_218_n393), .CI(
        DP_mult_218_n391), .CO(DP_mult_218_n383), .S(DP_mult_218_n384) );
  FA_X1 DP_mult_218_U251 ( .A(DP_mult_218_n802), .B(DP_mult_218_n779), .CI(
        DP_mult_218_n384), .CO(DP_mult_218_n381), .S(DP_mult_218_n382) );
  FA_X1 DP_mult_218_U250 ( .A(DP_mult_218_n387), .B(DP_mult_218_n801), .CI(
        DP_mult_218_n734), .CO(DP_mult_218_n379), .S(DP_mult_218_n380) );
  FA_X1 DP_mult_218_U249 ( .A(DP_mult_218_n385), .B(DP_mult_218_n380), .CI(
        DP_mult_218_n755), .CO(DP_mult_218_n377), .S(DP_mult_218_n378) );
  FA_X1 DP_mult_218_U248 ( .A(DP_mult_218_n778), .B(DP_mult_218_n378), .CI(
        DP_mult_218_n383), .CO(DP_mult_218_n375), .S(DP_mult_218_n376) );
  FA_X1 DP_mult_218_U246 ( .A(DP_mult_218_n374), .B(DP_mult_218_n379), .CI(
        DP_mult_218_n754), .CO(DP_mult_218_n372), .S(DP_mult_218_n373) );
  FA_X1 DP_mult_218_U245 ( .A(DP_mult_218_n373), .B(DP_mult_218_n377), .CI(
        DP_mult_218_n777), .CO(DP_mult_218_n370), .S(DP_mult_218_n371) );
  FA_X1 DP_mult_218_U243 ( .A(DP_mult_218_n733), .B(DP_mult_218_n374), .CI(
        DP_mult_218_n372), .CO(DP_mult_218_n366), .S(DP_mult_218_n367) );
  FA_X1 DP_mult_218_U242 ( .A(DP_mult_218_n776), .B(DP_mult_218_n753), .CI(
        DP_mult_218_n367), .CO(DP_mult_218_n364), .S(DP_mult_218_n365) );
  FA_X1 DP_mult_218_U241 ( .A(DP_mult_218_n368), .B(DP_mult_218_n775), .CI(
        DP_mult_218_n732), .CO(DP_mult_218_n356), .S(DP_mult_218_n363) );
  FA_X1 DP_mult_218_U240 ( .A(DP_mult_218_n752), .B(DP_mult_218_n363), .CI(
        DP_mult_218_n366), .CO(DP_mult_218_n361), .S(DP_mult_218_n362) );
  FA_X1 DP_mult_218_U238 ( .A(DP_mult_218_n360), .B(DP_mult_218_n731), .CI(
        DP_mult_218_n751), .CO(DP_mult_218_n358), .S(DP_mult_218_n359) );
  FA_X1 DP_mult_218_U236 ( .A(DP_mult_218_n730), .B(DP_mult_218_n360), .CI(
        DP_mult_218_n750), .CO(DP_mult_218_n354), .S(DP_mult_218_n355) );
  FA_X1 DP_mult_218_U235 ( .A(DP_mult_218_n356), .B(DP_mult_218_n749), .CI(
        DP_mult_218_n729), .CO(DP_mult_218_n352), .S(DP_mult_218_n353) );
  FA_X1 DP_mult_218_U204 ( .A(DP_mult_218_n908), .B(DP_mult_218_n536), .CI(
        DP_mult_218_n326), .CO(DP_mult_218_n325), .S(DP_pipe0_coeff_pipe02[0])
         );
  FA_X1 DP_mult_218_U203 ( .A(DP_mult_218_n907), .B(DP_mult_218_n522), .CI(
        DP_mult_218_n325), .CO(DP_mult_218_n324), .S(DP_pipe0_coeff_pipe02[1])
         );
  FA_X1 DP_mult_218_U202 ( .A(DP_mult_218_n508), .B(DP_mult_218_n906), .CI(
        DP_mult_218_n324), .CO(DP_mult_218_n323), .S(DP_pipe0_coeff_pipe02[2])
         );
  FA_X1 DP_mult_218_U201 ( .A(DP_mult_218_n495), .B(DP_mult_218_n507), .CI(
        DP_mult_218_n323), .CO(DP_mult_218_n322), .S(DP_pipe0_coeff_pipe02[3])
         );
  FA_X1 DP_mult_218_U200 ( .A(DP_mult_218_n482), .B(DP_mult_218_n494), .CI(
        DP_mult_218_n322), .CO(DP_mult_218_n321), .S(DP_pipe0_coeff_pipe02[4])
         );
  FA_X1 DP_mult_218_U199 ( .A(DP_mult_218_n468), .B(DP_mult_218_n481), .CI(
        DP_mult_218_n321), .CO(DP_mult_218_n320), .S(DP_pipe0_coeff_pipe02[5])
         );
  FA_X1 DP_mult_218_U198 ( .A(DP_mult_218_n456), .B(DP_mult_218_n467), .CI(
        DP_mult_218_n320), .CO(DP_mult_218_n319), .S(DP_pipe0_coeff_pipe02[6])
         );
  FA_X1 DP_mult_218_U197 ( .A(DP_mult_218_n445), .B(DP_mult_218_n455), .CI(
        DP_mult_218_n319), .CO(DP_mult_218_n318), .S(DP_pipe0_coeff_pipe02[7])
         );
  FA_X1 DP_mult_218_U196 ( .A(DP_mult_218_n433), .B(DP_mult_218_n444), .CI(
        DP_mult_218_n318), .CO(DP_mult_218_n317), .S(DP_pipe0_coeff_pipe02[8])
         );
  FA_X1 DP_mult_218_U195 ( .A(DP_mult_218_n423), .B(DP_mult_218_n432), .CI(
        DP_mult_218_n317), .CO(DP_mult_218_n316), .S(DP_pipe0_coeff_pipe02[9])
         );
  FA_X1 DP_mult_218_U194 ( .A(DP_mult_218_n414), .B(DP_mult_218_n422), .CI(
        DP_mult_218_n316), .CO(DP_mult_218_n315), .S(DP_pipe0_coeff_pipe02[10]) );
  FA_X1 DP_mult_218_U193 ( .A(DP_mult_218_n404), .B(DP_mult_218_n413), .CI(
        DP_mult_218_n315), .CO(DP_mult_218_n314), .S(DP_pipe0_coeff_pipe02[11]) );
  FA_X1 DP_mult_218_U192 ( .A(DP_mult_218_n397), .B(DP_mult_218_n403), .CI(
        DP_mult_218_n314), .CO(DP_mult_218_n313), .S(DP_pipe0_coeff_pipe02[12]) );
  FA_X1 DP_mult_218_U191 ( .A(DP_mult_218_n390), .B(DP_mult_218_n396), .CI(
        DP_mult_218_n313), .CO(DP_mult_218_n312), .S(DP_pipe0_coeff_pipe02[13]) );
  FA_X1 DP_mult_218_U190 ( .A(DP_mult_218_n382), .B(DP_mult_218_n389), .CI(
        DP_mult_218_n312), .CO(DP_mult_218_n311), .S(DP_pipe0_coeff_pipe02[14]) );
  FA_X1 DP_mult_218_U189 ( .A(DP_mult_218_n376), .B(DP_mult_218_n381), .CI(
        DP_mult_218_n311), .CO(DP_mult_218_n310), .S(DP_pipe0_coeff_pipe02[15]) );
  FA_X1 DP_mult_218_U188 ( .A(DP_mult_218_n371), .B(DP_mult_218_n375), .CI(
        DP_mult_218_n310), .CO(DP_mult_218_n309), .S(DP_pipe0_coeff_pipe02[16]) );
  FA_X1 DP_mult_218_U187 ( .A(DP_mult_218_n365), .B(DP_mult_218_n370), .CI(
        DP_mult_218_n309), .CO(DP_mult_218_n308), .S(DP_pipe0_coeff_pipe02[17]) );
  FA_X1 DP_mult_218_U186 ( .A(DP_mult_218_n362), .B(DP_mult_218_n364), .CI(
        DP_mult_218_n308), .CO(DP_mult_218_n307), .S(DP_pipe0_coeff_pipe02[18]) );
  FA_X1 DP_mult_218_U185 ( .A(DP_mult_218_n359), .B(DP_mult_218_n361), .CI(
        DP_mult_218_n307), .CO(DP_mult_218_n306), .S(DP_pipe0_coeff_pipe02[19]) );
  FA_X1 DP_mult_218_U184 ( .A(DP_mult_218_n355), .B(DP_mult_218_n358), .CI(
        DP_mult_218_n306), .CO(DP_mult_218_n305), .S(DP_pipe0_coeff_pipe02[20]) );
  FA_X1 DP_mult_218_U183 ( .A(DP_mult_218_n353), .B(DP_mult_218_n354), .CI(
        DP_mult_218_n305), .CO(DP_mult_218_n304), .S(DP_pipe0_coeff_pipe02[21]) );
  FA_X1 DP_mult_218_U182 ( .A(DP_mult_218_n351), .B(DP_mult_218_n352), .CI(
        DP_mult_218_n304), .CO(DP_mult_218_n303), .S(DP_pipe0_coeff_pipe02[22]) );
  INV_X1 DP_mult_217_U1959 ( .A(DP_coeff_pipe01[1]), .ZN(DP_mult_217_n2159) );
  NOR2_X1 DP_mult_217_U1958 ( .A1(DP_mult_217_n2159), .A2(DP_coeff_pipe01[0]), 
        .ZN(DP_mult_217_n1636) );
  INV_X1 DP_mult_217_U1957 ( .A(DP_coeff_pipe01[2]), .ZN(DP_mult_217_n1742) );
  XNOR2_X1 DP_mult_217_U1956 ( .A(DP_coeff_pipe01[1]), .B(DP_mult_217_n1742), 
        .ZN(DP_mult_217_n2157) );
  AOI221_X1 DP_mult_217_U1955 ( .B1(DP_pipe01[1]), .B2(DP_mult_217_n1563), 
        .C1(DP_mult_217_n1396), .C2(DP_mult_217_n1554), .A(DP_mult_217_n1742), 
        .ZN(DP_mult_217_n2160) );
  INV_X1 DP_mult_217_U1954 ( .A(DP_coeff_pipe01[0]), .ZN(DP_mult_217_n2158) );
  INV_X1 DP_mult_217_U1953 ( .A(DP_pipe01[2]), .ZN(DP_mult_217_n1661) );
  INV_X1 DP_mult_217_U1952 ( .A(DP_mult_217_n1397), .ZN(DP_mult_217_n1650) );
  OAI22_X1 DP_mult_217_U1951 ( .A1(DP_mult_217_n1542), .A2(DP_mult_217_n1661), 
        .B1(DP_mult_217_n1564), .B2(DP_mult_217_n1650), .ZN(DP_mult_217_n2162)
         );
  AOI211_X1 DP_mult_217_U1950 ( .C1(DP_pipe01[1]), .C2(DP_mult_217_n1561), .A(
        DP_mult_217_n2162), .B(DP_pipe01[0]), .ZN(DP_mult_217_n2161) );
  AND2_X1 DP_mult_217_U1949 ( .A1(DP_mult_217_n2160), .A2(DP_mult_217_n2161), 
        .ZN(DP_mult_217_n2153) );
  INV_X1 DP_mult_217_U1948 ( .A(DP_mult_217_n1395), .ZN(DP_mult_217_n1657) );
  INV_X1 DP_mult_217_U1947 ( .A(DP_pipe01[1]), .ZN(DP_mult_217_n1649) );
  OAI22_X1 DP_mult_217_U1946 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1657), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1649), .ZN(DP_mult_217_n2156)
         );
  AOI221_X1 DP_mult_217_U1945 ( .B1(DP_pipe01[3]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[2]), .C2(DP_mult_217_n1563), .A(DP_mult_217_n2156), .ZN(
        DP_mult_217_n2155) );
  XNOR2_X1 DP_mult_217_U1944 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2155), 
        .ZN(DP_mult_217_n2154) );
  AOI222_X1 DP_mult_217_U1943 ( .A1(DP_mult_217_n2153), .A2(DP_mult_217_n2154), 
        .B1(DP_mult_217_n2153), .B2(DP_mult_217_n688), .C1(DP_mult_217_n688), 
        .C2(DP_mult_217_n2154), .ZN(DP_mult_217_n2148) );
  INV_X1 DP_mult_217_U1942 ( .A(DP_mult_217_n1394), .ZN(DP_mult_217_n1660) );
  OAI22_X1 DP_mult_217_U1941 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1660), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1661), .ZN(DP_mult_217_n2152)
         );
  AOI221_X1 DP_mult_217_U1940 ( .B1(DP_pipe01[4]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[3]), .C2(DP_mult_217_n1563), .A(DP_mult_217_n2152), .ZN(
        DP_mult_217_n2151) );
  XNOR2_X1 DP_mult_217_U1939 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2151), 
        .ZN(DP_mult_217_n2149) );
  INV_X1 DP_mult_217_U1938 ( .A(DP_mult_217_n686), .ZN(DP_mult_217_n2150) );
  OAI222_X1 DP_mult_217_U1937 ( .A1(DP_mult_217_n2148), .A2(DP_mult_217_n2149), 
        .B1(DP_mult_217_n2148), .B2(DP_mult_217_n2150), .C1(DP_mult_217_n2150), 
        .C2(DP_mult_217_n2149), .ZN(DP_mult_217_n2144) );
  INV_X1 DP_mult_217_U1936 ( .A(DP_mult_217_n1393), .ZN(DP_mult_217_n1664) );
  INV_X1 DP_mult_217_U1935 ( .A(DP_pipe01[3]), .ZN(DP_mult_217_n1665) );
  OAI22_X1 DP_mult_217_U1934 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1664), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1665), .ZN(DP_mult_217_n2147)
         );
  AOI221_X1 DP_mult_217_U1933 ( .B1(DP_pipe01[5]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[4]), .C2(DP_mult_217_n1563), .A(DP_mult_217_n2147), .ZN(
        DP_mult_217_n2146) );
  XNOR2_X1 DP_mult_217_U1932 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2146), 
        .ZN(DP_mult_217_n2145) );
  AOI222_X1 DP_mult_217_U1931 ( .A1(DP_mult_217_n2144), .A2(DP_mult_217_n2145), 
        .B1(DP_mult_217_n2144), .B2(DP_mult_217_n684), .C1(DP_mult_217_n684), 
        .C2(DP_mult_217_n2145), .ZN(DP_mult_217_n2139) );
  INV_X1 DP_mult_217_U1930 ( .A(DP_mult_217_n1392), .ZN(DP_mult_217_n1668) );
  INV_X1 DP_mult_217_U1929 ( .A(DP_pipe01[4]), .ZN(DP_mult_217_n1669) );
  OAI22_X1 DP_mult_217_U1928 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1668), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1669), .ZN(DP_mult_217_n2143)
         );
  AOI221_X1 DP_mult_217_U1927 ( .B1(DP_pipe01[6]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[5]), .C2(DP_mult_217_n1563), .A(DP_mult_217_n2143), .ZN(
        DP_mult_217_n2142) );
  XNOR2_X1 DP_mult_217_U1926 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2142), 
        .ZN(DP_mult_217_n2140) );
  INV_X1 DP_mult_217_U1925 ( .A(DP_mult_217_n680), .ZN(DP_mult_217_n2141) );
  OAI222_X1 DP_mult_217_U1924 ( .A1(DP_mult_217_n2139), .A2(DP_mult_217_n2140), 
        .B1(DP_mult_217_n2139), .B2(DP_mult_217_n2141), .C1(DP_mult_217_n2141), 
        .C2(DP_mult_217_n2140), .ZN(DP_mult_217_n2135) );
  INV_X1 DP_mult_217_U1923 ( .A(DP_mult_217_n1391), .ZN(DP_mult_217_n1672) );
  INV_X1 DP_mult_217_U1922 ( .A(DP_pipe01[5]), .ZN(DP_mult_217_n1673) );
  OAI22_X1 DP_mult_217_U1921 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1672), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1673), .ZN(DP_mult_217_n2138)
         );
  AOI221_X1 DP_mult_217_U1920 ( .B1(DP_pipe01[7]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[6]), .C2(DP_mult_217_n1563), .A(DP_mult_217_n2138), .ZN(
        DP_mult_217_n2137) );
  XNOR2_X1 DP_mult_217_U1919 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2137), 
        .ZN(DP_mult_217_n2136) );
  AOI222_X1 DP_mult_217_U1918 ( .A1(DP_mult_217_n2135), .A2(DP_mult_217_n2136), 
        .B1(DP_mult_217_n2135), .B2(DP_mult_217_n676), .C1(DP_mult_217_n676), 
        .C2(DP_mult_217_n2136), .ZN(DP_mult_217_n2130) );
  INV_X1 DP_mult_217_U1917 ( .A(DP_mult_217_n1390), .ZN(DP_mult_217_n1676) );
  INV_X1 DP_mult_217_U1916 ( .A(DP_pipe01[6]), .ZN(DP_mult_217_n1677) );
  OAI22_X1 DP_mult_217_U1915 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1676), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1677), .ZN(DP_mult_217_n2134)
         );
  AOI221_X1 DP_mult_217_U1914 ( .B1(DP_pipe01[8]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[7]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2134), .ZN(
        DP_mult_217_n2133) );
  XNOR2_X1 DP_mult_217_U1913 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2133), 
        .ZN(DP_mult_217_n2131) );
  INV_X1 DP_mult_217_U1912 ( .A(DP_mult_217_n672), .ZN(DP_mult_217_n2132) );
  OAI222_X1 DP_mult_217_U1911 ( .A1(DP_mult_217_n2130), .A2(DP_mult_217_n2131), 
        .B1(DP_mult_217_n2130), .B2(DP_mult_217_n2132), .C1(DP_mult_217_n2132), 
        .C2(DP_mult_217_n2131), .ZN(DP_mult_217_n2126) );
  INV_X1 DP_mult_217_U1910 ( .A(DP_mult_217_n1389), .ZN(DP_mult_217_n1680) );
  INV_X1 DP_mult_217_U1909 ( .A(DP_pipe01[7]), .ZN(DP_mult_217_n1681) );
  OAI22_X1 DP_mult_217_U1908 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1680), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1681), .ZN(DP_mult_217_n2129)
         );
  AOI221_X1 DP_mult_217_U1907 ( .B1(DP_pipe01[9]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[8]), .C2(DP_mult_217_n1563), .A(DP_mult_217_n2129), .ZN(
        DP_mult_217_n2128) );
  XNOR2_X1 DP_mult_217_U1906 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2128), 
        .ZN(DP_mult_217_n2127) );
  AOI222_X1 DP_mult_217_U1905 ( .A1(DP_mult_217_n2126), .A2(DP_mult_217_n2127), 
        .B1(DP_mult_217_n2126), .B2(DP_mult_217_n666), .C1(DP_mult_217_n666), 
        .C2(DP_mult_217_n2127), .ZN(DP_mult_217_n2121) );
  INV_X1 DP_mult_217_U1904 ( .A(DP_mult_217_n1388), .ZN(DP_mult_217_n1684) );
  INV_X1 DP_mult_217_U1903 ( .A(DP_pipe01[8]), .ZN(DP_mult_217_n1685) );
  OAI22_X1 DP_mult_217_U1902 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1684), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1685), .ZN(DP_mult_217_n2125)
         );
  AOI221_X1 DP_mult_217_U1901 ( .B1(DP_pipe01[10]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[9]), .C2(DP_mult_217_n1563), .A(DP_mult_217_n2125), .ZN(
        DP_mult_217_n2124) );
  XNOR2_X1 DP_mult_217_U1900 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2124), 
        .ZN(DP_mult_217_n2122) );
  INV_X1 DP_mult_217_U1899 ( .A(DP_mult_217_n660), .ZN(DP_mult_217_n2123) );
  OAI222_X1 DP_mult_217_U1898 ( .A1(DP_mult_217_n2121), .A2(DP_mult_217_n2122), 
        .B1(DP_mult_217_n2121), .B2(DP_mult_217_n2123), .C1(DP_mult_217_n2123), 
        .C2(DP_mult_217_n2122), .ZN(DP_mult_217_n2117) );
  INV_X1 DP_mult_217_U1897 ( .A(DP_mult_217_n1387), .ZN(DP_mult_217_n1688) );
  INV_X1 DP_mult_217_U1896 ( .A(DP_pipe01[9]), .ZN(DP_mult_217_n1689) );
  OAI22_X1 DP_mult_217_U1895 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1688), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1689), .ZN(DP_mult_217_n2120)
         );
  AOI221_X1 DP_mult_217_U1894 ( .B1(DP_pipe01[11]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[10]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2120), 
        .ZN(DP_mult_217_n2119) );
  XNOR2_X1 DP_mult_217_U1893 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2119), 
        .ZN(DP_mult_217_n2118) );
  AOI222_X1 DP_mult_217_U1892 ( .A1(DP_mult_217_n2117), .A2(DP_mult_217_n2118), 
        .B1(DP_mult_217_n2117), .B2(DP_mult_217_n654), .C1(DP_mult_217_n654), 
        .C2(DP_mult_217_n2118), .ZN(DP_mult_217_n2112) );
  INV_X1 DP_mult_217_U1891 ( .A(DP_mult_217_n1386), .ZN(DP_mult_217_n1692) );
  INV_X1 DP_mult_217_U1890 ( .A(DP_pipe01[10]), .ZN(DP_mult_217_n1693) );
  OAI22_X1 DP_mult_217_U1889 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1692), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1693), .ZN(DP_mult_217_n2116)
         );
  AOI221_X1 DP_mult_217_U1888 ( .B1(DP_pipe01[12]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[11]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2116), 
        .ZN(DP_mult_217_n2115) );
  XNOR2_X1 DP_mult_217_U1887 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2115), 
        .ZN(DP_mult_217_n2113) );
  INV_X1 DP_mult_217_U1886 ( .A(DP_mult_217_n646), .ZN(DP_mult_217_n2114) );
  OAI222_X1 DP_mult_217_U1885 ( .A1(DP_mult_217_n2112), .A2(DP_mult_217_n2113), 
        .B1(DP_mult_217_n2112), .B2(DP_mult_217_n2114), .C1(DP_mult_217_n2114), 
        .C2(DP_mult_217_n2113), .ZN(DP_mult_217_n2108) );
  INV_X1 DP_mult_217_U1884 ( .A(DP_mult_217_n1385), .ZN(DP_mult_217_n1696) );
  INV_X1 DP_mult_217_U1883 ( .A(DP_pipe01[11]), .ZN(DP_mult_217_n1697) );
  OAI22_X1 DP_mult_217_U1882 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1696), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1697), .ZN(DP_mult_217_n2111)
         );
  AOI221_X1 DP_mult_217_U1881 ( .B1(DP_pipe01[13]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[12]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2111), 
        .ZN(DP_mult_217_n2110) );
  XNOR2_X1 DP_mult_217_U1880 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2110), 
        .ZN(DP_mult_217_n2109) );
  AOI222_X1 DP_mult_217_U1879 ( .A1(DP_mult_217_n2108), .A2(DP_mult_217_n2109), 
        .B1(DP_mult_217_n2108), .B2(DP_mult_217_n638), .C1(DP_mult_217_n638), 
        .C2(DP_mult_217_n2109), .ZN(DP_mult_217_n2103) );
  INV_X1 DP_mult_217_U1878 ( .A(DP_mult_217_n1384), .ZN(DP_mult_217_n1700) );
  INV_X1 DP_mult_217_U1877 ( .A(DP_pipe01[12]), .ZN(DP_mult_217_n1701) );
  OAI22_X1 DP_mult_217_U1876 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1700), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1701), .ZN(DP_mult_217_n2107)
         );
  AOI221_X1 DP_mult_217_U1875 ( .B1(DP_pipe01[14]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[13]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2107), 
        .ZN(DP_mult_217_n2106) );
  XNOR2_X1 DP_mult_217_U1874 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2106), 
        .ZN(DP_mult_217_n2104) );
  INV_X1 DP_mult_217_U1873 ( .A(DP_mult_217_n630), .ZN(DP_mult_217_n2105) );
  OAI222_X1 DP_mult_217_U1872 ( .A1(DP_mult_217_n2103), .A2(DP_mult_217_n2104), 
        .B1(DP_mult_217_n2103), .B2(DP_mult_217_n2105), .C1(DP_mult_217_n2105), 
        .C2(DP_mult_217_n2104), .ZN(DP_mult_217_n2099) );
  INV_X1 DP_mult_217_U1871 ( .A(DP_mult_217_n1383), .ZN(DP_mult_217_n1704) );
  INV_X1 DP_mult_217_U1870 ( .A(DP_pipe01[13]), .ZN(DP_mult_217_n1705) );
  OAI22_X1 DP_mult_217_U1869 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1704), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1705), .ZN(DP_mult_217_n2102)
         );
  AOI221_X1 DP_mult_217_U1868 ( .B1(DP_pipe01[15]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[14]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2102), 
        .ZN(DP_mult_217_n2101) );
  XNOR2_X1 DP_mult_217_U1867 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2101), 
        .ZN(DP_mult_217_n2100) );
  AOI222_X1 DP_mult_217_U1866 ( .A1(DP_mult_217_n2099), .A2(DP_mult_217_n2100), 
        .B1(DP_mult_217_n2099), .B2(DP_mult_217_n620), .C1(DP_mult_217_n620), 
        .C2(DP_mult_217_n2100), .ZN(DP_mult_217_n2094) );
  INV_X1 DP_mult_217_U1865 ( .A(DP_mult_217_n1382), .ZN(DP_mult_217_n1708) );
  INV_X1 DP_mult_217_U1864 ( .A(DP_pipe01[14]), .ZN(DP_mult_217_n1709) );
  OAI22_X1 DP_mult_217_U1863 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1708), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1709), .ZN(DP_mult_217_n2098)
         );
  AOI221_X1 DP_mult_217_U1862 ( .B1(DP_pipe01[16]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[15]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2098), 
        .ZN(DP_mult_217_n2097) );
  XNOR2_X1 DP_mult_217_U1861 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2097), 
        .ZN(DP_mult_217_n2095) );
  INV_X1 DP_mult_217_U1860 ( .A(DP_mult_217_n610), .ZN(DP_mult_217_n2096) );
  OAI222_X1 DP_mult_217_U1859 ( .A1(DP_mult_217_n2094), .A2(DP_mult_217_n2095), 
        .B1(DP_mult_217_n2094), .B2(DP_mult_217_n2096), .C1(DP_mult_217_n2096), 
        .C2(DP_mult_217_n2095), .ZN(DP_mult_217_n2090) );
  INV_X1 DP_mult_217_U1858 ( .A(DP_mult_217_n1381), .ZN(DP_mult_217_n1712) );
  INV_X1 DP_mult_217_U1857 ( .A(DP_pipe01[15]), .ZN(DP_mult_217_n1713) );
  OAI22_X1 DP_mult_217_U1856 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1712), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1713), .ZN(DP_mult_217_n2093)
         );
  AOI221_X1 DP_mult_217_U1855 ( .B1(DP_pipe01[17]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[16]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2093), 
        .ZN(DP_mult_217_n2092) );
  XNOR2_X1 DP_mult_217_U1854 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2092), 
        .ZN(DP_mult_217_n2091) );
  AOI222_X1 DP_mult_217_U1853 ( .A1(DP_mult_217_n2090), .A2(DP_mult_217_n2091), 
        .B1(DP_mult_217_n2090), .B2(DP_mult_217_n600), .C1(DP_mult_217_n600), 
        .C2(DP_mult_217_n2091), .ZN(DP_mult_217_n2085) );
  INV_X1 DP_mult_217_U1852 ( .A(DP_mult_217_n1380), .ZN(DP_mult_217_n1716) );
  INV_X1 DP_mult_217_U1851 ( .A(DP_pipe01[16]), .ZN(DP_mult_217_n1717) );
  OAI22_X1 DP_mult_217_U1850 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1716), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1717), .ZN(DP_mult_217_n2089)
         );
  AOI221_X1 DP_mult_217_U1849 ( .B1(DP_pipe01[18]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[17]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2089), 
        .ZN(DP_mult_217_n2088) );
  XNOR2_X1 DP_mult_217_U1848 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2088), 
        .ZN(DP_mult_217_n2086) );
  INV_X1 DP_mult_217_U1847 ( .A(DP_mult_217_n588), .ZN(DP_mult_217_n2087) );
  OAI222_X1 DP_mult_217_U1846 ( .A1(DP_mult_217_n2085), .A2(DP_mult_217_n2086), 
        .B1(DP_mult_217_n2085), .B2(DP_mult_217_n2087), .C1(DP_mult_217_n2087), 
        .C2(DP_mult_217_n2086), .ZN(DP_mult_217_n2081) );
  INV_X1 DP_mult_217_U1845 ( .A(DP_mult_217_n1379), .ZN(DP_mult_217_n1720) );
  INV_X1 DP_mult_217_U1844 ( .A(DP_pipe01[17]), .ZN(DP_mult_217_n1721) );
  OAI22_X1 DP_mult_217_U1843 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1720), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1721), .ZN(DP_mult_217_n2084)
         );
  AOI221_X1 DP_mult_217_U1842 ( .B1(DP_pipe01[19]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[18]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2084), 
        .ZN(DP_mult_217_n2083) );
  XNOR2_X1 DP_mult_217_U1841 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2083), 
        .ZN(DP_mult_217_n2082) );
  AOI222_X1 DP_mult_217_U1840 ( .A1(DP_mult_217_n2081), .A2(DP_mult_217_n2082), 
        .B1(DP_mult_217_n2081), .B2(DP_mult_217_n576), .C1(DP_mult_217_n576), 
        .C2(DP_mult_217_n2082), .ZN(DP_mult_217_n2080) );
  INV_X1 DP_mult_217_U1839 ( .A(DP_mult_217_n2080), .ZN(DP_mult_217_n2076) );
  INV_X1 DP_mult_217_U1838 ( .A(DP_mult_217_n1378), .ZN(DP_mult_217_n1724) );
  INV_X1 DP_mult_217_U1837 ( .A(DP_pipe01[18]), .ZN(DP_mult_217_n1725) );
  OAI22_X1 DP_mult_217_U1836 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1724), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1725), .ZN(DP_mult_217_n2079)
         );
  AOI221_X1 DP_mult_217_U1835 ( .B1(DP_pipe01[20]), .B2(DP_mult_217_n1561), 
        .C1(DP_pipe01[19]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2079), 
        .ZN(DP_mult_217_n2078) );
  XNOR2_X1 DP_mult_217_U1834 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n2078), 
        .ZN(DP_mult_217_n2077) );
  AOI222_X1 DP_mult_217_U1833 ( .A1(DP_mult_217_n2076), .A2(DP_mult_217_n2077), 
        .B1(DP_mult_217_n2076), .B2(DP_mult_217_n564), .C1(DP_mult_217_n564), 
        .C2(DP_mult_217_n2077), .ZN(DP_mult_217_n2071) );
  INV_X1 DP_mult_217_U1832 ( .A(DP_mult_217_n1377), .ZN(DP_mult_217_n1728) );
  INV_X1 DP_mult_217_U1831 ( .A(DP_pipe01[19]), .ZN(DP_mult_217_n1729) );
  OAI22_X1 DP_mult_217_U1830 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1728), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1729), .ZN(DP_mult_217_n2075)
         );
  AOI221_X1 DP_mult_217_U1829 ( .B1(DP_mult_217_n1561), .B2(DP_pipe01[21]), 
        .C1(DP_pipe01[20]), .C2(DP_mult_217_n1562), .A(DP_mult_217_n2075), 
        .ZN(DP_mult_217_n2074) );
  XNOR2_X1 DP_mult_217_U1828 ( .A(DP_mult_217_n1742), .B(DP_mult_217_n2074), 
        .ZN(DP_mult_217_n2072) );
  INV_X1 DP_mult_217_U1827 ( .A(DP_mult_217_n550), .ZN(DP_mult_217_n2073) );
  OAI222_X1 DP_mult_217_U1826 ( .A1(DP_mult_217_n2071), .A2(DP_mult_217_n2072), 
        .B1(DP_mult_217_n2071), .B2(DP_mult_217_n2073), .C1(DP_mult_217_n2073), 
        .C2(DP_mult_217_n2072), .ZN(DP_mult_217_n326) );
  XNOR2_X1 DP_mult_217_U1825 ( .A(DP_coeff_pipe01[21]), .B(DP_mult_217_n1608), 
        .ZN(DP_mult_217_n2067) );
  INV_X1 DP_mult_217_U1824 ( .A(DP_mult_217_n2067), .ZN(DP_mult_217_n2070) );
  XNOR2_X1 DP_mult_217_U1823 ( .A(DP_coeff_pipe01[21]), .B(DP_coeff_pipe01[22]), .ZN(DP_mult_217_n2069) );
  XNOR2_X1 DP_mult_217_U1822 ( .A(DP_coeff_pipe01[22]), .B(DP_mult_217_n1611), 
        .ZN(DP_mult_217_n2068) );
  NAND3_X1 DP_mult_217_U1821 ( .A1(DP_mult_217_n2067), .A2(DP_mult_217_n2068), 
        .A3(DP_mult_217_n2069), .ZN(DP_mult_217_n1629) );
  INV_X1 DP_mult_217_U1820 ( .A(DP_pipe01[21]), .ZN(DP_mult_217_n1643) );
  OAI22_X1 DP_mult_217_U1819 ( .A1(DP_mult_217_n1544), .A2(DP_mult_217_n1619), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1643), .ZN(DP_mult_217_n2066)
         );
  AOI221_X1 DP_mult_217_U1818 ( .B1(DP_pipe01[22]), .B2(DP_mult_217_n1560), 
        .C1(DP_mult_217_n1375), .C2(DP_mult_217_n1553), .A(DP_mult_217_n2066), 
        .ZN(DP_mult_217_n2065) );
  XOR2_X1 DP_mult_217_U1817 ( .A(DP_mult_217_n1611), .B(DP_mult_217_n2065), 
        .Z(DP_mult_217_n1627) );
  INV_X1 DP_mult_217_U1816 ( .A(DP_mult_217_n1627), .ZN(DP_mult_217_n351) );
  INV_X1 DP_mult_217_U1815 ( .A(DP_mult_217_n356), .ZN(DP_mult_217_n360) );
  OAI22_X1 DP_mult_217_U1814 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1712), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1713), .ZN(DP_mult_217_n2064)
         );
  AOI221_X1 DP_mult_217_U1813 ( .B1(DP_pipe01[17]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[16]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2064), 
        .ZN(DP_mult_217_n2063) );
  XOR2_X1 DP_mult_217_U1812 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2063), 
        .Z(DP_mult_217_n374) );
  INV_X1 DP_mult_217_U1811 ( .A(DP_mult_217_n374), .ZN(DP_mult_217_n368) );
  INV_X1 DP_mult_217_U1810 ( .A(DP_mult_217_n387), .ZN(DP_mult_217_n395) );
  OAI22_X1 DP_mult_217_U1809 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1688), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1689), .ZN(DP_mult_217_n2062)
         );
  AOI221_X1 DP_mult_217_U1808 ( .B1(DP_pipe01[11]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[10]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2062), 
        .ZN(DP_mult_217_n2061) );
  XOR2_X1 DP_mult_217_U1807 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2061), 
        .Z(DP_mult_217_n421) );
  INV_X1 DP_mult_217_U1806 ( .A(DP_mult_217_n421), .ZN(DP_mult_217_n411) );
  OAI22_X1 DP_mult_217_U1805 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1676), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1677), .ZN(DP_mult_217_n2060)
         );
  AOI221_X1 DP_mult_217_U1804 ( .B1(DP_pipe01[8]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[7]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2060), .ZN(
        DP_mult_217_n2059) );
  XOR2_X1 DP_mult_217_U1803 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2059), 
        .Z(DP_mult_217_n454) );
  INV_X1 DP_mult_217_U1802 ( .A(DP_mult_217_n454), .ZN(DP_mult_217_n442) );
  OAI21_X1 DP_mult_217_U1801 ( .B1(DP_mult_217_n1561), .B2(DP_mult_217_n1563), 
        .A(DP_mult_217_n1615), .ZN(DP_mult_217_n2058) );
  OAI221_X1 DP_mult_217_U1800 ( .B1(DP_mult_217_n1619), .B2(DP_mult_217_n1639), 
        .C1(DP_mult_217_n1620), .C2(DP_mult_217_n1564), .A(DP_mult_217_n2058), 
        .ZN(DP_mult_217_n2057) );
  XOR2_X1 DP_mult_217_U1799 ( .A(DP_mult_217_n2057), .B(DP_mult_217_n1742), 
        .Z(DP_mult_217_n2056) );
  NOR2_X1 DP_mult_217_U1798 ( .A1(DP_mult_217_n2056), .A2(DP_mult_217_n519), 
        .ZN(DP_mult_217_n493) );
  INV_X1 DP_mult_217_U1797 ( .A(DP_mult_217_n493), .ZN(DP_mult_217_n479) );
  XNOR2_X1 DP_mult_217_U1796 ( .A(DP_mult_217_n519), .B(DP_mult_217_n2056), 
        .ZN(DP_mult_217_n506) );
  INV_X1 DP_mult_217_U1795 ( .A(DP_pipe01[20]), .ZN(DP_mult_217_n1640) );
  OAI22_X1 DP_mult_217_U1794 ( .A1(DP_mult_217_n1556), .A2(DP_mult_217_n1640), 
        .B1(DP_mult_217_n1550), .B2(DP_mult_217_n1643), .ZN(DP_mult_217_n2055)
         );
  AOI221_X1 DP_mult_217_U1793 ( .B1(DP_pipe01[22]), .B2(DP_mult_217_n1559), 
        .C1(DP_mult_217_n1376), .C2(DP_mult_217_n1553), .A(DP_mult_217_n2055), 
        .ZN(DP_mult_217_n2054) );
  XNOR2_X1 DP_mult_217_U1792 ( .A(DP_coeff_pipe01[23]), .B(DP_mult_217_n2054), 
        .ZN(DP_mult_217_n729) );
  OAI22_X1 DP_mult_217_U1791 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1728), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1729), .ZN(DP_mult_217_n2053)
         );
  AOI221_X1 DP_mult_217_U1790 ( .B1(DP_pipe01[21]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[20]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2053), 
        .ZN(DP_mult_217_n2052) );
  XNOR2_X1 DP_mult_217_U1789 ( .A(DP_coeff_pipe01[23]), .B(DP_mult_217_n2052), 
        .ZN(DP_mult_217_n730) );
  OAI22_X1 DP_mult_217_U1788 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1724), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1725), .ZN(DP_mult_217_n2051)
         );
  AOI221_X1 DP_mult_217_U1787 ( .B1(DP_pipe01[20]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[19]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2051), 
        .ZN(DP_mult_217_n2050) );
  XNOR2_X1 DP_mult_217_U1786 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2050), 
        .ZN(DP_mult_217_n731) );
  OAI22_X1 DP_mult_217_U1785 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1720), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1721), .ZN(DP_mult_217_n2049)
         );
  AOI221_X1 DP_mult_217_U1784 ( .B1(DP_pipe01[19]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[18]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2049), 
        .ZN(DP_mult_217_n2048) );
  XNOR2_X1 DP_mult_217_U1783 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2048), 
        .ZN(DP_mult_217_n732) );
  OAI22_X1 DP_mult_217_U1782 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1716), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1717), .ZN(DP_mult_217_n2047)
         );
  AOI221_X1 DP_mult_217_U1781 ( .B1(DP_pipe01[18]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[17]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2047), 
        .ZN(DP_mult_217_n2046) );
  XNOR2_X1 DP_mult_217_U1780 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2046), 
        .ZN(DP_mult_217_n733) );
  OAI22_X1 DP_mult_217_U1779 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1708), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1709), .ZN(DP_mult_217_n2045)
         );
  AOI221_X1 DP_mult_217_U1778 ( .B1(DP_pipe01[16]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[15]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2045), 
        .ZN(DP_mult_217_n2044) );
  XNOR2_X1 DP_mult_217_U1777 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2044), 
        .ZN(DP_mult_217_n734) );
  OAI22_X1 DP_mult_217_U1776 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1704), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1705), .ZN(DP_mult_217_n2043)
         );
  AOI221_X1 DP_mult_217_U1775 ( .B1(DP_pipe01[15]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[14]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2043), 
        .ZN(DP_mult_217_n2042) );
  XNOR2_X1 DP_mult_217_U1774 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2042), 
        .ZN(DP_mult_217_n735) );
  OAI22_X1 DP_mult_217_U1773 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1700), 
        .B1(DP_mult_217_n1556), .B2(DP_mult_217_n1701), .ZN(DP_mult_217_n2041)
         );
  AOI221_X1 DP_mult_217_U1772 ( .B1(DP_pipe01[14]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[13]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2041), 
        .ZN(DP_mult_217_n2040) );
  XNOR2_X1 DP_mult_217_U1771 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2040), 
        .ZN(DP_mult_217_n736) );
  OAI22_X1 DP_mult_217_U1770 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1696), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1697), .ZN(DP_mult_217_n2039)
         );
  AOI221_X1 DP_mult_217_U1769 ( .B1(DP_pipe01[13]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[12]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2039), 
        .ZN(DP_mult_217_n2038) );
  XNOR2_X1 DP_mult_217_U1768 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2038), 
        .ZN(DP_mult_217_n737) );
  OAI22_X1 DP_mult_217_U1767 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1692), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1693), .ZN(DP_mult_217_n2037)
         );
  AOI221_X1 DP_mult_217_U1766 ( .B1(DP_pipe01[12]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[11]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2037), 
        .ZN(DP_mult_217_n2036) );
  XNOR2_X1 DP_mult_217_U1765 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2036), 
        .ZN(DP_mult_217_n738) );
  OAI22_X1 DP_mult_217_U1764 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1684), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1685), .ZN(DP_mult_217_n2035)
         );
  AOI221_X1 DP_mult_217_U1763 ( .B1(DP_pipe01[10]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[9]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2035), .ZN(
        DP_mult_217_n2034) );
  XNOR2_X1 DP_mult_217_U1762 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2034), 
        .ZN(DP_mult_217_n739) );
  OAI22_X1 DP_mult_217_U1761 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1680), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1681), .ZN(DP_mult_217_n2033)
         );
  AOI221_X1 DP_mult_217_U1760 ( .B1(DP_pipe01[9]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[8]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2033), .ZN(
        DP_mult_217_n2032) );
  XNOR2_X1 DP_mult_217_U1759 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2032), 
        .ZN(DP_mult_217_n740) );
  OAI22_X1 DP_mult_217_U1758 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1672), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1673), .ZN(DP_mult_217_n2031)
         );
  AOI221_X1 DP_mult_217_U1757 ( .B1(DP_pipe01[7]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[6]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2031), .ZN(
        DP_mult_217_n2030) );
  XNOR2_X1 DP_mult_217_U1756 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2030), 
        .ZN(DP_mult_217_n741) );
  OAI22_X1 DP_mult_217_U1755 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1668), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1669), .ZN(DP_mult_217_n2029)
         );
  AOI221_X1 DP_mult_217_U1754 ( .B1(DP_pipe01[6]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[5]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2029), .ZN(
        DP_mult_217_n2028) );
  XNOR2_X1 DP_mult_217_U1753 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2028), 
        .ZN(DP_mult_217_n742) );
  OAI22_X1 DP_mult_217_U1752 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1664), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1665), .ZN(DP_mult_217_n2027)
         );
  AOI221_X1 DP_mult_217_U1751 ( .B1(DP_pipe01[5]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[4]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2027), .ZN(
        DP_mult_217_n2026) );
  XNOR2_X1 DP_mult_217_U1750 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2026), 
        .ZN(DP_mult_217_n743) );
  OAI22_X1 DP_mult_217_U1749 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1660), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1661), .ZN(DP_mult_217_n2025)
         );
  AOI221_X1 DP_mult_217_U1748 ( .B1(DP_pipe01[4]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[3]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2025), .ZN(
        DP_mult_217_n2024) );
  XNOR2_X1 DP_mult_217_U1747 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2024), 
        .ZN(DP_mult_217_n744) );
  OAI22_X1 DP_mult_217_U1746 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1657), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1649), .ZN(DP_mult_217_n2023)
         );
  AOI221_X1 DP_mult_217_U1745 ( .B1(DP_pipe01[3]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[2]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2023), .ZN(
        DP_mult_217_n2022) );
  XNOR2_X1 DP_mult_217_U1744 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2022), 
        .ZN(DP_mult_217_n745) );
  INV_X1 DP_mult_217_U1743 ( .A(DP_mult_217_n1396), .ZN(DP_mult_217_n1653) );
  INV_X1 DP_mult_217_U1742 ( .A(DP_pipe01[0]), .ZN(DP_mult_217_n1647) );
  OAI22_X1 DP_mult_217_U1741 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1653), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1567), .ZN(DP_mult_217_n2021)
         );
  AOI221_X1 DP_mult_217_U1740 ( .B1(DP_pipe01[2]), .B2(DP_mult_217_n1559), 
        .C1(DP_pipe01[1]), .C2(DP_mult_217_n1560), .A(DP_mult_217_n2021), .ZN(
        DP_mult_217_n2020) );
  XNOR2_X1 DP_mult_217_U1739 ( .A(DP_mult_217_n1610), .B(DP_mult_217_n2020), 
        .ZN(DP_mult_217_n746) );
  OAI222_X1 DP_mult_217_U1738 ( .A1(DP_mult_217_n1544), .A2(DP_mult_217_n1649), 
        .B1(DP_mult_217_n1550), .B2(DP_mult_217_n1566), .C1(DP_mult_217_n1558), 
        .C2(DP_mult_217_n1650), .ZN(DP_mult_217_n2019) );
  XNOR2_X1 DP_mult_217_U1737 ( .A(DP_mult_217_n2019), .B(DP_mult_217_n1611), 
        .ZN(DP_mult_217_n747) );
  OAI22_X1 DP_mult_217_U1736 ( .A1(DP_mult_217_n1544), .A2(DP_mult_217_n1567), 
        .B1(DP_mult_217_n1558), .B2(DP_mult_217_n1567), .ZN(DP_mult_217_n2018)
         );
  XNOR2_X1 DP_mult_217_U1735 ( .A(DP_mult_217_n2018), .B(DP_mult_217_n1611), 
        .ZN(DP_mult_217_n748) );
  XOR2_X1 DP_mult_217_U1734 ( .A(DP_coeff_pipe01[18]), .B(DP_mult_217_n1607), 
        .Z(DP_mult_217_n2017) );
  XOR2_X1 DP_mult_217_U1733 ( .A(DP_coeff_pipe01[19]), .B(DP_mult_217_n1608), 
        .Z(DP_mult_217_n2016) );
  XNOR2_X1 DP_mult_217_U1732 ( .A(DP_coeff_pipe01[18]), .B(DP_coeff_pipe01[19]), .ZN(DP_mult_217_n2015) );
  NAND3_X1 DP_mult_217_U1731 ( .A1(DP_mult_217_n2017), .A2(DP_mult_217_n2016), 
        .A3(DP_mult_217_n2015), .ZN(DP_mult_217_n1967) );
  INV_X1 DP_mult_217_U1730 ( .A(DP_mult_217_n2017), .ZN(DP_mult_217_n2014) );
  OAI21_X1 DP_mult_217_U1729 ( .B1(DP_mult_217_n1594), .B2(DP_mult_217_n1595), 
        .A(DP_mult_217_n1615), .ZN(DP_mult_217_n2013) );
  OAI221_X1 DP_mult_217_U1728 ( .B1(DP_mult_217_n1617), .B2(DP_mult_217_n1597), 
        .C1(DP_mult_217_n1620), .C2(DP_mult_217_n1593), .A(DP_mult_217_n2013), 
        .ZN(DP_mult_217_n2012) );
  XNOR2_X1 DP_mult_217_U1727 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n2012), 
        .ZN(DP_mult_217_n749) );
  INV_X1 DP_mult_217_U1726 ( .A(DP_mult_217_n1374), .ZN(DP_mult_217_n1633) );
  INV_X1 DP_mult_217_U1725 ( .A(DP_pipe01[22]), .ZN(DP_mult_217_n1634) );
  OAI22_X1 DP_mult_217_U1724 ( .A1(DP_mult_217_n1633), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1634), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n2011)
         );
  AOI221_X1 DP_mult_217_U1723 ( .B1(DP_mult_217_n1594), .B2(DP_mult_217_n1614), 
        .C1(DP_mult_217_n1595), .C2(DP_mult_217_n1615), .A(DP_mult_217_n2011), 
        .ZN(DP_mult_217_n2010) );
  XNOR2_X1 DP_mult_217_U1722 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n2010), 
        .ZN(DP_mult_217_n750) );
  OAI22_X1 DP_mult_217_U1721 ( .A1(DP_mult_217_n1617), .A2(DP_mult_217_n1543), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n2009)
         );
  AOI221_X1 DP_mult_217_U1720 ( .B1(DP_mult_217_n1595), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1547), .C2(DP_mult_217_n1375), .A(DP_mult_217_n2009), 
        .ZN(DP_mult_217_n2008) );
  XNOR2_X1 DP_mult_217_U1719 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n2008), 
        .ZN(DP_mult_217_n751) );
  OAI22_X1 DP_mult_217_U1718 ( .A1(DP_mult_217_n1640), .A2(DP_mult_217_n1597), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1552), .ZN(DP_mult_217_n2007)
         );
  AOI221_X1 DP_mult_217_U1717 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1547), .C2(DP_mult_217_n1376), .A(DP_mult_217_n2007), 
        .ZN(DP_mult_217_n2006) );
  XNOR2_X1 DP_mult_217_U1716 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n2006), 
        .ZN(DP_mult_217_n752) );
  OAI22_X1 DP_mult_217_U1715 ( .A1(DP_mult_217_n1728), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1729), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n2005)
         );
  AOI221_X1 DP_mult_217_U1714 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[21]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[20]), .A(DP_mult_217_n2005), 
        .ZN(DP_mult_217_n2004) );
  XNOR2_X1 DP_mult_217_U1713 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n2004), 
        .ZN(DP_mult_217_n753) );
  OAI22_X1 DP_mult_217_U1712 ( .A1(DP_mult_217_n1724), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1725), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n2003)
         );
  AOI221_X1 DP_mult_217_U1711 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[20]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[19]), .A(DP_mult_217_n2003), 
        .ZN(DP_mult_217_n2002) );
  XNOR2_X1 DP_mult_217_U1710 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n2002), 
        .ZN(DP_mult_217_n754) );
  OAI22_X1 DP_mult_217_U1709 ( .A1(DP_mult_217_n1720), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1721), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n2001)
         );
  AOI221_X1 DP_mult_217_U1708 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[19]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[18]), .A(DP_mult_217_n2001), 
        .ZN(DP_mult_217_n2000) );
  XNOR2_X1 DP_mult_217_U1707 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n2000), 
        .ZN(DP_mult_217_n755) );
  OAI22_X1 DP_mult_217_U1706 ( .A1(DP_mult_217_n1716), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1717), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n1999)
         );
  AOI221_X1 DP_mult_217_U1705 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[18]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[17]), .A(DP_mult_217_n1999), 
        .ZN(DP_mult_217_n1998) );
  XNOR2_X1 DP_mult_217_U1704 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n1998), 
        .ZN(DP_mult_217_n756) );
  OAI22_X1 DP_mult_217_U1703 ( .A1(DP_mult_217_n1712), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1713), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n1997)
         );
  AOI221_X1 DP_mult_217_U1702 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[17]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[16]), .A(DP_mult_217_n1997), 
        .ZN(DP_mult_217_n1996) );
  XNOR2_X1 DP_mult_217_U1701 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n1996), 
        .ZN(DP_mult_217_n757) );
  OAI22_X1 DP_mult_217_U1700 ( .A1(DP_mult_217_n1708), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1709), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n1995)
         );
  AOI221_X1 DP_mult_217_U1699 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[16]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[15]), .A(DP_mult_217_n1995), 
        .ZN(DP_mult_217_n1994) );
  XNOR2_X1 DP_mult_217_U1698 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n1994), 
        .ZN(DP_mult_217_n758) );
  OAI22_X1 DP_mult_217_U1697 ( .A1(DP_mult_217_n1704), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1705), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n1993)
         );
  AOI221_X1 DP_mult_217_U1696 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[15]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[14]), .A(DP_mult_217_n1993), 
        .ZN(DP_mult_217_n1992) );
  XNOR2_X1 DP_mult_217_U1695 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n1992), 
        .ZN(DP_mult_217_n759) );
  OAI22_X1 DP_mult_217_U1694 ( .A1(DP_mult_217_n1700), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1701), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n1991)
         );
  AOI221_X1 DP_mult_217_U1693 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[14]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[13]), .A(DP_mult_217_n1991), 
        .ZN(DP_mult_217_n1990) );
  XNOR2_X1 DP_mult_217_U1692 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n1990), 
        .ZN(DP_mult_217_n760) );
  OAI22_X1 DP_mult_217_U1691 ( .A1(DP_mult_217_n1696), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1697), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n1989)
         );
  AOI221_X1 DP_mult_217_U1690 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[13]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[12]), .A(DP_mult_217_n1989), 
        .ZN(DP_mult_217_n1988) );
  XNOR2_X1 DP_mult_217_U1689 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n1988), 
        .ZN(DP_mult_217_n761) );
  OAI22_X1 DP_mult_217_U1688 ( .A1(DP_mult_217_n1692), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1693), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1987)
         );
  AOI221_X1 DP_mult_217_U1687 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[12]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[11]), .A(DP_mult_217_n1987), 
        .ZN(DP_mult_217_n1986) );
  XNOR2_X1 DP_mult_217_U1686 ( .A(DP_mult_217_n1609), .B(DP_mult_217_n1986), 
        .ZN(DP_mult_217_n762) );
  OAI22_X1 DP_mult_217_U1685 ( .A1(DP_mult_217_n1688), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1689), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1985)
         );
  AOI221_X1 DP_mult_217_U1684 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[11]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[10]), .A(DP_mult_217_n1985), 
        .ZN(DP_mult_217_n1984) );
  XNOR2_X1 DP_mult_217_U1683 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1984), 
        .ZN(DP_mult_217_n763) );
  OAI22_X1 DP_mult_217_U1682 ( .A1(DP_mult_217_n1684), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1685), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1983)
         );
  AOI221_X1 DP_mult_217_U1681 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[10]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[9]), .A(DP_mult_217_n1983), .ZN(
        DP_mult_217_n1982) );
  XNOR2_X1 DP_mult_217_U1680 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1982), 
        .ZN(DP_mult_217_n764) );
  OAI22_X1 DP_mult_217_U1679 ( .A1(DP_mult_217_n1680), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1681), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1981)
         );
  AOI221_X1 DP_mult_217_U1678 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[9]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[8]), .A(DP_mult_217_n1981), .ZN(
        DP_mult_217_n1980) );
  XNOR2_X1 DP_mult_217_U1677 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1980), 
        .ZN(DP_mult_217_n765) );
  OAI22_X1 DP_mult_217_U1676 ( .A1(DP_mult_217_n1676), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1677), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1979)
         );
  AOI221_X1 DP_mult_217_U1675 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[8]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[7]), .A(DP_mult_217_n1979), .ZN(
        DP_mult_217_n1978) );
  XNOR2_X1 DP_mult_217_U1674 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1978), 
        .ZN(DP_mult_217_n766) );
  OAI22_X1 DP_mult_217_U1673 ( .A1(DP_mult_217_n1672), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1673), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1977)
         );
  AOI221_X1 DP_mult_217_U1672 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[7]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[6]), .A(DP_mult_217_n1977), .ZN(
        DP_mult_217_n1976) );
  XNOR2_X1 DP_mult_217_U1671 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1976), 
        .ZN(DP_mult_217_n767) );
  OAI22_X1 DP_mult_217_U1670 ( .A1(DP_mult_217_n1668), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1669), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1975)
         );
  AOI221_X1 DP_mult_217_U1669 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[6]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[5]), .A(DP_mult_217_n1975), .ZN(
        DP_mult_217_n1974) );
  XNOR2_X1 DP_mult_217_U1668 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1974), 
        .ZN(DP_mult_217_n768) );
  OAI22_X1 DP_mult_217_U1667 ( .A1(DP_mult_217_n1664), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1665), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1973)
         );
  AOI221_X1 DP_mult_217_U1666 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[5]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[4]), .A(DP_mult_217_n1973), .ZN(
        DP_mult_217_n1972) );
  XNOR2_X1 DP_mult_217_U1665 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1972), 
        .ZN(DP_mult_217_n769) );
  OAI22_X1 DP_mult_217_U1664 ( .A1(DP_mult_217_n1660), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1661), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1971)
         );
  AOI221_X1 DP_mult_217_U1663 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[4]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[3]), .A(DP_mult_217_n1971), .ZN(
        DP_mult_217_n1970) );
  XNOR2_X1 DP_mult_217_U1662 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1970), 
        .ZN(DP_mult_217_n770) );
  OAI22_X1 DP_mult_217_U1661 ( .A1(DP_mult_217_n1657), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1649), .B2(DP_mult_217_n1597), .ZN(DP_mult_217_n1969)
         );
  AOI221_X1 DP_mult_217_U1660 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[3]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[2]), .A(DP_mult_217_n1969), .ZN(
        DP_mult_217_n1968) );
  XNOR2_X1 DP_mult_217_U1659 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1968), 
        .ZN(DP_mult_217_n771) );
  OAI22_X1 DP_mult_217_U1658 ( .A1(DP_mult_217_n1653), .A2(DP_mult_217_n1593), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1596), .ZN(DP_mult_217_n1966)
         );
  AOI221_X1 DP_mult_217_U1657 ( .B1(DP_mult_217_n1594), .B2(DP_pipe01[2]), 
        .C1(DP_mult_217_n1595), .C2(DP_pipe01[1]), .A(DP_mult_217_n1966), .ZN(
        DP_mult_217_n1965) );
  XNOR2_X1 DP_mult_217_U1656 ( .A(DP_mult_217_n1608), .B(DP_mult_217_n1965), 
        .ZN(DP_mult_217_n772) );
  OAI222_X1 DP_mult_217_U1655 ( .A1(DP_mult_217_n1649), .A2(DP_mult_217_n1543), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1552), .C1(DP_mult_217_n1650), 
        .C2(DP_mult_217_n1593), .ZN(DP_mult_217_n1964) );
  XOR2_X1 DP_mult_217_U1654 ( .A(DP_mult_217_n1964), .B(DP_mult_217_n1608), 
        .Z(DP_mult_217_n773) );
  OAI22_X1 DP_mult_217_U1653 ( .A1(DP_mult_217_n1565), .A2(DP_mult_217_n1543), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1593), .ZN(DP_mult_217_n1963)
         );
  XOR2_X1 DP_mult_217_U1652 ( .A(DP_mult_217_n1963), .B(DP_mult_217_n1608), 
        .Z(DP_mult_217_n774) );
  XOR2_X1 DP_mult_217_U1651 ( .A(DP_coeff_pipe01[15]), .B(DP_mult_217_n1605), 
        .Z(DP_mult_217_n1962) );
  XNOR2_X1 DP_mult_217_U1650 ( .A(DP_coeff_pipe01[16]), .B(DP_mult_217_n1607), 
        .ZN(DP_mult_217_n1961) );
  XNOR2_X1 DP_mult_217_U1649 ( .A(DP_coeff_pipe01[15]), .B(DP_coeff_pipe01[16]), .ZN(DP_mult_217_n1960) );
  NAND3_X1 DP_mult_217_U1648 ( .A1(DP_mult_217_n1962), .A2(DP_mult_217_n1961), 
        .A3(DP_mult_217_n1960), .ZN(DP_mult_217_n1912) );
  INV_X1 DP_mult_217_U1647 ( .A(DP_mult_217_n1962), .ZN(DP_mult_217_n1959) );
  OAI21_X1 DP_mult_217_U1646 ( .B1(DP_mult_217_n1589), .B2(DP_mult_217_n1590), 
        .A(DP_mult_217_n1615), .ZN(DP_mult_217_n1958) );
  OAI221_X1 DP_mult_217_U1645 ( .B1(DP_mult_217_n1619), .B2(DP_mult_217_n1592), 
        .C1(DP_mult_217_n1617), .C2(DP_mult_217_n1588), .A(DP_mult_217_n1958), 
        .ZN(DP_mult_217_n1957) );
  XNOR2_X1 DP_mult_217_U1644 ( .A(DP_coeff_pipe01[17]), .B(DP_mult_217_n1957), 
        .ZN(DP_mult_217_n775) );
  OAI22_X1 DP_mult_217_U1643 ( .A1(DP_mult_217_n1633), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1634), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1956)
         );
  AOI221_X1 DP_mult_217_U1642 ( .B1(DP_mult_217_n1589), .B2(DP_mult_217_n1614), 
        .C1(DP_mult_217_n1590), .C2(DP_mult_217_n1615), .A(DP_mult_217_n1956), 
        .ZN(DP_mult_217_n1955) );
  XNOR2_X1 DP_mult_217_U1641 ( .A(DP_coeff_pipe01[17]), .B(DP_mult_217_n1955), 
        .ZN(DP_mult_217_n776) );
  OAI22_X1 DP_mult_217_U1640 ( .A1(DP_mult_217_n1617), .A2(DP_mult_217_n1546), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1954)
         );
  AOI221_X1 DP_mult_217_U1639 ( .B1(DP_mult_217_n1590), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1549), .C2(DP_mult_217_n1375), .A(DP_mult_217_n1954), 
        .ZN(DP_mult_217_n1953) );
  XNOR2_X1 DP_mult_217_U1638 ( .A(DP_coeff_pipe01[17]), .B(DP_mult_217_n1953), 
        .ZN(DP_mult_217_n777) );
  OAI22_X1 DP_mult_217_U1637 ( .A1(DP_mult_217_n1640), .A2(DP_mult_217_n1592), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1551), .ZN(DP_mult_217_n1952)
         );
  AOI221_X1 DP_mult_217_U1636 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1549), .C2(DP_mult_217_n1376), .A(DP_mult_217_n1952), 
        .ZN(DP_mult_217_n1951) );
  XNOR2_X1 DP_mult_217_U1635 ( .A(DP_coeff_pipe01[17]), .B(DP_mult_217_n1951), 
        .ZN(DP_mult_217_n778) );
  OAI22_X1 DP_mult_217_U1634 ( .A1(DP_mult_217_n1728), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1729), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1950)
         );
  AOI221_X1 DP_mult_217_U1633 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[21]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[20]), .A(DP_mult_217_n1950), 
        .ZN(DP_mult_217_n1949) );
  XNOR2_X1 DP_mult_217_U1632 ( .A(DP_coeff_pipe01[17]), .B(DP_mult_217_n1949), 
        .ZN(DP_mult_217_n779) );
  OAI22_X1 DP_mult_217_U1631 ( .A1(DP_mult_217_n1724), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1725), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1948)
         );
  AOI221_X1 DP_mult_217_U1630 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[20]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[19]), .A(DP_mult_217_n1948), 
        .ZN(DP_mult_217_n1947) );
  XNOR2_X1 DP_mult_217_U1629 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1947), 
        .ZN(DP_mult_217_n780) );
  OAI22_X1 DP_mult_217_U1628 ( .A1(DP_mult_217_n1720), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1721), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1946)
         );
  AOI221_X1 DP_mult_217_U1627 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[19]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[18]), .A(DP_mult_217_n1946), 
        .ZN(DP_mult_217_n1945) );
  XNOR2_X1 DP_mult_217_U1626 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1945), 
        .ZN(DP_mult_217_n781) );
  OAI22_X1 DP_mult_217_U1625 ( .A1(DP_mult_217_n1716), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1717), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1944)
         );
  AOI221_X1 DP_mult_217_U1624 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[18]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[17]), .A(DP_mult_217_n1944), 
        .ZN(DP_mult_217_n1943) );
  XNOR2_X1 DP_mult_217_U1623 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1943), 
        .ZN(DP_mult_217_n782) );
  OAI22_X1 DP_mult_217_U1622 ( .A1(DP_mult_217_n1712), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1713), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1942)
         );
  AOI221_X1 DP_mult_217_U1621 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[17]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[16]), .A(DP_mult_217_n1942), 
        .ZN(DP_mult_217_n1941) );
  XNOR2_X1 DP_mult_217_U1620 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1941), 
        .ZN(DP_mult_217_n783) );
  OAI22_X1 DP_mult_217_U1619 ( .A1(DP_mult_217_n1708), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1709), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1940)
         );
  AOI221_X1 DP_mult_217_U1618 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[16]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[15]), .A(DP_mult_217_n1940), 
        .ZN(DP_mult_217_n1939) );
  XNOR2_X1 DP_mult_217_U1617 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1939), 
        .ZN(DP_mult_217_n784) );
  OAI22_X1 DP_mult_217_U1616 ( .A1(DP_mult_217_n1704), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1705), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1938)
         );
  AOI221_X1 DP_mult_217_U1615 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[15]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[14]), .A(DP_mult_217_n1938), 
        .ZN(DP_mult_217_n1937) );
  XNOR2_X1 DP_mult_217_U1614 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1937), 
        .ZN(DP_mult_217_n785) );
  OAI22_X1 DP_mult_217_U1613 ( .A1(DP_mult_217_n1700), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1701), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1936)
         );
  AOI221_X1 DP_mult_217_U1612 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[14]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[13]), .A(DP_mult_217_n1936), 
        .ZN(DP_mult_217_n1935) );
  XNOR2_X1 DP_mult_217_U1611 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1935), 
        .ZN(DP_mult_217_n786) );
  OAI22_X1 DP_mult_217_U1610 ( .A1(DP_mult_217_n1696), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1697), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1934)
         );
  AOI221_X1 DP_mult_217_U1609 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[13]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[12]), .A(DP_mult_217_n1934), 
        .ZN(DP_mult_217_n1933) );
  XNOR2_X1 DP_mult_217_U1608 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1933), 
        .ZN(DP_mult_217_n787) );
  OAI22_X1 DP_mult_217_U1607 ( .A1(DP_mult_217_n1692), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1693), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1932)
         );
  AOI221_X1 DP_mult_217_U1606 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[12]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[11]), .A(DP_mult_217_n1932), 
        .ZN(DP_mult_217_n1931) );
  XNOR2_X1 DP_mult_217_U1605 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1931), 
        .ZN(DP_mult_217_n788) );
  OAI22_X1 DP_mult_217_U1604 ( .A1(DP_mult_217_n1688), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1689), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1930)
         );
  AOI221_X1 DP_mult_217_U1603 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[11]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[10]), .A(DP_mult_217_n1930), 
        .ZN(DP_mult_217_n1929) );
  XNOR2_X1 DP_mult_217_U1602 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1929), 
        .ZN(DP_mult_217_n789) );
  OAI22_X1 DP_mult_217_U1601 ( .A1(DP_mult_217_n1684), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1685), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1928)
         );
  AOI221_X1 DP_mult_217_U1600 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[10]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[9]), .A(DP_mult_217_n1928), .ZN(
        DP_mult_217_n1927) );
  XNOR2_X1 DP_mult_217_U1599 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1927), 
        .ZN(DP_mult_217_n790) );
  OAI22_X1 DP_mult_217_U1598 ( .A1(DP_mult_217_n1680), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1681), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1926)
         );
  AOI221_X1 DP_mult_217_U1597 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[9]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[8]), .A(DP_mult_217_n1926), .ZN(
        DP_mult_217_n1925) );
  XNOR2_X1 DP_mult_217_U1596 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1925), 
        .ZN(DP_mult_217_n791) );
  OAI22_X1 DP_mult_217_U1595 ( .A1(DP_mult_217_n1676), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1677), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1924)
         );
  AOI221_X1 DP_mult_217_U1594 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[8]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[7]), .A(DP_mult_217_n1924), .ZN(
        DP_mult_217_n1923) );
  XNOR2_X1 DP_mult_217_U1593 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1923), 
        .ZN(DP_mult_217_n792) );
  OAI22_X1 DP_mult_217_U1592 ( .A1(DP_mult_217_n1672), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1673), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1922)
         );
  AOI221_X1 DP_mult_217_U1591 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[7]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[6]), .A(DP_mult_217_n1922), .ZN(
        DP_mult_217_n1921) );
  XNOR2_X1 DP_mult_217_U1590 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1921), 
        .ZN(DP_mult_217_n793) );
  OAI22_X1 DP_mult_217_U1589 ( .A1(DP_mult_217_n1668), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1669), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1920)
         );
  AOI221_X1 DP_mult_217_U1588 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[6]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[5]), .A(DP_mult_217_n1920), .ZN(
        DP_mult_217_n1919) );
  XNOR2_X1 DP_mult_217_U1587 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1919), 
        .ZN(DP_mult_217_n794) );
  OAI22_X1 DP_mult_217_U1586 ( .A1(DP_mult_217_n1664), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1665), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1918)
         );
  AOI221_X1 DP_mult_217_U1585 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[5]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[4]), .A(DP_mult_217_n1918), .ZN(
        DP_mult_217_n1917) );
  XNOR2_X1 DP_mult_217_U1584 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1917), 
        .ZN(DP_mult_217_n795) );
  OAI22_X1 DP_mult_217_U1583 ( .A1(DP_mult_217_n1660), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1661), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1916)
         );
  AOI221_X1 DP_mult_217_U1582 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[4]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[3]), .A(DP_mult_217_n1916), .ZN(
        DP_mult_217_n1915) );
  XNOR2_X1 DP_mult_217_U1581 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1915), 
        .ZN(DP_mult_217_n796) );
  OAI22_X1 DP_mult_217_U1580 ( .A1(DP_mult_217_n1657), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1649), .B2(DP_mult_217_n1592), .ZN(DP_mult_217_n1914)
         );
  AOI221_X1 DP_mult_217_U1579 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[3]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[2]), .A(DP_mult_217_n1914), .ZN(
        DP_mult_217_n1913) );
  XNOR2_X1 DP_mult_217_U1578 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1913), 
        .ZN(DP_mult_217_n797) );
  OAI22_X1 DP_mult_217_U1577 ( .A1(DP_mult_217_n1653), .A2(DP_mult_217_n1588), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1591), .ZN(DP_mult_217_n1911)
         );
  AOI221_X1 DP_mult_217_U1576 ( .B1(DP_mult_217_n1589), .B2(DP_pipe01[2]), 
        .C1(DP_mult_217_n1590), .C2(DP_pipe01[1]), .A(DP_mult_217_n1911), .ZN(
        DP_mult_217_n1910) );
  XNOR2_X1 DP_mult_217_U1575 ( .A(DP_mult_217_n1606), .B(DP_mult_217_n1910), 
        .ZN(DP_mult_217_n798) );
  OAI222_X1 DP_mult_217_U1574 ( .A1(DP_mult_217_n1649), .A2(DP_mult_217_n1546), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1551), .C1(DP_mult_217_n1650), 
        .C2(DP_mult_217_n1588), .ZN(DP_mult_217_n1909) );
  XNOR2_X1 DP_mult_217_U1573 ( .A(DP_mult_217_n1909), .B(DP_mult_217_n1607), 
        .ZN(DP_mult_217_n799) );
  OAI22_X1 DP_mult_217_U1572 ( .A1(DP_mult_217_n1565), .A2(DP_mult_217_n1546), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1588), .ZN(DP_mult_217_n1908)
         );
  XNOR2_X1 DP_mult_217_U1571 ( .A(DP_mult_217_n1908), .B(DP_mult_217_n1607), 
        .ZN(DP_mult_217_n800) );
  XOR2_X1 DP_mult_217_U1570 ( .A(DP_coeff_pipe01[12]), .B(DP_mult_217_n1603), 
        .Z(DP_mult_217_n1907) );
  XNOR2_X1 DP_mult_217_U1569 ( .A(DP_coeff_pipe01[13]), .B(DP_mult_217_n1605), 
        .ZN(DP_mult_217_n1906) );
  XNOR2_X1 DP_mult_217_U1568 ( .A(DP_coeff_pipe01[12]), .B(DP_coeff_pipe01[13]), .ZN(DP_mult_217_n1905) );
  NAND3_X1 DP_mult_217_U1567 ( .A1(DP_mult_217_n1907), .A2(DP_mult_217_n1906), 
        .A3(DP_mult_217_n1905), .ZN(DP_mult_217_n1857) );
  INV_X1 DP_mult_217_U1566 ( .A(DP_mult_217_n1907), .ZN(DP_mult_217_n1904) );
  OAI21_X1 DP_mult_217_U1565 ( .B1(DP_mult_217_n1584), .B2(DP_mult_217_n1585), 
        .A(DP_mult_217_n1615), .ZN(DP_mult_217_n1903) );
  OAI221_X1 DP_mult_217_U1564 ( .B1(DP_mult_217_n1617), .B2(DP_mult_217_n1587), 
        .C1(DP_mult_217_n1620), .C2(DP_mult_217_n1583), .A(DP_mult_217_n1903), 
        .ZN(DP_mult_217_n1902) );
  XNOR2_X1 DP_mult_217_U1563 ( .A(DP_coeff_pipe01[14]), .B(DP_mult_217_n1902), 
        .ZN(DP_mult_217_n801) );
  OAI22_X1 DP_mult_217_U1562 ( .A1(DP_mult_217_n1633), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1634), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1901)
         );
  AOI221_X1 DP_mult_217_U1561 ( .B1(DP_mult_217_n1584), .B2(DP_mult_217_n1615), 
        .C1(DP_mult_217_n1585), .C2(DP_mult_217_n1615), .A(DP_mult_217_n1901), 
        .ZN(DP_mult_217_n1900) );
  XNOR2_X1 DP_mult_217_U1560 ( .A(DP_coeff_pipe01[14]), .B(DP_mult_217_n1900), 
        .ZN(DP_mult_217_n802) );
  OAI22_X1 DP_mult_217_U1559 ( .A1(DP_mult_217_n1617), .A2(DP_mult_217_n1545), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1899)
         );
  AOI221_X1 DP_mult_217_U1558 ( .B1(DP_mult_217_n1585), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1548), .C2(DP_mult_217_n1375), .A(DP_mult_217_n1899), 
        .ZN(DP_mult_217_n1898) );
  XNOR2_X1 DP_mult_217_U1557 ( .A(DP_coeff_pipe01[14]), .B(DP_mult_217_n1898), 
        .ZN(DP_mult_217_n803) );
  OAI22_X1 DP_mult_217_U1556 ( .A1(DP_mult_217_n1640), .A2(DP_mult_217_n1587), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1555), .ZN(DP_mult_217_n1897)
         );
  AOI221_X1 DP_mult_217_U1555 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1548), .C2(DP_mult_217_n1376), .A(DP_mult_217_n1897), 
        .ZN(DP_mult_217_n1896) );
  XNOR2_X1 DP_mult_217_U1554 ( .A(DP_coeff_pipe01[14]), .B(DP_mult_217_n1896), 
        .ZN(DP_mult_217_n804) );
  OAI22_X1 DP_mult_217_U1553 ( .A1(DP_mult_217_n1728), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1729), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1895)
         );
  AOI221_X1 DP_mult_217_U1552 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[21]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[20]), .A(DP_mult_217_n1895), 
        .ZN(DP_mult_217_n1894) );
  XNOR2_X1 DP_mult_217_U1551 ( .A(DP_coeff_pipe01[14]), .B(DP_mult_217_n1894), 
        .ZN(DP_mult_217_n805) );
  OAI22_X1 DP_mult_217_U1550 ( .A1(DP_mult_217_n1724), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1725), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1893)
         );
  AOI221_X1 DP_mult_217_U1549 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[20]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[19]), .A(DP_mult_217_n1893), 
        .ZN(DP_mult_217_n1892) );
  XNOR2_X1 DP_mult_217_U1548 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1892), 
        .ZN(DP_mult_217_n806) );
  OAI22_X1 DP_mult_217_U1547 ( .A1(DP_mult_217_n1720), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1721), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1891)
         );
  AOI221_X1 DP_mult_217_U1546 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[19]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[18]), .A(DP_mult_217_n1891), 
        .ZN(DP_mult_217_n1890) );
  XNOR2_X1 DP_mult_217_U1545 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1890), 
        .ZN(DP_mult_217_n807) );
  OAI22_X1 DP_mult_217_U1544 ( .A1(DP_mult_217_n1716), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1717), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1889)
         );
  AOI221_X1 DP_mult_217_U1543 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[18]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[17]), .A(DP_mult_217_n1889), 
        .ZN(DP_mult_217_n1888) );
  XNOR2_X1 DP_mult_217_U1542 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1888), 
        .ZN(DP_mult_217_n808) );
  OAI22_X1 DP_mult_217_U1541 ( .A1(DP_mult_217_n1712), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1713), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1887)
         );
  AOI221_X1 DP_mult_217_U1540 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[17]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[16]), .A(DP_mult_217_n1887), 
        .ZN(DP_mult_217_n1886) );
  XNOR2_X1 DP_mult_217_U1539 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1886), 
        .ZN(DP_mult_217_n809) );
  OAI22_X1 DP_mult_217_U1538 ( .A1(DP_mult_217_n1708), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1709), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1885)
         );
  AOI221_X1 DP_mult_217_U1537 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[16]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[15]), .A(DP_mult_217_n1885), 
        .ZN(DP_mult_217_n1884) );
  XNOR2_X1 DP_mult_217_U1536 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1884), 
        .ZN(DP_mult_217_n810) );
  OAI22_X1 DP_mult_217_U1535 ( .A1(DP_mult_217_n1704), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1705), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1883)
         );
  AOI221_X1 DP_mult_217_U1534 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[15]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[14]), .A(DP_mult_217_n1883), 
        .ZN(DP_mult_217_n1882) );
  XNOR2_X1 DP_mult_217_U1533 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1882), 
        .ZN(DP_mult_217_n811) );
  OAI22_X1 DP_mult_217_U1532 ( .A1(DP_mult_217_n1700), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1701), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1881)
         );
  AOI221_X1 DP_mult_217_U1531 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[14]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[13]), .A(DP_mult_217_n1881), 
        .ZN(DP_mult_217_n1880) );
  XNOR2_X1 DP_mult_217_U1530 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1880), 
        .ZN(DP_mult_217_n812) );
  OAI22_X1 DP_mult_217_U1529 ( .A1(DP_mult_217_n1696), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1697), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1879)
         );
  AOI221_X1 DP_mult_217_U1528 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[13]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[12]), .A(DP_mult_217_n1879), 
        .ZN(DP_mult_217_n1878) );
  XNOR2_X1 DP_mult_217_U1527 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1878), 
        .ZN(DP_mult_217_n813) );
  OAI22_X1 DP_mult_217_U1526 ( .A1(DP_mult_217_n1692), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1693), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1877)
         );
  AOI221_X1 DP_mult_217_U1525 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[12]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[11]), .A(DP_mult_217_n1877), 
        .ZN(DP_mult_217_n1876) );
  XNOR2_X1 DP_mult_217_U1524 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1876), 
        .ZN(DP_mult_217_n814) );
  OAI22_X1 DP_mult_217_U1523 ( .A1(DP_mult_217_n1688), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1689), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1875)
         );
  AOI221_X1 DP_mult_217_U1522 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[11]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[10]), .A(DP_mult_217_n1875), 
        .ZN(DP_mult_217_n1874) );
  XNOR2_X1 DP_mult_217_U1521 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1874), 
        .ZN(DP_mult_217_n815) );
  OAI22_X1 DP_mult_217_U1520 ( .A1(DP_mult_217_n1684), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1685), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1873)
         );
  AOI221_X1 DP_mult_217_U1519 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[10]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[9]), .A(DP_mult_217_n1873), .ZN(
        DP_mult_217_n1872) );
  XNOR2_X1 DP_mult_217_U1518 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1872), 
        .ZN(DP_mult_217_n816) );
  OAI22_X1 DP_mult_217_U1517 ( .A1(DP_mult_217_n1680), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1681), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1871)
         );
  AOI221_X1 DP_mult_217_U1516 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[9]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[8]), .A(DP_mult_217_n1871), .ZN(
        DP_mult_217_n1870) );
  XNOR2_X1 DP_mult_217_U1515 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1870), 
        .ZN(DP_mult_217_n817) );
  OAI22_X1 DP_mult_217_U1514 ( .A1(DP_mult_217_n1676), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1677), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1869)
         );
  AOI221_X1 DP_mult_217_U1513 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[8]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[7]), .A(DP_mult_217_n1869), .ZN(
        DP_mult_217_n1868) );
  XNOR2_X1 DP_mult_217_U1512 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1868), 
        .ZN(DP_mult_217_n818) );
  OAI22_X1 DP_mult_217_U1511 ( .A1(DP_mult_217_n1672), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1673), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1867)
         );
  AOI221_X1 DP_mult_217_U1510 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[7]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[6]), .A(DP_mult_217_n1867), .ZN(
        DP_mult_217_n1866) );
  XNOR2_X1 DP_mult_217_U1509 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1866), 
        .ZN(DP_mult_217_n819) );
  OAI22_X1 DP_mult_217_U1508 ( .A1(DP_mult_217_n1668), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1669), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1865)
         );
  AOI221_X1 DP_mult_217_U1507 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[6]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[5]), .A(DP_mult_217_n1865), .ZN(
        DP_mult_217_n1864) );
  XNOR2_X1 DP_mult_217_U1506 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1864), 
        .ZN(DP_mult_217_n820) );
  OAI22_X1 DP_mult_217_U1505 ( .A1(DP_mult_217_n1664), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1665), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1863)
         );
  AOI221_X1 DP_mult_217_U1504 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[5]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[4]), .A(DP_mult_217_n1863), .ZN(
        DP_mult_217_n1862) );
  XNOR2_X1 DP_mult_217_U1503 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1862), 
        .ZN(DP_mult_217_n821) );
  OAI22_X1 DP_mult_217_U1502 ( .A1(DP_mult_217_n1660), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1661), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1861)
         );
  AOI221_X1 DP_mult_217_U1501 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[4]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[3]), .A(DP_mult_217_n1861), .ZN(
        DP_mult_217_n1860) );
  XNOR2_X1 DP_mult_217_U1500 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1860), 
        .ZN(DP_mult_217_n822) );
  OAI22_X1 DP_mult_217_U1499 ( .A1(DP_mult_217_n1657), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1649), .B2(DP_mult_217_n1587), .ZN(DP_mult_217_n1859)
         );
  AOI221_X1 DP_mult_217_U1498 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[3]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[2]), .A(DP_mult_217_n1859), .ZN(
        DP_mult_217_n1858) );
  XNOR2_X1 DP_mult_217_U1497 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1858), 
        .ZN(DP_mult_217_n823) );
  OAI22_X1 DP_mult_217_U1496 ( .A1(DP_mult_217_n1653), .A2(DP_mult_217_n1583), 
        .B1(DP_mult_217_n1565), .B2(DP_mult_217_n1586), .ZN(DP_mult_217_n1856)
         );
  AOI221_X1 DP_mult_217_U1495 ( .B1(DP_mult_217_n1584), .B2(DP_pipe01[2]), 
        .C1(DP_mult_217_n1585), .C2(DP_pipe01[1]), .A(DP_mult_217_n1856), .ZN(
        DP_mult_217_n1855) );
  XNOR2_X1 DP_mult_217_U1494 ( .A(DP_mult_217_n1604), .B(DP_mult_217_n1855), 
        .ZN(DP_mult_217_n824) );
  OAI222_X1 DP_mult_217_U1493 ( .A1(DP_mult_217_n1649), .A2(DP_mult_217_n1545), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1555), .C1(DP_mult_217_n1650), 
        .C2(DP_mult_217_n1583), .ZN(DP_mult_217_n1854) );
  XNOR2_X1 DP_mult_217_U1492 ( .A(DP_mult_217_n1854), .B(DP_mult_217_n1605), 
        .ZN(DP_mult_217_n825) );
  OAI22_X1 DP_mult_217_U1491 ( .A1(DP_mult_217_n1565), .A2(DP_mult_217_n1545), 
        .B1(DP_mult_217_n1565), .B2(DP_mult_217_n1583), .ZN(DP_mult_217_n1853)
         );
  XNOR2_X1 DP_mult_217_U1490 ( .A(DP_mult_217_n1853), .B(DP_mult_217_n1605), 
        .ZN(DP_mult_217_n826) );
  XOR2_X1 DP_mult_217_U1489 ( .A(DP_coeff_pipe01[9]), .B(DP_mult_217_n1601), 
        .Z(DP_mult_217_n1852) );
  XNOR2_X1 DP_mult_217_U1488 ( .A(DP_coeff_pipe01[10]), .B(DP_mult_217_n1603), 
        .ZN(DP_mult_217_n1851) );
  XNOR2_X1 DP_mult_217_U1487 ( .A(DP_coeff_pipe01[10]), .B(DP_coeff_pipe01[9]), 
        .ZN(DP_mult_217_n1850) );
  NAND3_X1 DP_mult_217_U1486 ( .A1(DP_mult_217_n1852), .A2(DP_mult_217_n1851), 
        .A3(DP_mult_217_n1850), .ZN(DP_mult_217_n1802) );
  INV_X1 DP_mult_217_U1485 ( .A(DP_mult_217_n1852), .ZN(DP_mult_217_n1849) );
  OAI21_X1 DP_mult_217_U1484 ( .B1(DP_mult_217_n1579), .B2(DP_mult_217_n1580), 
        .A(DP_mult_217_n1615), .ZN(DP_mult_217_n1848) );
  OAI221_X1 DP_mult_217_U1483 ( .B1(DP_mult_217_n1618), .B2(DP_mult_217_n1582), 
        .C1(DP_mult_217_n1617), .C2(DP_mult_217_n1578), .A(DP_mult_217_n1848), 
        .ZN(DP_mult_217_n1847) );
  XNOR2_X1 DP_mult_217_U1482 ( .A(DP_coeff_pipe01[11]), .B(DP_mult_217_n1847), 
        .ZN(DP_mult_217_n827) );
  OAI22_X1 DP_mult_217_U1481 ( .A1(DP_mult_217_n1633), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1634), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1846)
         );
  AOI221_X1 DP_mult_217_U1480 ( .B1(DP_mult_217_n1579), .B2(DP_mult_217_n1615), 
        .C1(DP_mult_217_n1580), .C2(DP_mult_217_n1615), .A(DP_mult_217_n1846), 
        .ZN(DP_mult_217_n1845) );
  XNOR2_X1 DP_mult_217_U1479 ( .A(DP_coeff_pipe01[11]), .B(DP_mult_217_n1845), 
        .ZN(DP_mult_217_n828) );
  OAI22_X1 DP_mult_217_U1478 ( .A1(DP_mult_217_n1617), .A2(DP_mult_217_n1540), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1844)
         );
  AOI221_X1 DP_mult_217_U1477 ( .B1(DP_mult_217_n1580), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1541), .C2(DP_mult_217_n1375), .A(DP_mult_217_n1844), 
        .ZN(DP_mult_217_n1843) );
  XNOR2_X1 DP_mult_217_U1476 ( .A(DP_coeff_pipe01[11]), .B(DP_mult_217_n1843), 
        .ZN(DP_mult_217_n829) );
  OAI22_X1 DP_mult_217_U1475 ( .A1(DP_mult_217_n1640), .A2(DP_mult_217_n1582), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1533), .ZN(DP_mult_217_n1842)
         );
  AOI221_X1 DP_mult_217_U1474 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1541), .C2(DP_mult_217_n1376), .A(DP_mult_217_n1842), 
        .ZN(DP_mult_217_n1841) );
  XNOR2_X1 DP_mult_217_U1473 ( .A(DP_coeff_pipe01[11]), .B(DP_mult_217_n1841), 
        .ZN(DP_mult_217_n830) );
  OAI22_X1 DP_mult_217_U1472 ( .A1(DP_mult_217_n1728), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1729), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1840)
         );
  AOI221_X1 DP_mult_217_U1471 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[21]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[20]), .A(DP_mult_217_n1840), 
        .ZN(DP_mult_217_n1839) );
  XNOR2_X1 DP_mult_217_U1470 ( .A(DP_coeff_pipe01[11]), .B(DP_mult_217_n1839), 
        .ZN(DP_mult_217_n831) );
  OAI22_X1 DP_mult_217_U1469 ( .A1(DP_mult_217_n1724), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1725), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1838)
         );
  AOI221_X1 DP_mult_217_U1468 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[20]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[19]), .A(DP_mult_217_n1838), 
        .ZN(DP_mult_217_n1837) );
  XNOR2_X1 DP_mult_217_U1467 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1837), 
        .ZN(DP_mult_217_n832) );
  OAI22_X1 DP_mult_217_U1466 ( .A1(DP_mult_217_n1720), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1721), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1836)
         );
  AOI221_X1 DP_mult_217_U1465 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[19]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[18]), .A(DP_mult_217_n1836), 
        .ZN(DP_mult_217_n1835) );
  XNOR2_X1 DP_mult_217_U1464 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1835), 
        .ZN(DP_mult_217_n833) );
  OAI22_X1 DP_mult_217_U1463 ( .A1(DP_mult_217_n1716), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1717), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1834)
         );
  AOI221_X1 DP_mult_217_U1462 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[18]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[17]), .A(DP_mult_217_n1834), 
        .ZN(DP_mult_217_n1833) );
  XNOR2_X1 DP_mult_217_U1461 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1833), 
        .ZN(DP_mult_217_n834) );
  OAI22_X1 DP_mult_217_U1460 ( .A1(DP_mult_217_n1712), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1713), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1832)
         );
  AOI221_X1 DP_mult_217_U1459 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[17]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[16]), .A(DP_mult_217_n1832), 
        .ZN(DP_mult_217_n1831) );
  XNOR2_X1 DP_mult_217_U1458 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1831), 
        .ZN(DP_mult_217_n835) );
  OAI22_X1 DP_mult_217_U1457 ( .A1(DP_mult_217_n1708), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1709), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1830)
         );
  AOI221_X1 DP_mult_217_U1456 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[16]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[15]), .A(DP_mult_217_n1830), 
        .ZN(DP_mult_217_n1829) );
  XNOR2_X1 DP_mult_217_U1455 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1829), 
        .ZN(DP_mult_217_n836) );
  OAI22_X1 DP_mult_217_U1454 ( .A1(DP_mult_217_n1704), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1705), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1828)
         );
  AOI221_X1 DP_mult_217_U1453 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[15]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[14]), .A(DP_mult_217_n1828), 
        .ZN(DP_mult_217_n1827) );
  XNOR2_X1 DP_mult_217_U1452 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1827), 
        .ZN(DP_mult_217_n837) );
  OAI22_X1 DP_mult_217_U1451 ( .A1(DP_mult_217_n1700), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1701), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1826)
         );
  AOI221_X1 DP_mult_217_U1450 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[14]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[13]), .A(DP_mult_217_n1826), 
        .ZN(DP_mult_217_n1825) );
  XNOR2_X1 DP_mult_217_U1449 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1825), 
        .ZN(DP_mult_217_n838) );
  OAI22_X1 DP_mult_217_U1448 ( .A1(DP_mult_217_n1696), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1697), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1824)
         );
  AOI221_X1 DP_mult_217_U1447 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[13]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[12]), .A(DP_mult_217_n1824), 
        .ZN(DP_mult_217_n1823) );
  XNOR2_X1 DP_mult_217_U1446 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1823), 
        .ZN(DP_mult_217_n839) );
  OAI22_X1 DP_mult_217_U1445 ( .A1(DP_mult_217_n1692), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1693), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1822)
         );
  AOI221_X1 DP_mult_217_U1444 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[12]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[11]), .A(DP_mult_217_n1822), 
        .ZN(DP_mult_217_n1821) );
  XNOR2_X1 DP_mult_217_U1443 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1821), 
        .ZN(DP_mult_217_n840) );
  OAI22_X1 DP_mult_217_U1442 ( .A1(DP_mult_217_n1688), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1689), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1820)
         );
  AOI221_X1 DP_mult_217_U1441 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[11]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[10]), .A(DP_mult_217_n1820), 
        .ZN(DP_mult_217_n1819) );
  XNOR2_X1 DP_mult_217_U1440 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1819), 
        .ZN(DP_mult_217_n841) );
  OAI22_X1 DP_mult_217_U1439 ( .A1(DP_mult_217_n1684), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1685), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1818)
         );
  AOI221_X1 DP_mult_217_U1438 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[10]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[9]), .A(DP_mult_217_n1818), .ZN(
        DP_mult_217_n1817) );
  XNOR2_X1 DP_mult_217_U1437 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1817), 
        .ZN(DP_mult_217_n842) );
  OAI22_X1 DP_mult_217_U1436 ( .A1(DP_mult_217_n1680), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1681), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1816)
         );
  AOI221_X1 DP_mult_217_U1435 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[9]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[8]), .A(DP_mult_217_n1816), .ZN(
        DP_mult_217_n1815) );
  XNOR2_X1 DP_mult_217_U1434 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1815), 
        .ZN(DP_mult_217_n843) );
  OAI22_X1 DP_mult_217_U1433 ( .A1(DP_mult_217_n1676), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1677), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1814)
         );
  AOI221_X1 DP_mult_217_U1432 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[8]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[7]), .A(DP_mult_217_n1814), .ZN(
        DP_mult_217_n1813) );
  XNOR2_X1 DP_mult_217_U1431 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1813), 
        .ZN(DP_mult_217_n844) );
  OAI22_X1 DP_mult_217_U1430 ( .A1(DP_mult_217_n1672), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1673), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1812)
         );
  AOI221_X1 DP_mult_217_U1429 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[7]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[6]), .A(DP_mult_217_n1812), .ZN(
        DP_mult_217_n1811) );
  XNOR2_X1 DP_mult_217_U1428 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1811), 
        .ZN(DP_mult_217_n845) );
  OAI22_X1 DP_mult_217_U1427 ( .A1(DP_mult_217_n1668), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1669), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1810)
         );
  AOI221_X1 DP_mult_217_U1426 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[6]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[5]), .A(DP_mult_217_n1810), .ZN(
        DP_mult_217_n1809) );
  XNOR2_X1 DP_mult_217_U1425 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1809), 
        .ZN(DP_mult_217_n846) );
  OAI22_X1 DP_mult_217_U1424 ( .A1(DP_mult_217_n1664), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1665), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1808)
         );
  AOI221_X1 DP_mult_217_U1423 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[5]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[4]), .A(DP_mult_217_n1808), .ZN(
        DP_mult_217_n1807) );
  XNOR2_X1 DP_mult_217_U1422 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1807), 
        .ZN(DP_mult_217_n847) );
  OAI22_X1 DP_mult_217_U1421 ( .A1(DP_mult_217_n1660), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1661), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1806)
         );
  AOI221_X1 DP_mult_217_U1420 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[4]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[3]), .A(DP_mult_217_n1806), .ZN(
        DP_mult_217_n1805) );
  XNOR2_X1 DP_mult_217_U1419 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1805), 
        .ZN(DP_mult_217_n848) );
  OAI22_X1 DP_mult_217_U1418 ( .A1(DP_mult_217_n1657), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1649), .B2(DP_mult_217_n1582), .ZN(DP_mult_217_n1804)
         );
  AOI221_X1 DP_mult_217_U1417 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[3]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[2]), .A(DP_mult_217_n1804), .ZN(
        DP_mult_217_n1803) );
  XNOR2_X1 DP_mult_217_U1416 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1803), 
        .ZN(DP_mult_217_n849) );
  OAI22_X1 DP_mult_217_U1415 ( .A1(DP_mult_217_n1653), .A2(DP_mult_217_n1578), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1581), .ZN(DP_mult_217_n1801)
         );
  AOI221_X1 DP_mult_217_U1414 ( .B1(DP_mult_217_n1579), .B2(DP_pipe01[2]), 
        .C1(DP_mult_217_n1580), .C2(DP_pipe01[1]), .A(DP_mult_217_n1801), .ZN(
        DP_mult_217_n1800) );
  XNOR2_X1 DP_mult_217_U1413 ( .A(DP_mult_217_n1602), .B(DP_mult_217_n1800), 
        .ZN(DP_mult_217_n850) );
  OAI222_X1 DP_mult_217_U1412 ( .A1(DP_mult_217_n1649), .A2(DP_mult_217_n1540), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1533), .C1(DP_mult_217_n1650), 
        .C2(DP_mult_217_n1578), .ZN(DP_mult_217_n1799) );
  XNOR2_X1 DP_mult_217_U1411 ( .A(DP_mult_217_n1799), .B(DP_mult_217_n1603), 
        .ZN(DP_mult_217_n851) );
  OAI22_X1 DP_mult_217_U1410 ( .A1(DP_mult_217_n1565), .A2(DP_mult_217_n1540), 
        .B1(DP_mult_217_n1565), .B2(DP_mult_217_n1578), .ZN(DP_mult_217_n1798)
         );
  XNOR2_X1 DP_mult_217_U1409 ( .A(DP_mult_217_n1798), .B(DP_mult_217_n1603), 
        .ZN(DP_mult_217_n852) );
  XOR2_X1 DP_mult_217_U1408 ( .A(DP_coeff_pipe01[6]), .B(DP_mult_217_n1599), 
        .Z(DP_mult_217_n1797) );
  XNOR2_X1 DP_mult_217_U1407 ( .A(DP_coeff_pipe01[7]), .B(DP_mult_217_n1601), 
        .ZN(DP_mult_217_n1796) );
  XNOR2_X1 DP_mult_217_U1406 ( .A(DP_coeff_pipe01[6]), .B(DP_coeff_pipe01[7]), 
        .ZN(DP_mult_217_n1795) );
  NAND3_X1 DP_mult_217_U1405 ( .A1(DP_mult_217_n1797), .A2(DP_mult_217_n1796), 
        .A3(DP_mult_217_n1795), .ZN(DP_mult_217_n1747) );
  INV_X1 DP_mult_217_U1404 ( .A(DP_mult_217_n1797), .ZN(DP_mult_217_n1794) );
  OAI21_X1 DP_mult_217_U1403 ( .B1(DP_mult_217_n1574), .B2(DP_mult_217_n1575), 
        .A(DP_mult_217_n1615), .ZN(DP_mult_217_n1793) );
  OAI221_X1 DP_mult_217_U1402 ( .B1(DP_mult_217_n1618), .B2(DP_mult_217_n1577), 
        .C1(DP_mult_217_n1617), .C2(DP_mult_217_n1573), .A(DP_mult_217_n1793), 
        .ZN(DP_mult_217_n1792) );
  XNOR2_X1 DP_mult_217_U1401 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1792), 
        .ZN(DP_mult_217_n853) );
  OAI22_X1 DP_mult_217_U1400 ( .A1(DP_mult_217_n1633), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1634), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1791)
         );
  AOI221_X1 DP_mult_217_U1399 ( .B1(DP_mult_217_n1574), .B2(DP_mult_217_n1614), 
        .C1(DP_mult_217_n1575), .C2(DP_mult_217_n1615), .A(DP_mult_217_n1791), 
        .ZN(DP_mult_217_n1790) );
  XNOR2_X1 DP_mult_217_U1398 ( .A(DP_coeff_pipe01[8]), .B(DP_mult_217_n1790), 
        .ZN(DP_mult_217_n854) );
  OAI22_X1 DP_mult_217_U1397 ( .A1(DP_mult_217_n1617), .A2(DP_mult_217_n1534), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1789)
         );
  AOI221_X1 DP_mult_217_U1396 ( .B1(DP_mult_217_n1575), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1535), .C2(DP_mult_217_n1375), .A(DP_mult_217_n1789), 
        .ZN(DP_mult_217_n1788) );
  XNOR2_X1 DP_mult_217_U1395 ( .A(DP_coeff_pipe01[8]), .B(DP_mult_217_n1788), 
        .ZN(DP_mult_217_n855) );
  OAI22_X1 DP_mult_217_U1394 ( .A1(DP_mult_217_n1640), .A2(DP_mult_217_n1577), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1536), .ZN(DP_mult_217_n1787)
         );
  AOI221_X1 DP_mult_217_U1393 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1535), .C2(DP_mult_217_n1376), .A(DP_mult_217_n1787), 
        .ZN(DP_mult_217_n1786) );
  XNOR2_X1 DP_mult_217_U1392 ( .A(DP_coeff_pipe01[8]), .B(DP_mult_217_n1786), 
        .ZN(DP_mult_217_n856) );
  OAI22_X1 DP_mult_217_U1391 ( .A1(DP_mult_217_n1728), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1729), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1785)
         );
  AOI221_X1 DP_mult_217_U1390 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[21]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[20]), .A(DP_mult_217_n1785), 
        .ZN(DP_mult_217_n1784) );
  XNOR2_X1 DP_mult_217_U1389 ( .A(DP_coeff_pipe01[8]), .B(DP_mult_217_n1784), 
        .ZN(DP_mult_217_n857) );
  OAI22_X1 DP_mult_217_U1388 ( .A1(DP_mult_217_n1724), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1725), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1783)
         );
  AOI221_X1 DP_mult_217_U1387 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[20]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[19]), .A(DP_mult_217_n1783), 
        .ZN(DP_mult_217_n1782) );
  XNOR2_X1 DP_mult_217_U1386 ( .A(DP_coeff_pipe01[8]), .B(DP_mult_217_n1782), 
        .ZN(DP_mult_217_n858) );
  OAI22_X1 DP_mult_217_U1385 ( .A1(DP_mult_217_n1720), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1721), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1781)
         );
  AOI221_X1 DP_mult_217_U1384 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[19]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[18]), .A(DP_mult_217_n1781), 
        .ZN(DP_mult_217_n1780) );
  XNOR2_X1 DP_mult_217_U1383 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1780), 
        .ZN(DP_mult_217_n859) );
  OAI22_X1 DP_mult_217_U1382 ( .A1(DP_mult_217_n1716), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1717), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1779)
         );
  AOI221_X1 DP_mult_217_U1381 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[18]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[17]), .A(DP_mult_217_n1779), 
        .ZN(DP_mult_217_n1778) );
  XNOR2_X1 DP_mult_217_U1380 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1778), 
        .ZN(DP_mult_217_n860) );
  OAI22_X1 DP_mult_217_U1379 ( .A1(DP_mult_217_n1712), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1713), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1777)
         );
  AOI221_X1 DP_mult_217_U1378 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[17]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[16]), .A(DP_mult_217_n1777), 
        .ZN(DP_mult_217_n1776) );
  XNOR2_X1 DP_mult_217_U1377 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1776), 
        .ZN(DP_mult_217_n861) );
  OAI22_X1 DP_mult_217_U1376 ( .A1(DP_mult_217_n1708), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1709), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1775)
         );
  AOI221_X1 DP_mult_217_U1375 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[16]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[15]), .A(DP_mult_217_n1775), 
        .ZN(DP_mult_217_n1774) );
  XNOR2_X1 DP_mult_217_U1374 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1774), 
        .ZN(DP_mult_217_n862) );
  OAI22_X1 DP_mult_217_U1373 ( .A1(DP_mult_217_n1704), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1705), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1773)
         );
  AOI221_X1 DP_mult_217_U1372 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[15]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[14]), .A(DP_mult_217_n1773), 
        .ZN(DP_mult_217_n1772) );
  XNOR2_X1 DP_mult_217_U1371 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1772), 
        .ZN(DP_mult_217_n863) );
  OAI22_X1 DP_mult_217_U1370 ( .A1(DP_mult_217_n1700), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1701), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1771)
         );
  AOI221_X1 DP_mult_217_U1369 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[14]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[13]), .A(DP_mult_217_n1771), 
        .ZN(DP_mult_217_n1770) );
  XNOR2_X1 DP_mult_217_U1368 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1770), 
        .ZN(DP_mult_217_n864) );
  OAI22_X1 DP_mult_217_U1367 ( .A1(DP_mult_217_n1696), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1697), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1769)
         );
  AOI221_X1 DP_mult_217_U1366 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[13]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[12]), .A(DP_mult_217_n1769), 
        .ZN(DP_mult_217_n1768) );
  XNOR2_X1 DP_mult_217_U1365 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1768), 
        .ZN(DP_mult_217_n865) );
  OAI22_X1 DP_mult_217_U1364 ( .A1(DP_mult_217_n1692), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1693), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1767)
         );
  AOI221_X1 DP_mult_217_U1363 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[12]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[11]), .A(DP_mult_217_n1767), 
        .ZN(DP_mult_217_n1766) );
  XNOR2_X1 DP_mult_217_U1362 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1766), 
        .ZN(DP_mult_217_n866) );
  OAI22_X1 DP_mult_217_U1361 ( .A1(DP_mult_217_n1688), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1689), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1765)
         );
  AOI221_X1 DP_mult_217_U1360 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[11]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[10]), .A(DP_mult_217_n1765), 
        .ZN(DP_mult_217_n1764) );
  XNOR2_X1 DP_mult_217_U1359 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1764), 
        .ZN(DP_mult_217_n867) );
  OAI22_X1 DP_mult_217_U1358 ( .A1(DP_mult_217_n1684), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1685), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1763)
         );
  AOI221_X1 DP_mult_217_U1357 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[10]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[9]), .A(DP_mult_217_n1763), .ZN(
        DP_mult_217_n1762) );
  XNOR2_X1 DP_mult_217_U1356 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1762), 
        .ZN(DP_mult_217_n868) );
  OAI22_X1 DP_mult_217_U1355 ( .A1(DP_mult_217_n1680), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1681), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1761)
         );
  AOI221_X1 DP_mult_217_U1354 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[9]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[8]), .A(DP_mult_217_n1761), .ZN(
        DP_mult_217_n1760) );
  XNOR2_X1 DP_mult_217_U1353 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1760), 
        .ZN(DP_mult_217_n869) );
  OAI22_X1 DP_mult_217_U1352 ( .A1(DP_mult_217_n1676), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1677), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1759)
         );
  AOI221_X1 DP_mult_217_U1351 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[8]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[7]), .A(DP_mult_217_n1759), .ZN(
        DP_mult_217_n1758) );
  XNOR2_X1 DP_mult_217_U1350 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1758), 
        .ZN(DP_mult_217_n870) );
  OAI22_X1 DP_mult_217_U1349 ( .A1(DP_mult_217_n1672), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1673), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1757)
         );
  AOI221_X1 DP_mult_217_U1348 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[7]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[6]), .A(DP_mult_217_n1757), .ZN(
        DP_mult_217_n1756) );
  XNOR2_X1 DP_mult_217_U1347 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1756), 
        .ZN(DP_mult_217_n871) );
  OAI22_X1 DP_mult_217_U1346 ( .A1(DP_mult_217_n1668), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1669), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1755)
         );
  AOI221_X1 DP_mult_217_U1345 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[6]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[5]), .A(DP_mult_217_n1755), .ZN(
        DP_mult_217_n1754) );
  XNOR2_X1 DP_mult_217_U1344 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1754), 
        .ZN(DP_mult_217_n872) );
  OAI22_X1 DP_mult_217_U1343 ( .A1(DP_mult_217_n1664), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1665), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1753)
         );
  AOI221_X1 DP_mult_217_U1342 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[5]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[4]), .A(DP_mult_217_n1753), .ZN(
        DP_mult_217_n1752) );
  XNOR2_X1 DP_mult_217_U1341 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1752), 
        .ZN(DP_mult_217_n873) );
  OAI22_X1 DP_mult_217_U1340 ( .A1(DP_mult_217_n1660), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1661), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1751)
         );
  AOI221_X1 DP_mult_217_U1339 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[4]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[3]), .A(DP_mult_217_n1751), .ZN(
        DP_mult_217_n1750) );
  XNOR2_X1 DP_mult_217_U1338 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1750), 
        .ZN(DP_mult_217_n874) );
  OAI22_X1 DP_mult_217_U1337 ( .A1(DP_mult_217_n1657), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1649), .B2(DP_mult_217_n1577), .ZN(DP_mult_217_n1749)
         );
  AOI221_X1 DP_mult_217_U1336 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[3]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[2]), .A(DP_mult_217_n1749), .ZN(
        DP_mult_217_n1748) );
  XNOR2_X1 DP_mult_217_U1335 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1748), 
        .ZN(DP_mult_217_n875) );
  OAI22_X1 DP_mult_217_U1334 ( .A1(DP_mult_217_n1653), .A2(DP_mult_217_n1573), 
        .B1(DP_mult_217_n1565), .B2(DP_mult_217_n1576), .ZN(DP_mult_217_n1746)
         );
  AOI221_X1 DP_mult_217_U1333 ( .B1(DP_mult_217_n1574), .B2(DP_pipe01[2]), 
        .C1(DP_mult_217_n1575), .C2(DP_pipe01[1]), .A(DP_mult_217_n1746), .ZN(
        DP_mult_217_n1745) );
  XNOR2_X1 DP_mult_217_U1332 ( .A(DP_mult_217_n1600), .B(DP_mult_217_n1745), 
        .ZN(DP_mult_217_n876) );
  OAI222_X1 DP_mult_217_U1331 ( .A1(DP_mult_217_n1649), .A2(DP_mult_217_n1534), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1536), .C1(DP_mult_217_n1650), 
        .C2(DP_mult_217_n1573), .ZN(DP_mult_217_n1744) );
  XNOR2_X1 DP_mult_217_U1330 ( .A(DP_mult_217_n1744), .B(DP_mult_217_n1601), 
        .ZN(DP_mult_217_n877) );
  OAI22_X1 DP_mult_217_U1329 ( .A1(DP_mult_217_n1565), .A2(DP_mult_217_n1534), 
        .B1(DP_mult_217_n1565), .B2(DP_mult_217_n1573), .ZN(DP_mult_217_n1743)
         );
  XNOR2_X1 DP_mult_217_U1328 ( .A(DP_mult_217_n1743), .B(DP_mult_217_n1601), 
        .ZN(DP_mult_217_n878) );
  XOR2_X1 DP_mult_217_U1327 ( .A(DP_coeff_pipe01[3]), .B(DP_mult_217_n1742), 
        .Z(DP_mult_217_n1741) );
  XNOR2_X1 DP_mult_217_U1326 ( .A(DP_coeff_pipe01[4]), .B(DP_mult_217_n1599), 
        .ZN(DP_mult_217_n1740) );
  XNOR2_X1 DP_mult_217_U1325 ( .A(DP_coeff_pipe01[3]), .B(DP_coeff_pipe01[4]), 
        .ZN(DP_mult_217_n1739) );
  NAND3_X1 DP_mult_217_U1324 ( .A1(DP_mult_217_n1741), .A2(DP_mult_217_n1740), 
        .A3(DP_mult_217_n1739), .ZN(DP_mult_217_n1654) );
  INV_X1 DP_mult_217_U1323 ( .A(DP_mult_217_n1741), .ZN(DP_mult_217_n1738) );
  OAI21_X1 DP_mult_217_U1322 ( .B1(DP_mult_217_n1569), .B2(DP_mult_217_n1570), 
        .A(DP_mult_217_n1615), .ZN(DP_mult_217_n1737) );
  OAI221_X1 DP_mult_217_U1321 ( .B1(DP_mult_217_n1618), .B2(DP_mult_217_n1572), 
        .C1(DP_mult_217_n1618), .C2(DP_mult_217_n1568), .A(DP_mult_217_n1737), 
        .ZN(DP_mult_217_n1736) );
  XNOR2_X1 DP_mult_217_U1320 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1736), 
        .ZN(DP_mult_217_n879) );
  OAI22_X1 DP_mult_217_U1319 ( .A1(DP_mult_217_n1633), .A2(DP_mult_217_n1568), 
        .B1(DP_mult_217_n1634), .B2(DP_mult_217_n1572), .ZN(DP_mult_217_n1735)
         );
  AOI221_X1 DP_mult_217_U1318 ( .B1(DP_mult_217_n1569), .B2(DP_mult_217_n1614), 
        .C1(DP_mult_217_n1570), .C2(DP_mult_217_n1615), .A(DP_mult_217_n1735), 
        .ZN(DP_mult_217_n1734) );
  XNOR2_X1 DP_mult_217_U1317 ( .A(DP_coeff_pipe01[5]), .B(DP_mult_217_n1734), 
        .ZN(DP_mult_217_n880) );
  OAI22_X1 DP_mult_217_U1316 ( .A1(DP_mult_217_n1616), .A2(DP_mult_217_n1538), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1572), .ZN(DP_mult_217_n1733)
         );
  AOI221_X1 DP_mult_217_U1315 ( .B1(DP_mult_217_n1570), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1537), .C2(DP_mult_217_n1375), .A(DP_mult_217_n1733), 
        .ZN(DP_mult_217_n1732) );
  XNOR2_X1 DP_mult_217_U1314 ( .A(DP_coeff_pipe01[5]), .B(DP_mult_217_n1732), 
        .ZN(DP_mult_217_n881) );
  OAI22_X1 DP_mult_217_U1313 ( .A1(DP_mult_217_n1640), .A2(DP_mult_217_n1572), 
        .B1(DP_mult_217_n1643), .B2(DP_mult_217_n1539), .ZN(DP_mult_217_n1731)
         );
  AOI221_X1 DP_mult_217_U1312 ( .B1(DP_mult_217_n1569), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1537), .C2(DP_mult_217_n1376), .A(DP_mult_217_n1731), 
        .ZN(DP_mult_217_n1730) );
  XNOR2_X1 DP_mult_217_U1311 ( .A(DP_coeff_pipe01[5]), .B(DP_mult_217_n1730), 
        .ZN(DP_mult_217_n882) );
  OAI22_X1 DP_mult_217_U1310 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1728), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1729), .ZN(DP_mult_217_n1727)
         );
  AOI221_X1 DP_mult_217_U1309 ( .B1(DP_mult_217_n1569), .B2(DP_pipe01[21]), 
        .C1(DP_mult_217_n1570), .C2(DP_pipe01[20]), .A(DP_mult_217_n1727), 
        .ZN(DP_mult_217_n1726) );
  XNOR2_X1 DP_mult_217_U1308 ( .A(DP_coeff_pipe01[5]), .B(DP_mult_217_n1726), 
        .ZN(DP_mult_217_n883) );
  OAI22_X1 DP_mult_217_U1307 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1724), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1725), .ZN(DP_mult_217_n1723)
         );
  AOI221_X1 DP_mult_217_U1306 ( .B1(DP_mult_217_n1569), .B2(DP_pipe01[20]), 
        .C1(DP_pipe01[19]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1723), 
        .ZN(DP_mult_217_n1722) );
  XNOR2_X1 DP_mult_217_U1305 ( .A(DP_coeff_pipe01[5]), .B(DP_mult_217_n1722), 
        .ZN(DP_mult_217_n884) );
  OAI22_X1 DP_mult_217_U1304 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1720), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1721), .ZN(DP_mult_217_n1719)
         );
  AOI221_X1 DP_mult_217_U1303 ( .B1(DP_pipe01[19]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[18]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1719), 
        .ZN(DP_mult_217_n1718) );
  XNOR2_X1 DP_mult_217_U1302 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1718), 
        .ZN(DP_mult_217_n885) );
  OAI22_X1 DP_mult_217_U1301 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1716), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1717), .ZN(DP_mult_217_n1715)
         );
  AOI221_X1 DP_mult_217_U1300 ( .B1(DP_pipe01[18]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[17]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1715), 
        .ZN(DP_mult_217_n1714) );
  XNOR2_X1 DP_mult_217_U1299 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1714), 
        .ZN(DP_mult_217_n886) );
  OAI22_X1 DP_mult_217_U1298 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1712), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1713), .ZN(DP_mult_217_n1711)
         );
  AOI221_X1 DP_mult_217_U1297 ( .B1(DP_pipe01[17]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[16]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1711), 
        .ZN(DP_mult_217_n1710) );
  XNOR2_X1 DP_mult_217_U1296 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1710), 
        .ZN(DP_mult_217_n887) );
  OAI22_X1 DP_mult_217_U1295 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1708), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1709), .ZN(DP_mult_217_n1707)
         );
  AOI221_X1 DP_mult_217_U1294 ( .B1(DP_pipe01[16]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[15]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1707), 
        .ZN(DP_mult_217_n1706) );
  XNOR2_X1 DP_mult_217_U1293 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1706), 
        .ZN(DP_mult_217_n888) );
  OAI22_X1 DP_mult_217_U1292 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1704), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1705), .ZN(DP_mult_217_n1703)
         );
  AOI221_X1 DP_mult_217_U1291 ( .B1(DP_pipe01[15]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[14]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1703), 
        .ZN(DP_mult_217_n1702) );
  XNOR2_X1 DP_mult_217_U1290 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1702), 
        .ZN(DP_mult_217_n889) );
  OAI22_X1 DP_mult_217_U1289 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1700), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1701), .ZN(DP_mult_217_n1699)
         );
  AOI221_X1 DP_mult_217_U1288 ( .B1(DP_pipe01[14]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[13]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1699), 
        .ZN(DP_mult_217_n1698) );
  XNOR2_X1 DP_mult_217_U1287 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1698), 
        .ZN(DP_mult_217_n890) );
  OAI22_X1 DP_mult_217_U1286 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1696), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1697), .ZN(DP_mult_217_n1695)
         );
  AOI221_X1 DP_mult_217_U1285 ( .B1(DP_pipe01[13]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[12]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1695), 
        .ZN(DP_mult_217_n1694) );
  XNOR2_X1 DP_mult_217_U1284 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1694), 
        .ZN(DP_mult_217_n891) );
  OAI22_X1 DP_mult_217_U1283 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1692), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1693), .ZN(DP_mult_217_n1691)
         );
  AOI221_X1 DP_mult_217_U1282 ( .B1(DP_pipe01[12]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[11]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1691), 
        .ZN(DP_mult_217_n1690) );
  XNOR2_X1 DP_mult_217_U1281 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1690), 
        .ZN(DP_mult_217_n892) );
  OAI22_X1 DP_mult_217_U1280 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1688), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1689), .ZN(DP_mult_217_n1687)
         );
  AOI221_X1 DP_mult_217_U1279 ( .B1(DP_pipe01[11]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[10]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1687), 
        .ZN(DP_mult_217_n1686) );
  XNOR2_X1 DP_mult_217_U1278 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1686), 
        .ZN(DP_mult_217_n893) );
  OAI22_X1 DP_mult_217_U1277 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1684), 
        .B1(DP_mult_217_n1572), .B2(DP_mult_217_n1685), .ZN(DP_mult_217_n1683)
         );
  AOI221_X1 DP_mult_217_U1276 ( .B1(DP_pipe01[10]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[9]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1683), .ZN(
        DP_mult_217_n1682) );
  XNOR2_X1 DP_mult_217_U1275 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1682), 
        .ZN(DP_mult_217_n894) );
  OAI22_X1 DP_mult_217_U1274 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1680), 
        .B1(DP_mult_217_n1572), .B2(DP_mult_217_n1681), .ZN(DP_mult_217_n1679)
         );
  AOI221_X1 DP_mult_217_U1273 ( .B1(DP_pipe01[9]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[8]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1679), .ZN(
        DP_mult_217_n1678) );
  XNOR2_X1 DP_mult_217_U1272 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1678), 
        .ZN(DP_mult_217_n895) );
  OAI22_X1 DP_mult_217_U1271 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1676), 
        .B1(DP_mult_217_n1571), .B2(DP_mult_217_n1677), .ZN(DP_mult_217_n1675)
         );
  AOI221_X1 DP_mult_217_U1270 ( .B1(DP_pipe01[8]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[7]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1675), .ZN(
        DP_mult_217_n1674) );
  XNOR2_X1 DP_mult_217_U1269 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1674), 
        .ZN(DP_mult_217_n896) );
  OAI22_X1 DP_mult_217_U1268 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1672), 
        .B1(DP_mult_217_n1572), .B2(DP_mult_217_n1673), .ZN(DP_mult_217_n1671)
         );
  AOI221_X1 DP_mult_217_U1267 ( .B1(DP_pipe01[7]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[6]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1671), .ZN(
        DP_mult_217_n1670) );
  XNOR2_X1 DP_mult_217_U1266 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1670), 
        .ZN(DP_mult_217_n897) );
  OAI22_X1 DP_mult_217_U1265 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1668), 
        .B1(DP_mult_217_n1572), .B2(DP_mult_217_n1669), .ZN(DP_mult_217_n1667)
         );
  AOI221_X1 DP_mult_217_U1264 ( .B1(DP_pipe01[6]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[5]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1667), .ZN(
        DP_mult_217_n1666) );
  XNOR2_X1 DP_mult_217_U1263 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1666), 
        .ZN(DP_mult_217_n898) );
  OAI22_X1 DP_mult_217_U1262 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1664), 
        .B1(DP_mult_217_n1572), .B2(DP_mult_217_n1665), .ZN(DP_mult_217_n1663)
         );
  AOI221_X1 DP_mult_217_U1261 ( .B1(DP_pipe01[5]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[4]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1663), .ZN(
        DP_mult_217_n1662) );
  XNOR2_X1 DP_mult_217_U1260 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1662), 
        .ZN(DP_mult_217_n899) );
  OAI22_X1 DP_mult_217_U1259 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1660), 
        .B1(DP_mult_217_n1661), .B2(DP_mult_217_n1572), .ZN(DP_mult_217_n1659)
         );
  AOI221_X1 DP_mult_217_U1258 ( .B1(DP_pipe01[4]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[3]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1659), .ZN(
        DP_mult_217_n1658) );
  XNOR2_X1 DP_mult_217_U1257 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1658), 
        .ZN(DP_mult_217_n900) );
  OAI22_X1 DP_mult_217_U1256 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1657), 
        .B1(DP_mult_217_n1649), .B2(DP_mult_217_n1572), .ZN(DP_mult_217_n1656)
         );
  AOI221_X1 DP_mult_217_U1255 ( .B1(DP_pipe01[3]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[2]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1656), .ZN(
        DP_mult_217_n1655) );
  XNOR2_X1 DP_mult_217_U1254 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1655), 
        .ZN(DP_mult_217_n901) );
  OAI22_X1 DP_mult_217_U1253 ( .A1(DP_mult_217_n1568), .A2(DP_mult_217_n1653), 
        .B1(DP_mult_217_n1565), .B2(DP_mult_217_n1572), .ZN(DP_mult_217_n1652)
         );
  AOI221_X1 DP_mult_217_U1252 ( .B1(DP_pipe01[2]), .B2(DP_mult_217_n1569), 
        .C1(DP_pipe01[1]), .C2(DP_mult_217_n1570), .A(DP_mult_217_n1652), .ZN(
        DP_mult_217_n1651) );
  XNOR2_X1 DP_mult_217_U1251 ( .A(DP_mult_217_n1598), .B(DP_mult_217_n1651), 
        .ZN(DP_mult_217_n902) );
  OAI222_X1 DP_mult_217_U1250 ( .A1(DP_mult_217_n1538), .A2(DP_mult_217_n1649), 
        .B1(DP_mult_217_n1566), .B2(DP_mult_217_n1539), .C1(DP_mult_217_n1568), 
        .C2(DP_mult_217_n1650), .ZN(DP_mult_217_n1648) );
  XNOR2_X1 DP_mult_217_U1249 ( .A(DP_mult_217_n1648), .B(DP_mult_217_n1599), 
        .ZN(DP_mult_217_n903) );
  OAI22_X1 DP_mult_217_U1248 ( .A1(DP_mult_217_n1565), .A2(DP_mult_217_n1538), 
        .B1(DP_mult_217_n1568), .B2(DP_mult_217_n1567), .ZN(DP_mult_217_n1646)
         );
  XNOR2_X1 DP_mult_217_U1247 ( .A(DP_mult_217_n1646), .B(DP_mult_217_n1599), 
        .ZN(DP_mult_217_n904) );
  OAI22_X1 DP_mult_217_U1246 ( .A1(DP_mult_217_n1633), .A2(DP_mult_217_n1564), 
        .B1(DP_mult_217_n1634), .B2(DP_mult_217_n1639), .ZN(DP_mult_217_n1645)
         );
  AOI221_X1 DP_mult_217_U1245 ( .B1(DP_mult_217_n1561), .B2(DP_mult_217_n1614), 
        .C1(DP_mult_217_n1563), .C2(DP_mult_217_n1615), .A(DP_mult_217_n1645), 
        .ZN(DP_mult_217_n1644) );
  XNOR2_X1 DP_mult_217_U1244 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n1644), 
        .ZN(DP_mult_217_n906) );
  OAI22_X1 DP_mult_217_U1243 ( .A1(DP_mult_217_n1643), .A2(DP_mult_217_n1639), 
        .B1(DP_mult_217_n1617), .B2(DP_mult_217_n1542), .ZN(DP_mult_217_n1642)
         );
  AOI221_X1 DP_mult_217_U1242 ( .B1(DP_mult_217_n1563), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1554), .C2(DP_mult_217_n1375), .A(DP_mult_217_n1642), 
        .ZN(DP_mult_217_n1641) );
  XNOR2_X1 DP_mult_217_U1241 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n1641), 
        .ZN(DP_mult_217_n907) );
  INV_X1 DP_mult_217_U1240 ( .A(DP_mult_217_n1376), .ZN(DP_mult_217_n1638) );
  OAI22_X1 DP_mult_217_U1239 ( .A1(DP_mult_217_n1564), .A2(DP_mult_217_n1638), 
        .B1(DP_mult_217_n1639), .B2(DP_mult_217_n1640), .ZN(DP_mult_217_n1637)
         );
  AOI221_X1 DP_mult_217_U1238 ( .B1(DP_mult_217_n1561), .B2(DP_pipe01[22]), 
        .C1(DP_mult_217_n1563), .C2(DP_pipe01[21]), .A(DP_mult_217_n1637), 
        .ZN(DP_mult_217_n1635) );
  XNOR2_X1 DP_mult_217_U1237 ( .A(DP_coeff_pipe01[2]), .B(DP_mult_217_n1635), 
        .ZN(DP_mult_217_n908) );
  OAI22_X1 DP_mult_217_U1236 ( .A1(DP_mult_217_n1558), .A2(DP_mult_217_n1633), 
        .B1(DP_mult_217_n1557), .B2(DP_mult_217_n1634), .ZN(DP_mult_217_n1632)
         );
  AOI221_X1 DP_mult_217_U1235 ( .B1(DP_mult_217_n1613), .B2(DP_mult_217_n1559), 
        .C1(DP_mult_217_n1560), .C2(DP_mult_217_n1615), .A(DP_mult_217_n1632), 
        .ZN(DP_mult_217_n1631) );
  XOR2_X1 DP_mult_217_U1234 ( .A(DP_coeff_pipe01[23]), .B(DP_mult_217_n1631), 
        .Z(DP_mult_217_n1625) );
  INV_X1 DP_mult_217_U1233 ( .A(DP_mult_217_n1625), .ZN(DP_mult_217_n1621) );
  OAI21_X1 DP_mult_217_U1232 ( .B1(DP_mult_217_n1559), .B2(DP_mult_217_n1560), 
        .A(DP_mult_217_n1615), .ZN(DP_mult_217_n1630) );
  OAI221_X1 DP_mult_217_U1231 ( .B1(DP_mult_217_n1617), .B2(DP_mult_217_n1557), 
        .C1(DP_mult_217_n1617), .C2(DP_mult_217_n1558), .A(DP_mult_217_n1630), 
        .ZN(DP_mult_217_n1628) );
  XOR2_X1 DP_mult_217_U1230 ( .A(DP_mult_217_n1628), .B(DP_mult_217_n1611), 
        .Z(DP_mult_217_n1622) );
  AOI222_X1 DP_mult_217_U1229 ( .A1(DP_mult_217_n1627), .A2(DP_mult_217_n303), 
        .B1(DP_mult_217_n1625), .B2(DP_mult_217_n303), .C1(DP_mult_217_n1627), 
        .C2(DP_mult_217_n1625), .ZN(DP_mult_217_n1624) );
  INV_X1 DP_mult_217_U1228 ( .A(DP_mult_217_n1622), .ZN(DP_mult_217_n1626) );
  OAI22_X1 DP_mult_217_U1227 ( .A1(DP_mult_217_n1624), .A2(DP_mult_217_n1625), 
        .B1(DP_mult_217_n1624), .B2(DP_mult_217_n1626), .ZN(DP_mult_217_n1623)
         );
  AOI21_X1 DP_mult_217_U1226 ( .B1(DP_mult_217_n1621), .B2(DP_mult_217_n1622), 
        .A(DP_mult_217_n1623), .ZN(DP_pipe0_coeff_pipe01[23]) );
  INV_X1 DP_mult_217_U1225 ( .A(DP_mult_217_n1614), .ZN(DP_mult_217_n1620) );
  INV_X1 DP_mult_217_U1224 ( .A(DP_mult_217_n1613), .ZN(DP_mult_217_n1619) );
  INV_X1 DP_mult_217_U1223 ( .A(DP_mult_217_n1613), .ZN(DP_mult_217_n1618) );
  INV_X1 DP_mult_217_U1222 ( .A(DP_mult_217_n1612), .ZN(DP_mult_217_n1617) );
  INV_X1 DP_mult_217_U1221 ( .A(DP_mult_217_n1612), .ZN(DP_mult_217_n1616) );
  CLKBUF_X1 DP_mult_217_U1220 ( .A(DP_pipe01[23]), .Z(DP_mult_217_n1614) );
  CLKBUF_X1 DP_mult_217_U1219 ( .A(DP_pipe01[23]), .Z(DP_mult_217_n1613) );
  CLKBUF_X1 DP_mult_217_U1218 ( .A(DP_pipe01[23]), .Z(DP_mult_217_n1612) );
  INV_X1 DP_mult_217_U1217 ( .A(DP_coeff_pipe01[23]), .ZN(DP_mult_217_n1611)
         );
  BUF_X1 DP_mult_217_U1216 ( .A(DP_mult_217_n1647), .Z(DP_mult_217_n1567) );
  BUF_X1 DP_mult_217_U1215 ( .A(DP_mult_217_n1647), .Z(DP_mult_217_n1566) );
  BUF_X1 DP_mult_217_U1214 ( .A(DP_mult_217_n1647), .Z(DP_mult_217_n1565) );
  BUF_X1 DP_mult_217_U1213 ( .A(DP_coeff_pipe01[20]), .Z(DP_mult_217_n1609) );
  INV_X1 DP_mult_217_U1212 ( .A(DP_coeff_pipe01[17]), .ZN(DP_mult_217_n1607)
         );
  INV_X1 DP_mult_217_U1211 ( .A(DP_coeff_pipe01[14]), .ZN(DP_mult_217_n1605)
         );
  INV_X1 DP_mult_217_U1210 ( .A(DP_coeff_pipe01[11]), .ZN(DP_mult_217_n1603)
         );
  BUF_X1 DP_mult_217_U1209 ( .A(DP_coeff_pipe01[20]), .Z(DP_mult_217_n1608) );
  INV_X1 DP_mult_217_U1208 ( .A(DP_mult_217_n1611), .ZN(DP_mult_217_n1610) );
  INV_X1 DP_mult_217_U1207 ( .A(DP_mult_217_n1616), .ZN(DP_mult_217_n1615) );
  OR2_X1 DP_mult_217_U1206 ( .A1(DP_mult_217_n1904), .A2(DP_mult_217_n1905), 
        .ZN(DP_mult_217_n1555) );
  AND2_X1 DP_mult_217_U1205 ( .A1(DP_coeff_pipe01[0]), .A2(DP_mult_217_n2157), 
        .ZN(DP_mult_217_n1554) );
  INV_X1 DP_mult_217_U1204 ( .A(DP_mult_217_n1603), .ZN(DP_mult_217_n1602) );
  AND2_X1 DP_mult_217_U1203 ( .A1(DP_mult_217_n2070), .A2(DP_mult_217_n2068), 
        .ZN(DP_mult_217_n1553) );
  OR2_X1 DP_mult_217_U1202 ( .A1(DP_mult_217_n2014), .A2(DP_mult_217_n2015), 
        .ZN(DP_mult_217_n1552) );
  OR2_X1 DP_mult_217_U1201 ( .A1(DP_mult_217_n1959), .A2(DP_mult_217_n1960), 
        .ZN(DP_mult_217_n1551) );
  OR2_X1 DP_mult_217_U1200 ( .A1(DP_mult_217_n2070), .A2(DP_mult_217_n2069), 
        .ZN(DP_mult_217_n1550) );
  AND2_X1 DP_mult_217_U1199 ( .A1(DP_mult_217_n1959), .A2(DP_mult_217_n1961), 
        .ZN(DP_mult_217_n1549) );
  AND2_X1 DP_mult_217_U1198 ( .A1(DP_mult_217_n1904), .A2(DP_mult_217_n1906), 
        .ZN(DP_mult_217_n1548) );
  AND2_X1 DP_mult_217_U1197 ( .A1(DP_mult_217_n2014), .A2(DP_mult_217_n2016), 
        .ZN(DP_mult_217_n1547) );
  OR2_X1 DP_mult_217_U1196 ( .A1(DP_mult_217_n1961), .A2(DP_mult_217_n1962), 
        .ZN(DP_mult_217_n1546) );
  OR2_X1 DP_mult_217_U1195 ( .A1(DP_mult_217_n1906), .A2(DP_mult_217_n1907), 
        .ZN(DP_mult_217_n1545) );
  OR2_X1 DP_mult_217_U1194 ( .A1(DP_mult_217_n2068), .A2(DP_mult_217_n2067), 
        .ZN(DP_mult_217_n1544) );
  OR2_X1 DP_mult_217_U1193 ( .A1(DP_mult_217_n2016), .A2(DP_mult_217_n2017), 
        .ZN(DP_mult_217_n1543) );
  INV_X1 DP_mult_217_U1192 ( .A(DP_mult_217_n1607), .ZN(DP_mult_217_n1606) );
  INV_X1 DP_mult_217_U1191 ( .A(DP_mult_217_n1605), .ZN(DP_mult_217_n1604) );
  BUF_X1 DP_mult_217_U1190 ( .A(DP_mult_217_n1636), .Z(DP_mult_217_n1562) );
  OR2_X1 DP_mult_217_U1189 ( .A1(DP_mult_217_n2158), .A2(DP_mult_217_n2157), 
        .ZN(DP_mult_217_n1542) );
  BUF_X1 DP_mult_217_U1188 ( .A(DP_mult_217_n1629), .Z(DP_mult_217_n1556) );
  BUF_X1 DP_mult_217_U1187 ( .A(DP_mult_217_n1636), .Z(DP_mult_217_n1563) );
  INV_X1 DP_mult_217_U1186 ( .A(DP_mult_217_n1554), .ZN(DP_mult_217_n1564) );
  INV_X1 DP_mult_217_U1185 ( .A(DP_mult_217_n1543), .ZN(DP_mult_217_n1594) );
  INV_X1 DP_mult_217_U1184 ( .A(DP_mult_217_n1546), .ZN(DP_mult_217_n1589) );
  INV_X1 DP_mult_217_U1183 ( .A(DP_mult_217_n1545), .ZN(DP_mult_217_n1584) );
  INV_X1 DP_mult_217_U1182 ( .A(DP_mult_217_n1555), .ZN(DP_mult_217_n1585) );
  NAND3_X1 DP_mult_217_U1181 ( .A1(DP_mult_217_n2157), .A2(DP_mult_217_n2158), 
        .A3(DP_mult_217_n2159), .ZN(DP_mult_217_n1639) );
  AND2_X1 DP_mult_217_U1180 ( .A1(DP_mult_217_n1849), .A2(DP_mult_217_n1851), 
        .ZN(DP_mult_217_n1541) );
  OR2_X1 DP_mult_217_U1179 ( .A1(DP_mult_217_n1851), .A2(DP_mult_217_n1852), 
        .ZN(DP_mult_217_n1540) );
  BUF_X1 DP_mult_217_U1178 ( .A(DP_mult_217_n1967), .Z(DP_mult_217_n1597) );
  BUF_X1 DP_mult_217_U1177 ( .A(DP_mult_217_n1912), .Z(DP_mult_217_n1592) );
  BUF_X1 DP_mult_217_U1176 ( .A(DP_mult_217_n1857), .Z(DP_mult_217_n1587) );
  BUF_X1 DP_mult_217_U1175 ( .A(DP_mult_217_n1912), .Z(DP_mult_217_n1591) );
  BUF_X1 DP_mult_217_U1174 ( .A(DP_mult_217_n1967), .Z(DP_mult_217_n1596) );
  BUF_X1 DP_mult_217_U1173 ( .A(DP_mult_217_n1857), .Z(DP_mult_217_n1586) );
  BUF_X1 DP_mult_217_U1172 ( .A(DP_mult_217_n1629), .Z(DP_mult_217_n1557) );
  INV_X1 DP_mult_217_U1171 ( .A(DP_mult_217_n1547), .ZN(DP_mult_217_n1593) );
  INV_X1 DP_mult_217_U1170 ( .A(DP_mult_217_n1548), .ZN(DP_mult_217_n1583) );
  INV_X1 DP_mult_217_U1169 ( .A(DP_mult_217_n1549), .ZN(DP_mult_217_n1588) );
  INV_X1 DP_mult_217_U1168 ( .A(DP_mult_217_n1544), .ZN(DP_mult_217_n1559) );
  INV_X1 DP_mult_217_U1167 ( .A(DP_mult_217_n1552), .ZN(DP_mult_217_n1595) );
  INV_X1 DP_mult_217_U1166 ( .A(DP_mult_217_n1551), .ZN(DP_mult_217_n1590) );
  INV_X1 DP_mult_217_U1165 ( .A(DP_mult_217_n1553), .ZN(DP_mult_217_n1558) );
  INV_X1 DP_mult_217_U1164 ( .A(DP_mult_217_n1550), .ZN(DP_mult_217_n1560) );
  INV_X1 DP_mult_217_U1163 ( .A(DP_mult_217_n1540), .ZN(DP_mult_217_n1579) );
  INV_X1 DP_mult_217_U1162 ( .A(DP_coeff_pipe01[8]), .ZN(DP_mult_217_n1601) );
  INV_X1 DP_mult_217_U1161 ( .A(DP_coeff_pipe01[5]), .ZN(DP_mult_217_n1599) );
  BUF_X1 DP_mult_217_U1160 ( .A(DP_mult_217_n1802), .Z(DP_mult_217_n1582) );
  BUF_X1 DP_mult_217_U1159 ( .A(DP_mult_217_n1802), .Z(DP_mult_217_n1581) );
  OR2_X1 DP_mult_217_U1158 ( .A1(DP_mult_217_n1738), .A2(DP_mult_217_n1739), 
        .ZN(DP_mult_217_n1539) );
  OR2_X1 DP_mult_217_U1157 ( .A1(DP_mult_217_n1740), .A2(DP_mult_217_n1741), 
        .ZN(DP_mult_217_n1538) );
  INV_X1 DP_mult_217_U1156 ( .A(DP_mult_217_n1542), .ZN(DP_mult_217_n1561) );
  INV_X1 DP_mult_217_U1155 ( .A(DP_mult_217_n1541), .ZN(DP_mult_217_n1578) );
  AND2_X1 DP_mult_217_U1154 ( .A1(DP_mult_217_n1738), .A2(DP_mult_217_n1740), 
        .ZN(DP_mult_217_n1537) );
  BUF_X1 DP_mult_217_U1153 ( .A(DP_mult_217_n1654), .Z(DP_mult_217_n1572) );
  BUF_X1 DP_mult_217_U1152 ( .A(DP_mult_217_n1654), .Z(DP_mult_217_n1571) );
  INV_X1 DP_mult_217_U1151 ( .A(DP_mult_217_n1538), .ZN(DP_mult_217_n1569) );
  INV_X1 DP_mult_217_U1150 ( .A(DP_mult_217_n1539), .ZN(DP_mult_217_n1570) );
  INV_X1 DP_mult_217_U1149 ( .A(DP_mult_217_n1601), .ZN(DP_mult_217_n1600) );
  INV_X1 DP_mult_217_U1148 ( .A(DP_mult_217_n1599), .ZN(DP_mult_217_n1598) );
  OR2_X1 DP_mult_217_U1147 ( .A1(DP_mult_217_n1794), .A2(DP_mult_217_n1795), 
        .ZN(DP_mult_217_n1536) );
  AND2_X1 DP_mult_217_U1146 ( .A1(DP_mult_217_n1794), .A2(DP_mult_217_n1796), 
        .ZN(DP_mult_217_n1535) );
  OR2_X1 DP_mult_217_U1145 ( .A1(DP_mult_217_n1796), .A2(DP_mult_217_n1797), 
        .ZN(DP_mult_217_n1534) );
  INV_X1 DP_mult_217_U1144 ( .A(DP_mult_217_n1537), .ZN(DP_mult_217_n1568) );
  INV_X1 DP_mult_217_U1143 ( .A(DP_mult_217_n1534), .ZN(DP_mult_217_n1574) );
  OR2_X1 DP_mult_217_U1142 ( .A1(DP_mult_217_n1849), .A2(DP_mult_217_n1850), 
        .ZN(DP_mult_217_n1533) );
  BUF_X1 DP_mult_217_U1141 ( .A(DP_mult_217_n1747), .Z(DP_mult_217_n1577) );
  BUF_X1 DP_mult_217_U1140 ( .A(DP_mult_217_n1747), .Z(DP_mult_217_n1576) );
  INV_X1 DP_mult_217_U1139 ( .A(DP_mult_217_n1535), .ZN(DP_mult_217_n1573) );
  INV_X1 DP_mult_217_U1138 ( .A(DP_mult_217_n1536), .ZN(DP_mult_217_n1575) );
  INV_X1 DP_mult_217_U1137 ( .A(DP_mult_217_n1533), .ZN(DP_mult_217_n1580) );
  HA_X1 DP_mult_217_U1134 ( .A(DP_pipe01[0]), .B(DP_pipe01[1]), .CO(
        DP_mult_217_n727), .S(DP_mult_217_n1397) );
  FA_X1 DP_mult_217_U1133 ( .A(DP_pipe01[1]), .B(DP_pipe01[2]), .CI(
        DP_mult_217_n727), .CO(DP_mult_217_n726), .S(DP_mult_217_n1396) );
  FA_X1 DP_mult_217_U1132 ( .A(DP_pipe01[2]), .B(DP_pipe01[3]), .CI(
        DP_mult_217_n726), .CO(DP_mult_217_n725), .S(DP_mult_217_n1395) );
  FA_X1 DP_mult_217_U1131 ( .A(DP_pipe01[3]), .B(DP_pipe01[4]), .CI(
        DP_mult_217_n725), .CO(DP_mult_217_n724), .S(DP_mult_217_n1394) );
  FA_X1 DP_mult_217_U1130 ( .A(DP_pipe01[4]), .B(DP_pipe01[5]), .CI(
        DP_mult_217_n724), .CO(DP_mult_217_n723), .S(DP_mult_217_n1393) );
  FA_X1 DP_mult_217_U1129 ( .A(DP_pipe01[5]), .B(DP_pipe01[6]), .CI(
        DP_mult_217_n723), .CO(DP_mult_217_n722), .S(DP_mult_217_n1392) );
  FA_X1 DP_mult_217_U1128 ( .A(DP_pipe01[6]), .B(DP_pipe01[7]), .CI(
        DP_mult_217_n722), .CO(DP_mult_217_n721), .S(DP_mult_217_n1391) );
  FA_X1 DP_mult_217_U1127 ( .A(DP_pipe01[7]), .B(DP_pipe01[8]), .CI(
        DP_mult_217_n721), .CO(DP_mult_217_n720), .S(DP_mult_217_n1390) );
  FA_X1 DP_mult_217_U1126 ( .A(DP_pipe01[8]), .B(DP_pipe01[9]), .CI(
        DP_mult_217_n720), .CO(DP_mult_217_n719), .S(DP_mult_217_n1389) );
  FA_X1 DP_mult_217_U1125 ( .A(DP_pipe01[9]), .B(DP_pipe01[10]), .CI(
        DP_mult_217_n719), .CO(DP_mult_217_n718), .S(DP_mult_217_n1388) );
  FA_X1 DP_mult_217_U1124 ( .A(DP_pipe01[10]), .B(DP_pipe01[11]), .CI(
        DP_mult_217_n718), .CO(DP_mult_217_n717), .S(DP_mult_217_n1387) );
  FA_X1 DP_mult_217_U1123 ( .A(DP_pipe01[11]), .B(DP_pipe01[12]), .CI(
        DP_mult_217_n717), .CO(DP_mult_217_n716), .S(DP_mult_217_n1386) );
  FA_X1 DP_mult_217_U1122 ( .A(DP_pipe01[12]), .B(DP_pipe01[13]), .CI(
        DP_mult_217_n716), .CO(DP_mult_217_n715), .S(DP_mult_217_n1385) );
  FA_X1 DP_mult_217_U1121 ( .A(DP_pipe01[13]), .B(DP_pipe01[14]), .CI(
        DP_mult_217_n715), .CO(DP_mult_217_n714), .S(DP_mult_217_n1384) );
  FA_X1 DP_mult_217_U1120 ( .A(DP_pipe01[14]), .B(DP_pipe01[15]), .CI(
        DP_mult_217_n714), .CO(DP_mult_217_n713), .S(DP_mult_217_n1383) );
  FA_X1 DP_mult_217_U1119 ( .A(DP_pipe01[15]), .B(DP_pipe01[16]), .CI(
        DP_mult_217_n713), .CO(DP_mult_217_n712), .S(DP_mult_217_n1382) );
  FA_X1 DP_mult_217_U1118 ( .A(DP_pipe01[16]), .B(DP_pipe01[17]), .CI(
        DP_mult_217_n712), .CO(DP_mult_217_n711), .S(DP_mult_217_n1381) );
  FA_X1 DP_mult_217_U1117 ( .A(DP_pipe01[17]), .B(DP_pipe01[18]), .CI(
        DP_mult_217_n711), .CO(DP_mult_217_n710), .S(DP_mult_217_n1380) );
  FA_X1 DP_mult_217_U1116 ( .A(DP_pipe01[18]), .B(DP_pipe01[19]), .CI(
        DP_mult_217_n710), .CO(DP_mult_217_n709), .S(DP_mult_217_n1379) );
  FA_X1 DP_mult_217_U1115 ( .A(DP_pipe01[19]), .B(DP_pipe01[20]), .CI(
        DP_mult_217_n709), .CO(DP_mult_217_n708), .S(DP_mult_217_n1378) );
  FA_X1 DP_mult_217_U1114 ( .A(DP_pipe01[20]), .B(DP_pipe01[21]), .CI(
        DP_mult_217_n708), .CO(DP_mult_217_n707), .S(DP_mult_217_n1377) );
  FA_X1 DP_mult_217_U1113 ( .A(DP_pipe01[21]), .B(DP_pipe01[22]), .CI(
        DP_mult_217_n707), .CO(DP_mult_217_n706), .S(DP_mult_217_n1376) );
  FA_X1 DP_mult_217_U1112 ( .A(DP_pipe01[22]), .B(DP_mult_217_n1615), .CI(
        DP_mult_217_n706), .CO(DP_mult_217_n1374), .S(DP_mult_217_n1375) );
  HA_X1 DP_mult_217_U408 ( .A(DP_mult_217_n904), .B(DP_mult_217_n1598), .CO(
        DP_mult_217_n687), .S(DP_mult_217_n688) );
  HA_X1 DP_mult_217_U407 ( .A(DP_mult_217_n687), .B(DP_mult_217_n903), .CO(
        DP_mult_217_n685), .S(DP_mult_217_n686) );
  HA_X1 DP_mult_217_U406 ( .A(DP_mult_217_n685), .B(DP_mult_217_n902), .CO(
        DP_mult_217_n683), .S(DP_mult_217_n684) );
  HA_X1 DP_mult_217_U405 ( .A(DP_mult_217_n878), .B(DP_mult_217_n1600), .CO(
        DP_mult_217_n681), .S(DP_mult_217_n682) );
  FA_X1 DP_mult_217_U404 ( .A(DP_mult_217_n901), .B(DP_mult_217_n682), .CI(
        DP_mult_217_n683), .CO(DP_mult_217_n679), .S(DP_mult_217_n680) );
  HA_X1 DP_mult_217_U403 ( .A(DP_mult_217_n681), .B(DP_mult_217_n877), .CO(
        DP_mult_217_n677), .S(DP_mult_217_n678) );
  FA_X1 DP_mult_217_U402 ( .A(DP_mult_217_n900), .B(DP_mult_217_n678), .CI(
        DP_mult_217_n679), .CO(DP_mult_217_n675), .S(DP_mult_217_n676) );
  HA_X1 DP_mult_217_U401 ( .A(DP_mult_217_n677), .B(DP_mult_217_n876), .CO(
        DP_mult_217_n673), .S(DP_mult_217_n674) );
  FA_X1 DP_mult_217_U400 ( .A(DP_mult_217_n899), .B(DP_mult_217_n674), .CI(
        DP_mult_217_n675), .CO(DP_mult_217_n671), .S(DP_mult_217_n672) );
  HA_X1 DP_mult_217_U399 ( .A(DP_mult_217_n852), .B(DP_mult_217_n1602), .CO(
        DP_mult_217_n669), .S(DP_mult_217_n670) );
  FA_X1 DP_mult_217_U398 ( .A(DP_mult_217_n875), .B(DP_mult_217_n670), .CI(
        DP_mult_217_n673), .CO(DP_mult_217_n667), .S(DP_mult_217_n668) );
  FA_X1 DP_mult_217_U397 ( .A(DP_mult_217_n898), .B(DP_mult_217_n668), .CI(
        DP_mult_217_n671), .CO(DP_mult_217_n665), .S(DP_mult_217_n666) );
  HA_X1 DP_mult_217_U396 ( .A(DP_mult_217_n669), .B(DP_mult_217_n851), .CO(
        DP_mult_217_n663), .S(DP_mult_217_n664) );
  FA_X1 DP_mult_217_U395 ( .A(DP_mult_217_n874), .B(DP_mult_217_n664), .CI(
        DP_mult_217_n667), .CO(DP_mult_217_n661), .S(DP_mult_217_n662) );
  FA_X1 DP_mult_217_U394 ( .A(DP_mult_217_n897), .B(DP_mult_217_n662), .CI(
        DP_mult_217_n665), .CO(DP_mult_217_n659), .S(DP_mult_217_n660) );
  HA_X1 DP_mult_217_U393 ( .A(DP_mult_217_n663), .B(DP_mult_217_n850), .CO(
        DP_mult_217_n657), .S(DP_mult_217_n658) );
  FA_X1 DP_mult_217_U392 ( .A(DP_mult_217_n873), .B(DP_mult_217_n658), .CI(
        DP_mult_217_n661), .CO(DP_mult_217_n655), .S(DP_mult_217_n656) );
  FA_X1 DP_mult_217_U391 ( .A(DP_mult_217_n896), .B(DP_mult_217_n656), .CI(
        DP_mult_217_n659), .CO(DP_mult_217_n653), .S(DP_mult_217_n654) );
  HA_X1 DP_mult_217_U390 ( .A(DP_mult_217_n826), .B(DP_mult_217_n1604), .CO(
        DP_mult_217_n651), .S(DP_mult_217_n652) );
  FA_X1 DP_mult_217_U389 ( .A(DP_mult_217_n849), .B(DP_mult_217_n652), .CI(
        DP_mult_217_n657), .CO(DP_mult_217_n649), .S(DP_mult_217_n650) );
  FA_X1 DP_mult_217_U388 ( .A(DP_mult_217_n872), .B(DP_mult_217_n650), .CI(
        DP_mult_217_n655), .CO(DP_mult_217_n647), .S(DP_mult_217_n648) );
  FA_X1 DP_mult_217_U387 ( .A(DP_mult_217_n895), .B(DP_mult_217_n648), .CI(
        DP_mult_217_n653), .CO(DP_mult_217_n645), .S(DP_mult_217_n646) );
  HA_X1 DP_mult_217_U386 ( .A(DP_mult_217_n651), .B(DP_mult_217_n825), .CO(
        DP_mult_217_n643), .S(DP_mult_217_n644) );
  FA_X1 DP_mult_217_U385 ( .A(DP_mult_217_n848), .B(DP_mult_217_n644), .CI(
        DP_mult_217_n649), .CO(DP_mult_217_n641), .S(DP_mult_217_n642) );
  FA_X1 DP_mult_217_U384 ( .A(DP_mult_217_n871), .B(DP_mult_217_n642), .CI(
        DP_mult_217_n647), .CO(DP_mult_217_n639), .S(DP_mult_217_n640) );
  FA_X1 DP_mult_217_U383 ( .A(DP_mult_217_n894), .B(DP_mult_217_n640), .CI(
        DP_mult_217_n645), .CO(DP_mult_217_n637), .S(DP_mult_217_n638) );
  HA_X1 DP_mult_217_U382 ( .A(DP_mult_217_n643), .B(DP_mult_217_n824), .CO(
        DP_mult_217_n635), .S(DP_mult_217_n636) );
  FA_X1 DP_mult_217_U381 ( .A(DP_mult_217_n847), .B(DP_mult_217_n636), .CI(
        DP_mult_217_n641), .CO(DP_mult_217_n633), .S(DP_mult_217_n634) );
  FA_X1 DP_mult_217_U380 ( .A(DP_mult_217_n870), .B(DP_mult_217_n634), .CI(
        DP_mult_217_n639), .CO(DP_mult_217_n631), .S(DP_mult_217_n632) );
  FA_X1 DP_mult_217_U379 ( .A(DP_mult_217_n893), .B(DP_mult_217_n632), .CI(
        DP_mult_217_n637), .CO(DP_mult_217_n629), .S(DP_mult_217_n630) );
  HA_X1 DP_mult_217_U378 ( .A(DP_mult_217_n800), .B(DP_mult_217_n1606), .CO(
        DP_mult_217_n627), .S(DP_mult_217_n628) );
  FA_X1 DP_mult_217_U377 ( .A(DP_mult_217_n823), .B(DP_mult_217_n628), .CI(
        DP_mult_217_n635), .CO(DP_mult_217_n625), .S(DP_mult_217_n626) );
  FA_X1 DP_mult_217_U376 ( .A(DP_mult_217_n846), .B(DP_mult_217_n626), .CI(
        DP_mult_217_n633), .CO(DP_mult_217_n623), .S(DP_mult_217_n624) );
  FA_X1 DP_mult_217_U375 ( .A(DP_mult_217_n869), .B(DP_mult_217_n624), .CI(
        DP_mult_217_n631), .CO(DP_mult_217_n621), .S(DP_mult_217_n622) );
  FA_X1 DP_mult_217_U374 ( .A(DP_mult_217_n892), .B(DP_mult_217_n622), .CI(
        DP_mult_217_n629), .CO(DP_mult_217_n619), .S(DP_mult_217_n620) );
  HA_X1 DP_mult_217_U373 ( .A(DP_mult_217_n627), .B(DP_mult_217_n799), .CO(
        DP_mult_217_n617), .S(DP_mult_217_n618) );
  FA_X1 DP_mult_217_U372 ( .A(DP_mult_217_n822), .B(DP_mult_217_n618), .CI(
        DP_mult_217_n625), .CO(DP_mult_217_n615), .S(DP_mult_217_n616) );
  FA_X1 DP_mult_217_U371 ( .A(DP_mult_217_n845), .B(DP_mult_217_n616), .CI(
        DP_mult_217_n623), .CO(DP_mult_217_n613), .S(DP_mult_217_n614) );
  FA_X1 DP_mult_217_U370 ( .A(DP_mult_217_n868), .B(DP_mult_217_n614), .CI(
        DP_mult_217_n621), .CO(DP_mult_217_n611), .S(DP_mult_217_n612) );
  FA_X1 DP_mult_217_U369 ( .A(DP_mult_217_n891), .B(DP_mult_217_n612), .CI(
        DP_mult_217_n619), .CO(DP_mult_217_n609), .S(DP_mult_217_n610) );
  HA_X1 DP_mult_217_U368 ( .A(DP_mult_217_n617), .B(DP_mult_217_n798), .CO(
        DP_mult_217_n607), .S(DP_mult_217_n608) );
  FA_X1 DP_mult_217_U367 ( .A(DP_mult_217_n821), .B(DP_mult_217_n608), .CI(
        DP_mult_217_n615), .CO(DP_mult_217_n605), .S(DP_mult_217_n606) );
  FA_X1 DP_mult_217_U366 ( .A(DP_mult_217_n844), .B(DP_mult_217_n606), .CI(
        DP_mult_217_n613), .CO(DP_mult_217_n603), .S(DP_mult_217_n604) );
  FA_X1 DP_mult_217_U365 ( .A(DP_mult_217_n867), .B(DP_mult_217_n604), .CI(
        DP_mult_217_n611), .CO(DP_mult_217_n601), .S(DP_mult_217_n602) );
  FA_X1 DP_mult_217_U364 ( .A(DP_mult_217_n890), .B(DP_mult_217_n602), .CI(
        DP_mult_217_n609), .CO(DP_mult_217_n599), .S(DP_mult_217_n600) );
  HA_X1 DP_mult_217_U363 ( .A(DP_mult_217_n774), .B(DP_mult_217_n1608), .CO(
        DP_mult_217_n597), .S(DP_mult_217_n598) );
  FA_X1 DP_mult_217_U362 ( .A(DP_mult_217_n797), .B(DP_mult_217_n598), .CI(
        DP_mult_217_n607), .CO(DP_mult_217_n595), .S(DP_mult_217_n596) );
  FA_X1 DP_mult_217_U361 ( .A(DP_mult_217_n820), .B(DP_mult_217_n596), .CI(
        DP_mult_217_n605), .CO(DP_mult_217_n593), .S(DP_mult_217_n594) );
  FA_X1 DP_mult_217_U360 ( .A(DP_mult_217_n843), .B(DP_mult_217_n594), .CI(
        DP_mult_217_n603), .CO(DP_mult_217_n591), .S(DP_mult_217_n592) );
  FA_X1 DP_mult_217_U359 ( .A(DP_mult_217_n866), .B(DP_mult_217_n592), .CI(
        DP_mult_217_n601), .CO(DP_mult_217_n589), .S(DP_mult_217_n590) );
  FA_X1 DP_mult_217_U358 ( .A(DP_mult_217_n889), .B(DP_mult_217_n590), .CI(
        DP_mult_217_n599), .CO(DP_mult_217_n587), .S(DP_mult_217_n588) );
  HA_X1 DP_mult_217_U357 ( .A(DP_mult_217_n597), .B(DP_mult_217_n773), .CO(
        DP_mult_217_n585), .S(DP_mult_217_n586) );
  FA_X1 DP_mult_217_U356 ( .A(DP_mult_217_n796), .B(DP_mult_217_n586), .CI(
        DP_mult_217_n595), .CO(DP_mult_217_n583), .S(DP_mult_217_n584) );
  FA_X1 DP_mult_217_U355 ( .A(DP_mult_217_n819), .B(DP_mult_217_n584), .CI(
        DP_mult_217_n593), .CO(DP_mult_217_n581), .S(DP_mult_217_n582) );
  FA_X1 DP_mult_217_U354 ( .A(DP_mult_217_n842), .B(DP_mult_217_n582), .CI(
        DP_mult_217_n591), .CO(DP_mult_217_n579), .S(DP_mult_217_n580) );
  FA_X1 DP_mult_217_U353 ( .A(DP_mult_217_n865), .B(DP_mult_217_n580), .CI(
        DP_mult_217_n589), .CO(DP_mult_217_n577), .S(DP_mult_217_n578) );
  FA_X1 DP_mult_217_U352 ( .A(DP_mult_217_n888), .B(DP_mult_217_n578), .CI(
        DP_mult_217_n587), .CO(DP_mult_217_n575), .S(DP_mult_217_n576) );
  HA_X1 DP_mult_217_U351 ( .A(DP_mult_217_n585), .B(DP_mult_217_n772), .CO(
        DP_mult_217_n573), .S(DP_mult_217_n574) );
  FA_X1 DP_mult_217_U350 ( .A(DP_mult_217_n795), .B(DP_mult_217_n574), .CI(
        DP_mult_217_n583), .CO(DP_mult_217_n571), .S(DP_mult_217_n572) );
  FA_X1 DP_mult_217_U349 ( .A(DP_mult_217_n818), .B(DP_mult_217_n572), .CI(
        DP_mult_217_n581), .CO(DP_mult_217_n569), .S(DP_mult_217_n570) );
  FA_X1 DP_mult_217_U348 ( .A(DP_mult_217_n841), .B(DP_mult_217_n570), .CI(
        DP_mult_217_n579), .CO(DP_mult_217_n567), .S(DP_mult_217_n568) );
  FA_X1 DP_mult_217_U347 ( .A(DP_mult_217_n864), .B(DP_mult_217_n568), .CI(
        DP_mult_217_n577), .CO(DP_mult_217_n565), .S(DP_mult_217_n566) );
  FA_X1 DP_mult_217_U346 ( .A(DP_mult_217_n887), .B(DP_mult_217_n566), .CI(
        DP_mult_217_n575), .CO(DP_mult_217_n563), .S(DP_mult_217_n564) );
  HA_X1 DP_mult_217_U345 ( .A(DP_mult_217_n748), .B(DP_mult_217_n1610), .CO(
        DP_mult_217_n561), .S(DP_mult_217_n562) );
  FA_X1 DP_mult_217_U344 ( .A(DP_mult_217_n771), .B(DP_mult_217_n562), .CI(
        DP_mult_217_n573), .CO(DP_mult_217_n559), .S(DP_mult_217_n560) );
  FA_X1 DP_mult_217_U343 ( .A(DP_mult_217_n794), .B(DP_mult_217_n560), .CI(
        DP_mult_217_n571), .CO(DP_mult_217_n557), .S(DP_mult_217_n558) );
  FA_X1 DP_mult_217_U342 ( .A(DP_mult_217_n817), .B(DP_mult_217_n558), .CI(
        DP_mult_217_n569), .CO(DP_mult_217_n555), .S(DP_mult_217_n556) );
  FA_X1 DP_mult_217_U341 ( .A(DP_mult_217_n840), .B(DP_mult_217_n556), .CI(
        DP_mult_217_n567), .CO(DP_mult_217_n553), .S(DP_mult_217_n554) );
  FA_X1 DP_mult_217_U340 ( .A(DP_mult_217_n863), .B(DP_mult_217_n554), .CI(
        DP_mult_217_n565), .CO(DP_mult_217_n551), .S(DP_mult_217_n552) );
  FA_X1 DP_mult_217_U339 ( .A(DP_mult_217_n886), .B(DP_mult_217_n552), .CI(
        DP_mult_217_n563), .CO(DP_mult_217_n549), .S(DP_mult_217_n550) );
  HA_X1 DP_mult_217_U338 ( .A(DP_mult_217_n561), .B(DP_mult_217_n747), .CO(
        DP_mult_217_n547), .S(DP_mult_217_n548) );
  FA_X1 DP_mult_217_U337 ( .A(DP_mult_217_n770), .B(DP_mult_217_n548), .CI(
        DP_mult_217_n559), .CO(DP_mult_217_n545), .S(DP_mult_217_n546) );
  FA_X1 DP_mult_217_U336 ( .A(DP_mult_217_n793), .B(DP_mult_217_n546), .CI(
        DP_mult_217_n557), .CO(DP_mult_217_n543), .S(DP_mult_217_n544) );
  FA_X1 DP_mult_217_U335 ( .A(DP_mult_217_n816), .B(DP_mult_217_n544), .CI(
        DP_mult_217_n555), .CO(DP_mult_217_n541), .S(DP_mult_217_n542) );
  FA_X1 DP_mult_217_U334 ( .A(DP_mult_217_n839), .B(DP_mult_217_n542), .CI(
        DP_mult_217_n553), .CO(DP_mult_217_n539), .S(DP_mult_217_n540) );
  FA_X1 DP_mult_217_U333 ( .A(DP_mult_217_n862), .B(DP_mult_217_n540), .CI(
        DP_mult_217_n551), .CO(DP_mult_217_n537), .S(DP_mult_217_n538) );
  FA_X1 DP_mult_217_U332 ( .A(DP_mult_217_n885), .B(DP_mult_217_n538), .CI(
        DP_mult_217_n549), .CO(DP_mult_217_n535), .S(DP_mult_217_n536) );
  HA_X1 DP_mult_217_U331 ( .A(DP_mult_217_n547), .B(DP_mult_217_n746), .CO(
        DP_mult_217_n533), .S(DP_mult_217_n534) );
  FA_X1 DP_mult_217_U330 ( .A(DP_mult_217_n769), .B(DP_mult_217_n534), .CI(
        DP_mult_217_n545), .CO(DP_mult_217_n531), .S(DP_mult_217_n532) );
  FA_X1 DP_mult_217_U329 ( .A(DP_mult_217_n792), .B(DP_mult_217_n532), .CI(
        DP_mult_217_n543), .CO(DP_mult_217_n529), .S(DP_mult_217_n530) );
  FA_X1 DP_mult_217_U328 ( .A(DP_mult_217_n815), .B(DP_mult_217_n530), .CI(
        DP_mult_217_n541), .CO(DP_mult_217_n527), .S(DP_mult_217_n528) );
  FA_X1 DP_mult_217_U327 ( .A(DP_mult_217_n838), .B(DP_mult_217_n528), .CI(
        DP_mult_217_n539), .CO(DP_mult_217_n525), .S(DP_mult_217_n526) );
  FA_X1 DP_mult_217_U326 ( .A(DP_mult_217_n861), .B(DP_mult_217_n526), .CI(
        DP_mult_217_n537), .CO(DP_mult_217_n523), .S(DP_mult_217_n524) );
  FA_X1 DP_mult_217_U325 ( .A(DP_mult_217_n884), .B(DP_mult_217_n524), .CI(
        DP_mult_217_n535), .CO(DP_mult_217_n521), .S(DP_mult_217_n522) );
  HA_X1 DP_mult_217_U324 ( .A(DP_mult_217_n533), .B(DP_mult_217_n745), .CO(
        DP_mult_217_n519), .S(DP_mult_217_n520) );
  FA_X1 DP_mult_217_U323 ( .A(DP_mult_217_n768), .B(DP_mult_217_n520), .CI(
        DP_mult_217_n531), .CO(DP_mult_217_n517), .S(DP_mult_217_n518) );
  FA_X1 DP_mult_217_U322 ( .A(DP_mult_217_n791), .B(DP_mult_217_n518), .CI(
        DP_mult_217_n529), .CO(DP_mult_217_n515), .S(DP_mult_217_n516) );
  FA_X1 DP_mult_217_U321 ( .A(DP_mult_217_n814), .B(DP_mult_217_n516), .CI(
        DP_mult_217_n527), .CO(DP_mult_217_n513), .S(DP_mult_217_n514) );
  FA_X1 DP_mult_217_U320 ( .A(DP_mult_217_n837), .B(DP_mult_217_n514), .CI(
        DP_mult_217_n525), .CO(DP_mult_217_n511), .S(DP_mult_217_n512) );
  FA_X1 DP_mult_217_U319 ( .A(DP_mult_217_n860), .B(DP_mult_217_n512), .CI(
        DP_mult_217_n523), .CO(DP_mult_217_n509), .S(DP_mult_217_n510) );
  FA_X1 DP_mult_217_U318 ( .A(DP_mult_217_n883), .B(DP_mult_217_n510), .CI(
        DP_mult_217_n521), .CO(DP_mult_217_n507), .S(DP_mult_217_n508) );
  FA_X1 DP_mult_217_U315 ( .A(DP_mult_217_n506), .B(DP_mult_217_n744), .CI(
        DP_mult_217_n767), .CO(DP_mult_217_n504), .S(DP_mult_217_n505) );
  FA_X1 DP_mult_217_U314 ( .A(DP_mult_217_n505), .B(DP_mult_217_n517), .CI(
        DP_mult_217_n790), .CO(DP_mult_217_n502), .S(DP_mult_217_n503) );
  FA_X1 DP_mult_217_U313 ( .A(DP_mult_217_n503), .B(DP_mult_217_n515), .CI(
        DP_mult_217_n813), .CO(DP_mult_217_n500), .S(DP_mult_217_n501) );
  FA_X1 DP_mult_217_U312 ( .A(DP_mult_217_n501), .B(DP_mult_217_n513), .CI(
        DP_mult_217_n836), .CO(DP_mult_217_n498), .S(DP_mult_217_n499) );
  FA_X1 DP_mult_217_U311 ( .A(DP_mult_217_n499), .B(DP_mult_217_n511), .CI(
        DP_mult_217_n859), .CO(DP_mult_217_n496), .S(DP_mult_217_n497) );
  FA_X1 DP_mult_217_U310 ( .A(DP_mult_217_n497), .B(DP_mult_217_n509), .CI(
        DP_mult_217_n882), .CO(DP_mult_217_n494), .S(DP_mult_217_n495) );
  FA_X1 DP_mult_217_U308 ( .A(DP_mult_217_n743), .B(DP_mult_217_n493), .CI(
        DP_mult_217_n766), .CO(DP_mult_217_n491), .S(DP_mult_217_n492) );
  FA_X1 DP_mult_217_U307 ( .A(DP_mult_217_n492), .B(DP_mult_217_n504), .CI(
        DP_mult_217_n789), .CO(DP_mult_217_n489), .S(DP_mult_217_n490) );
  FA_X1 DP_mult_217_U306 ( .A(DP_mult_217_n490), .B(DP_mult_217_n502), .CI(
        DP_mult_217_n500), .CO(DP_mult_217_n487), .S(DP_mult_217_n488) );
  FA_X1 DP_mult_217_U305 ( .A(DP_mult_217_n488), .B(DP_mult_217_n812), .CI(
        DP_mult_217_n835), .CO(DP_mult_217_n485), .S(DP_mult_217_n486) );
  FA_X1 DP_mult_217_U304 ( .A(DP_mult_217_n486), .B(DP_mult_217_n498), .CI(
        DP_mult_217_n496), .CO(DP_mult_217_n483), .S(DP_mult_217_n484) );
  FA_X1 DP_mult_217_U303 ( .A(DP_mult_217_n484), .B(DP_mult_217_n858), .CI(
        DP_mult_217_n881), .CO(DP_mult_217_n481), .S(DP_mult_217_n482) );
  FA_X1 DP_mult_217_U301 ( .A(DP_mult_217_n742), .B(DP_mult_217_n493), .CI(
        DP_mult_217_n491), .CO(DP_mult_217_n477), .S(DP_mult_217_n478) );
  FA_X1 DP_mult_217_U300 ( .A(DP_mult_217_n478), .B(DP_mult_217_n765), .CI(
        DP_mult_217_n788), .CO(DP_mult_217_n475), .S(DP_mult_217_n476) );
  FA_X1 DP_mult_217_U299 ( .A(DP_mult_217_n476), .B(DP_mult_217_n489), .CI(
        DP_mult_217_n487), .CO(DP_mult_217_n473), .S(DP_mult_217_n474) );
  FA_X1 DP_mult_217_U298 ( .A(DP_mult_217_n474), .B(DP_mult_217_n811), .CI(
        DP_mult_217_n834), .CO(DP_mult_217_n471), .S(DP_mult_217_n472) );
  FA_X1 DP_mult_217_U297 ( .A(DP_mult_217_n472), .B(DP_mult_217_n485), .CI(
        DP_mult_217_n483), .CO(DP_mult_217_n469), .S(DP_mult_217_n470) );
  FA_X1 DP_mult_217_U296 ( .A(DP_mult_217_n880), .B(DP_mult_217_n857), .CI(
        DP_mult_217_n470), .CO(DP_mult_217_n467), .S(DP_mult_217_n468) );
  FA_X1 DP_mult_217_U295 ( .A(DP_mult_217_n479), .B(DP_mult_217_n879), .CI(
        DP_mult_217_n741), .CO(DP_mult_217_n465), .S(DP_mult_217_n466) );
  FA_X1 DP_mult_217_U294 ( .A(DP_mult_217_n764), .B(DP_mult_217_n466), .CI(
        DP_mult_217_n477), .CO(DP_mult_217_n463), .S(DP_mult_217_n464) );
  FA_X1 DP_mult_217_U293 ( .A(DP_mult_217_n475), .B(DP_mult_217_n464), .CI(
        DP_mult_217_n787), .CO(DP_mult_217_n461), .S(DP_mult_217_n462) );
  FA_X1 DP_mult_217_U292 ( .A(DP_mult_217_n810), .B(DP_mult_217_n462), .CI(
        DP_mult_217_n473), .CO(DP_mult_217_n459), .S(DP_mult_217_n460) );
  FA_X1 DP_mult_217_U291 ( .A(DP_mult_217_n471), .B(DP_mult_217_n460), .CI(
        DP_mult_217_n833), .CO(DP_mult_217_n457), .S(DP_mult_217_n458) );
  FA_X1 DP_mult_217_U290 ( .A(DP_mult_217_n856), .B(DP_mult_217_n458), .CI(
        DP_mult_217_n469), .CO(DP_mult_217_n455), .S(DP_mult_217_n456) );
  FA_X1 DP_mult_217_U288 ( .A(DP_mult_217_n454), .B(DP_mult_217_n465), .CI(
        DP_mult_217_n763), .CO(DP_mult_217_n452), .S(DP_mult_217_n453) );
  FA_X1 DP_mult_217_U287 ( .A(DP_mult_217_n453), .B(DP_mult_217_n463), .CI(
        DP_mult_217_n786), .CO(DP_mult_217_n450), .S(DP_mult_217_n451) );
  FA_X1 DP_mult_217_U286 ( .A(DP_mult_217_n451), .B(DP_mult_217_n461), .CI(
        DP_mult_217_n809), .CO(DP_mult_217_n448), .S(DP_mult_217_n449) );
  FA_X1 DP_mult_217_U285 ( .A(DP_mult_217_n449), .B(DP_mult_217_n459), .CI(
        DP_mult_217_n832), .CO(DP_mult_217_n446), .S(DP_mult_217_n447) );
  FA_X1 DP_mult_217_U284 ( .A(DP_mult_217_n447), .B(DP_mult_217_n457), .CI(
        DP_mult_217_n855), .CO(DP_mult_217_n444), .S(DP_mult_217_n445) );
  FA_X1 DP_mult_217_U282 ( .A(DP_mult_217_n740), .B(DP_mult_217_n454), .CI(
        DP_mult_217_n762), .CO(DP_mult_217_n440), .S(DP_mult_217_n441) );
  FA_X1 DP_mult_217_U281 ( .A(DP_mult_217_n441), .B(DP_mult_217_n452), .CI(
        DP_mult_217_n450), .CO(DP_mult_217_n438), .S(DP_mult_217_n439) );
  FA_X1 DP_mult_217_U280 ( .A(DP_mult_217_n439), .B(DP_mult_217_n785), .CI(
        DP_mult_217_n808), .CO(DP_mult_217_n436), .S(DP_mult_217_n437) );
  FA_X1 DP_mult_217_U279 ( .A(DP_mult_217_n437), .B(DP_mult_217_n448), .CI(
        DP_mult_217_n446), .CO(DP_mult_217_n434), .S(DP_mult_217_n435) );
  FA_X1 DP_mult_217_U278 ( .A(DP_mult_217_n854), .B(DP_mult_217_n831), .CI(
        DP_mult_217_n435), .CO(DP_mult_217_n432), .S(DP_mult_217_n433) );
  FA_X1 DP_mult_217_U277 ( .A(DP_mult_217_n442), .B(DP_mult_217_n853), .CI(
        DP_mult_217_n739), .CO(DP_mult_217_n430), .S(DP_mult_217_n431) );
  FA_X1 DP_mult_217_U276 ( .A(DP_mult_217_n440), .B(DP_mult_217_n431), .CI(
        DP_mult_217_n761), .CO(DP_mult_217_n428), .S(DP_mult_217_n429) );
  FA_X1 DP_mult_217_U275 ( .A(DP_mult_217_n784), .B(DP_mult_217_n429), .CI(
        DP_mult_217_n438), .CO(DP_mult_217_n426), .S(DP_mult_217_n427) );
  FA_X1 DP_mult_217_U274 ( .A(DP_mult_217_n436), .B(DP_mult_217_n427), .CI(
        DP_mult_217_n807), .CO(DP_mult_217_n424), .S(DP_mult_217_n425) );
  FA_X1 DP_mult_217_U273 ( .A(DP_mult_217_n830), .B(DP_mult_217_n425), .CI(
        DP_mult_217_n434), .CO(DP_mult_217_n422), .S(DP_mult_217_n423) );
  FA_X1 DP_mult_217_U271 ( .A(DP_mult_217_n421), .B(DP_mult_217_n430), .CI(
        DP_mult_217_n760), .CO(DP_mult_217_n419), .S(DP_mult_217_n420) );
  FA_X1 DP_mult_217_U270 ( .A(DP_mult_217_n420), .B(DP_mult_217_n428), .CI(
        DP_mult_217_n783), .CO(DP_mult_217_n417), .S(DP_mult_217_n418) );
  FA_X1 DP_mult_217_U269 ( .A(DP_mult_217_n418), .B(DP_mult_217_n426), .CI(
        DP_mult_217_n806), .CO(DP_mult_217_n415), .S(DP_mult_217_n416) );
  FA_X1 DP_mult_217_U268 ( .A(DP_mult_217_n416), .B(DP_mult_217_n424), .CI(
        DP_mult_217_n829), .CO(DP_mult_217_n413), .S(DP_mult_217_n414) );
  FA_X1 DP_mult_217_U266 ( .A(DP_mult_217_n738), .B(DP_mult_217_n421), .CI(
        DP_mult_217_n419), .CO(DP_mult_217_n409), .S(DP_mult_217_n410) );
  FA_X1 DP_mult_217_U265 ( .A(DP_mult_217_n410), .B(DP_mult_217_n759), .CI(
        DP_mult_217_n782), .CO(DP_mult_217_n407), .S(DP_mult_217_n408) );
  FA_X1 DP_mult_217_U264 ( .A(DP_mult_217_n408), .B(DP_mult_217_n417), .CI(
        DP_mult_217_n415), .CO(DP_mult_217_n405), .S(DP_mult_217_n406) );
  FA_X1 DP_mult_217_U263 ( .A(DP_mult_217_n828), .B(DP_mult_217_n805), .CI(
        DP_mult_217_n406), .CO(DP_mult_217_n403), .S(DP_mult_217_n404) );
  FA_X1 DP_mult_217_U262 ( .A(DP_mult_217_n411), .B(DP_mult_217_n827), .CI(
        DP_mult_217_n737), .CO(DP_mult_217_n387), .S(DP_mult_217_n402) );
  FA_X1 DP_mult_217_U261 ( .A(DP_mult_217_n758), .B(DP_mult_217_n402), .CI(
        DP_mult_217_n409), .CO(DP_mult_217_n400), .S(DP_mult_217_n401) );
  FA_X1 DP_mult_217_U260 ( .A(DP_mult_217_n407), .B(DP_mult_217_n401), .CI(
        DP_mult_217_n781), .CO(DP_mult_217_n398), .S(DP_mult_217_n399) );
  FA_X1 DP_mult_217_U259 ( .A(DP_mult_217_n804), .B(DP_mult_217_n399), .CI(
        DP_mult_217_n405), .CO(DP_mult_217_n396), .S(DP_mult_217_n397) );
  FA_X1 DP_mult_217_U257 ( .A(DP_mult_217_n395), .B(DP_mult_217_n736), .CI(
        DP_mult_217_n757), .CO(DP_mult_217_n393), .S(DP_mult_217_n394) );
  FA_X1 DP_mult_217_U256 ( .A(DP_mult_217_n394), .B(DP_mult_217_n400), .CI(
        DP_mult_217_n780), .CO(DP_mult_217_n391), .S(DP_mult_217_n392) );
  FA_X1 DP_mult_217_U255 ( .A(DP_mult_217_n392), .B(DP_mult_217_n398), .CI(
        DP_mult_217_n803), .CO(DP_mult_217_n389), .S(DP_mult_217_n390) );
  FA_X1 DP_mult_217_U253 ( .A(DP_mult_217_n735), .B(DP_mult_217_n395), .CI(
        DP_mult_217_n756), .CO(DP_mult_217_n385), .S(DP_mult_217_n386) );
  FA_X1 DP_mult_217_U252 ( .A(DP_mult_217_n386), .B(DP_mult_217_n393), .CI(
        DP_mult_217_n391), .CO(DP_mult_217_n383), .S(DP_mult_217_n384) );
  FA_X1 DP_mult_217_U251 ( .A(DP_mult_217_n802), .B(DP_mult_217_n779), .CI(
        DP_mult_217_n384), .CO(DP_mult_217_n381), .S(DP_mult_217_n382) );
  FA_X1 DP_mult_217_U250 ( .A(DP_mult_217_n387), .B(DP_mult_217_n801), .CI(
        DP_mult_217_n734), .CO(DP_mult_217_n379), .S(DP_mult_217_n380) );
  FA_X1 DP_mult_217_U249 ( .A(DP_mult_217_n385), .B(DP_mult_217_n380), .CI(
        DP_mult_217_n755), .CO(DP_mult_217_n377), .S(DP_mult_217_n378) );
  FA_X1 DP_mult_217_U248 ( .A(DP_mult_217_n778), .B(DP_mult_217_n378), .CI(
        DP_mult_217_n383), .CO(DP_mult_217_n375), .S(DP_mult_217_n376) );
  FA_X1 DP_mult_217_U246 ( .A(DP_mult_217_n374), .B(DP_mult_217_n379), .CI(
        DP_mult_217_n754), .CO(DP_mult_217_n372), .S(DP_mult_217_n373) );
  FA_X1 DP_mult_217_U245 ( .A(DP_mult_217_n373), .B(DP_mult_217_n377), .CI(
        DP_mult_217_n777), .CO(DP_mult_217_n370), .S(DP_mult_217_n371) );
  FA_X1 DP_mult_217_U243 ( .A(DP_mult_217_n733), .B(DP_mult_217_n374), .CI(
        DP_mult_217_n372), .CO(DP_mult_217_n366), .S(DP_mult_217_n367) );
  FA_X1 DP_mult_217_U242 ( .A(DP_mult_217_n776), .B(DP_mult_217_n753), .CI(
        DP_mult_217_n367), .CO(DP_mult_217_n364), .S(DP_mult_217_n365) );
  FA_X1 DP_mult_217_U241 ( .A(DP_mult_217_n368), .B(DP_mult_217_n775), .CI(
        DP_mult_217_n732), .CO(DP_mult_217_n356), .S(DP_mult_217_n363) );
  FA_X1 DP_mult_217_U240 ( .A(DP_mult_217_n752), .B(DP_mult_217_n363), .CI(
        DP_mult_217_n366), .CO(DP_mult_217_n361), .S(DP_mult_217_n362) );
  FA_X1 DP_mult_217_U238 ( .A(DP_mult_217_n360), .B(DP_mult_217_n731), .CI(
        DP_mult_217_n751), .CO(DP_mult_217_n358), .S(DP_mult_217_n359) );
  FA_X1 DP_mult_217_U236 ( .A(DP_mult_217_n730), .B(DP_mult_217_n360), .CI(
        DP_mult_217_n750), .CO(DP_mult_217_n354), .S(DP_mult_217_n355) );
  FA_X1 DP_mult_217_U235 ( .A(DP_mult_217_n356), .B(DP_mult_217_n749), .CI(
        DP_mult_217_n729), .CO(DP_mult_217_n352), .S(DP_mult_217_n353) );
  FA_X1 DP_mult_217_U204 ( .A(DP_mult_217_n908), .B(DP_mult_217_n536), .CI(
        DP_mult_217_n326), .CO(DP_mult_217_n325), .S(DP_pipe0_coeff_pipe01[0])
         );
  FA_X1 DP_mult_217_U203 ( .A(DP_mult_217_n907), .B(DP_mult_217_n522), .CI(
        DP_mult_217_n325), .CO(DP_mult_217_n324), .S(DP_pipe0_coeff_pipe01[1])
         );
  FA_X1 DP_mult_217_U202 ( .A(DP_mult_217_n508), .B(DP_mult_217_n906), .CI(
        DP_mult_217_n324), .CO(DP_mult_217_n323), .S(DP_pipe0_coeff_pipe01[2])
         );
  FA_X1 DP_mult_217_U201 ( .A(DP_mult_217_n495), .B(DP_mult_217_n507), .CI(
        DP_mult_217_n323), .CO(DP_mult_217_n322), .S(DP_pipe0_coeff_pipe01[3])
         );
  FA_X1 DP_mult_217_U200 ( .A(DP_mult_217_n482), .B(DP_mult_217_n494), .CI(
        DP_mult_217_n322), .CO(DP_mult_217_n321), .S(DP_pipe0_coeff_pipe01[4])
         );
  FA_X1 DP_mult_217_U199 ( .A(DP_mult_217_n468), .B(DP_mult_217_n481), .CI(
        DP_mult_217_n321), .CO(DP_mult_217_n320), .S(DP_pipe0_coeff_pipe01[5])
         );
  FA_X1 DP_mult_217_U198 ( .A(DP_mult_217_n456), .B(DP_mult_217_n467), .CI(
        DP_mult_217_n320), .CO(DP_mult_217_n319), .S(DP_pipe0_coeff_pipe01[6])
         );
  FA_X1 DP_mult_217_U197 ( .A(DP_mult_217_n445), .B(DP_mult_217_n455), .CI(
        DP_mult_217_n319), .CO(DP_mult_217_n318), .S(DP_pipe0_coeff_pipe01[7])
         );
  FA_X1 DP_mult_217_U196 ( .A(DP_mult_217_n433), .B(DP_mult_217_n444), .CI(
        DP_mult_217_n318), .CO(DP_mult_217_n317), .S(DP_pipe0_coeff_pipe01[8])
         );
  FA_X1 DP_mult_217_U195 ( .A(DP_mult_217_n423), .B(DP_mult_217_n432), .CI(
        DP_mult_217_n317), .CO(DP_mult_217_n316), .S(DP_pipe0_coeff_pipe01[9])
         );
  FA_X1 DP_mult_217_U194 ( .A(DP_mult_217_n414), .B(DP_mult_217_n422), .CI(
        DP_mult_217_n316), .CO(DP_mult_217_n315), .S(DP_pipe0_coeff_pipe01[10]) );
  FA_X1 DP_mult_217_U193 ( .A(DP_mult_217_n404), .B(DP_mult_217_n413), .CI(
        DP_mult_217_n315), .CO(DP_mult_217_n314), .S(DP_pipe0_coeff_pipe01[11]) );
  FA_X1 DP_mult_217_U192 ( .A(DP_mult_217_n397), .B(DP_mult_217_n403), .CI(
        DP_mult_217_n314), .CO(DP_mult_217_n313), .S(DP_pipe0_coeff_pipe01[12]) );
  FA_X1 DP_mult_217_U191 ( .A(DP_mult_217_n390), .B(DP_mult_217_n396), .CI(
        DP_mult_217_n313), .CO(DP_mult_217_n312), .S(DP_pipe0_coeff_pipe01[13]) );
  FA_X1 DP_mult_217_U190 ( .A(DP_mult_217_n382), .B(DP_mult_217_n389), .CI(
        DP_mult_217_n312), .CO(DP_mult_217_n311), .S(DP_pipe0_coeff_pipe01[14]) );
  FA_X1 DP_mult_217_U189 ( .A(DP_mult_217_n376), .B(DP_mult_217_n381), .CI(
        DP_mult_217_n311), .CO(DP_mult_217_n310), .S(DP_pipe0_coeff_pipe01[15]) );
  FA_X1 DP_mult_217_U188 ( .A(DP_mult_217_n371), .B(DP_mult_217_n375), .CI(
        DP_mult_217_n310), .CO(DP_mult_217_n309), .S(DP_pipe0_coeff_pipe01[16]) );
  FA_X1 DP_mult_217_U187 ( .A(DP_mult_217_n365), .B(DP_mult_217_n370), .CI(
        DP_mult_217_n309), .CO(DP_mult_217_n308), .S(DP_pipe0_coeff_pipe01[17]) );
  FA_X1 DP_mult_217_U186 ( .A(DP_mult_217_n362), .B(DP_mult_217_n364), .CI(
        DP_mult_217_n308), .CO(DP_mult_217_n307), .S(DP_pipe0_coeff_pipe01[18]) );
  FA_X1 DP_mult_217_U185 ( .A(DP_mult_217_n359), .B(DP_mult_217_n361), .CI(
        DP_mult_217_n307), .CO(DP_mult_217_n306), .S(DP_pipe0_coeff_pipe01[19]) );
  FA_X1 DP_mult_217_U184 ( .A(DP_mult_217_n355), .B(DP_mult_217_n358), .CI(
        DP_mult_217_n306), .CO(DP_mult_217_n305), .S(DP_pipe0_coeff_pipe01[20]) );
  FA_X1 DP_mult_217_U183 ( .A(DP_mult_217_n353), .B(DP_mult_217_n354), .CI(
        DP_mult_217_n305), .CO(DP_mult_217_n304), .S(DP_pipe0_coeff_pipe01[21]) );
  FA_X1 DP_mult_217_U182 ( .A(DP_mult_217_n351), .B(DP_mult_217_n352), .CI(
        DP_mult_217_n304), .CO(DP_mult_217_n303), .S(DP_pipe0_coeff_pipe01[22]) );
  INV_X1 DP_mult_215_U1959 ( .A(DP_coeff_ret1[1]), .ZN(DP_mult_215_n2159) );
  NOR2_X1 DP_mult_215_U1958 ( .A1(DP_mult_215_n2159), .A2(DP_coeff_ret1[0]), 
        .ZN(DP_mult_215_n1636) );
  INV_X1 DP_mult_215_U1957 ( .A(DP_coeff_ret1[2]), .ZN(DP_mult_215_n1742) );
  XNOR2_X1 DP_mult_215_U1956 ( .A(DP_coeff_ret1[1]), .B(DP_mult_215_n1742), 
        .ZN(DP_mult_215_n2157) );
  AOI221_X1 DP_mult_215_U1955 ( .B1(DP_sw1_1_), .B2(DP_mult_215_n1563), .C1(
        DP_mult_215_n1396), .C2(DP_mult_215_n1555), .A(DP_mult_215_n1742), 
        .ZN(DP_mult_215_n2160) );
  INV_X1 DP_mult_215_U1954 ( .A(DP_coeff_ret1[0]), .ZN(DP_mult_215_n2158) );
  INV_X1 DP_mult_215_U1953 ( .A(DP_sw1_2_), .ZN(DP_mult_215_n1661) );
  INV_X1 DP_mult_215_U1952 ( .A(DP_mult_215_n1397), .ZN(DP_mult_215_n1650) );
  OAI22_X1 DP_mult_215_U1951 ( .A1(DP_mult_215_n1554), .A2(DP_mult_215_n1661), 
        .B1(DP_mult_215_n1564), .B2(DP_mult_215_n1650), .ZN(DP_mult_215_n2162)
         );
  AOI211_X1 DP_mult_215_U1950 ( .C1(DP_sw1_1_), .C2(DP_mult_215_n1561), .A(
        DP_mult_215_n2162), .B(DP_sw1_0_), .ZN(DP_mult_215_n2161) );
  AND2_X1 DP_mult_215_U1949 ( .A1(DP_mult_215_n2160), .A2(DP_mult_215_n2161), 
        .ZN(DP_mult_215_n2153) );
  INV_X1 DP_mult_215_U1948 ( .A(DP_mult_215_n1395), .ZN(DP_mult_215_n1657) );
  INV_X1 DP_mult_215_U1947 ( .A(DP_sw1_1_), .ZN(DP_mult_215_n1649) );
  OAI22_X1 DP_mult_215_U1946 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1657), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1649), .ZN(DP_mult_215_n2156)
         );
  AOI221_X1 DP_mult_215_U1945 ( .B1(DP_sw1_3_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_2_), .C2(DP_mult_215_n1563), .A(DP_mult_215_n2156), .ZN(
        DP_mult_215_n2155) );
  XNOR2_X1 DP_mult_215_U1944 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2155), 
        .ZN(DP_mult_215_n2154) );
  AOI222_X1 DP_mult_215_U1943 ( .A1(DP_mult_215_n2153), .A2(DP_mult_215_n2154), 
        .B1(DP_mult_215_n2153), .B2(DP_mult_215_n688), .C1(DP_mult_215_n688), 
        .C2(DP_mult_215_n2154), .ZN(DP_mult_215_n2148) );
  INV_X1 DP_mult_215_U1942 ( .A(DP_mult_215_n1394), .ZN(DP_mult_215_n1660) );
  OAI22_X1 DP_mult_215_U1941 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1660), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1661), .ZN(DP_mult_215_n2152)
         );
  AOI221_X1 DP_mult_215_U1940 ( .B1(DP_sw1_4_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_3_), .C2(DP_mult_215_n1563), .A(DP_mult_215_n2152), .ZN(
        DP_mult_215_n2151) );
  XNOR2_X1 DP_mult_215_U1939 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2151), 
        .ZN(DP_mult_215_n2149) );
  INV_X1 DP_mult_215_U1938 ( .A(DP_mult_215_n686), .ZN(DP_mult_215_n2150) );
  OAI222_X1 DP_mult_215_U1937 ( .A1(DP_mult_215_n2148), .A2(DP_mult_215_n2149), 
        .B1(DP_mult_215_n2148), .B2(DP_mult_215_n2150), .C1(DP_mult_215_n2150), 
        .C2(DP_mult_215_n2149), .ZN(DP_mult_215_n2144) );
  INV_X1 DP_mult_215_U1936 ( .A(DP_mult_215_n1393), .ZN(DP_mult_215_n1664) );
  INV_X1 DP_mult_215_U1935 ( .A(DP_sw1_3_), .ZN(DP_mult_215_n1665) );
  OAI22_X1 DP_mult_215_U1934 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1664), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1665), .ZN(DP_mult_215_n2147)
         );
  AOI221_X1 DP_mult_215_U1933 ( .B1(DP_sw1_5_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_4_), .C2(DP_mult_215_n1563), .A(DP_mult_215_n2147), .ZN(
        DP_mult_215_n2146) );
  XNOR2_X1 DP_mult_215_U1932 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2146), 
        .ZN(DP_mult_215_n2145) );
  AOI222_X1 DP_mult_215_U1931 ( .A1(DP_mult_215_n2144), .A2(DP_mult_215_n2145), 
        .B1(DP_mult_215_n2144), .B2(DP_mult_215_n684), .C1(DP_mult_215_n684), 
        .C2(DP_mult_215_n2145), .ZN(DP_mult_215_n2139) );
  INV_X1 DP_mult_215_U1930 ( .A(DP_mult_215_n1392), .ZN(DP_mult_215_n1668) );
  INV_X1 DP_mult_215_U1929 ( .A(DP_sw1_4_), .ZN(DP_mult_215_n1669) );
  OAI22_X1 DP_mult_215_U1928 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1668), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1669), .ZN(DP_mult_215_n2143)
         );
  AOI221_X1 DP_mult_215_U1927 ( .B1(DP_sw1_6_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_5_), .C2(DP_mult_215_n1563), .A(DP_mult_215_n2143), .ZN(
        DP_mult_215_n2142) );
  XNOR2_X1 DP_mult_215_U1926 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2142), 
        .ZN(DP_mult_215_n2140) );
  INV_X1 DP_mult_215_U1925 ( .A(DP_mult_215_n680), .ZN(DP_mult_215_n2141) );
  OAI222_X1 DP_mult_215_U1924 ( .A1(DP_mult_215_n2139), .A2(DP_mult_215_n2140), 
        .B1(DP_mult_215_n2139), .B2(DP_mult_215_n2141), .C1(DP_mult_215_n2141), 
        .C2(DP_mult_215_n2140), .ZN(DP_mult_215_n2135) );
  INV_X1 DP_mult_215_U1923 ( .A(DP_mult_215_n1391), .ZN(DP_mult_215_n1672) );
  INV_X1 DP_mult_215_U1922 ( .A(DP_sw1_5_), .ZN(DP_mult_215_n1673) );
  OAI22_X1 DP_mult_215_U1921 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1672), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1673), .ZN(DP_mult_215_n2138)
         );
  AOI221_X1 DP_mult_215_U1920 ( .B1(DP_sw1_7_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_6_), .C2(DP_mult_215_n1563), .A(DP_mult_215_n2138), .ZN(
        DP_mult_215_n2137) );
  XNOR2_X1 DP_mult_215_U1919 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2137), 
        .ZN(DP_mult_215_n2136) );
  AOI222_X1 DP_mult_215_U1918 ( .A1(DP_mult_215_n2135), .A2(DP_mult_215_n2136), 
        .B1(DP_mult_215_n2135), .B2(DP_mult_215_n676), .C1(DP_mult_215_n676), 
        .C2(DP_mult_215_n2136), .ZN(DP_mult_215_n2130) );
  INV_X1 DP_mult_215_U1917 ( .A(DP_mult_215_n1390), .ZN(DP_mult_215_n1676) );
  INV_X1 DP_mult_215_U1916 ( .A(DP_sw1_6_), .ZN(DP_mult_215_n1677) );
  OAI22_X1 DP_mult_215_U1915 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1676), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1677), .ZN(DP_mult_215_n2134)
         );
  AOI221_X1 DP_mult_215_U1914 ( .B1(DP_sw1_8_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_7_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2134), .ZN(
        DP_mult_215_n2133) );
  XNOR2_X1 DP_mult_215_U1913 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2133), 
        .ZN(DP_mult_215_n2131) );
  INV_X1 DP_mult_215_U1912 ( .A(DP_mult_215_n672), .ZN(DP_mult_215_n2132) );
  OAI222_X1 DP_mult_215_U1911 ( .A1(DP_mult_215_n2130), .A2(DP_mult_215_n2131), 
        .B1(DP_mult_215_n2130), .B2(DP_mult_215_n2132), .C1(DP_mult_215_n2132), 
        .C2(DP_mult_215_n2131), .ZN(DP_mult_215_n2126) );
  INV_X1 DP_mult_215_U1910 ( .A(DP_mult_215_n1389), .ZN(DP_mult_215_n1680) );
  INV_X1 DP_mult_215_U1909 ( .A(DP_sw1_7_), .ZN(DP_mult_215_n1681) );
  OAI22_X1 DP_mult_215_U1908 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1680), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1681), .ZN(DP_mult_215_n2129)
         );
  AOI221_X1 DP_mult_215_U1907 ( .B1(DP_sw1_9_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_8_), .C2(DP_mult_215_n1563), .A(DP_mult_215_n2129), .ZN(
        DP_mult_215_n2128) );
  XNOR2_X1 DP_mult_215_U1906 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2128), 
        .ZN(DP_mult_215_n2127) );
  AOI222_X1 DP_mult_215_U1905 ( .A1(DP_mult_215_n2126), .A2(DP_mult_215_n2127), 
        .B1(DP_mult_215_n2126), .B2(DP_mult_215_n666), .C1(DP_mult_215_n666), 
        .C2(DP_mult_215_n2127), .ZN(DP_mult_215_n2121) );
  INV_X1 DP_mult_215_U1904 ( .A(DP_mult_215_n1388), .ZN(DP_mult_215_n1684) );
  INV_X1 DP_mult_215_U1903 ( .A(DP_sw1_8_), .ZN(DP_mult_215_n1685) );
  OAI22_X1 DP_mult_215_U1902 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1684), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1685), .ZN(DP_mult_215_n2125)
         );
  AOI221_X1 DP_mult_215_U1901 ( .B1(DP_sw1_10_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_9_), .C2(DP_mult_215_n1563), .A(DP_mult_215_n2125), .ZN(
        DP_mult_215_n2124) );
  XNOR2_X1 DP_mult_215_U1900 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2124), 
        .ZN(DP_mult_215_n2122) );
  INV_X1 DP_mult_215_U1899 ( .A(DP_mult_215_n660), .ZN(DP_mult_215_n2123) );
  OAI222_X1 DP_mult_215_U1898 ( .A1(DP_mult_215_n2121), .A2(DP_mult_215_n2122), 
        .B1(DP_mult_215_n2121), .B2(DP_mult_215_n2123), .C1(DP_mult_215_n2123), 
        .C2(DP_mult_215_n2122), .ZN(DP_mult_215_n2117) );
  INV_X1 DP_mult_215_U1897 ( .A(DP_mult_215_n1387), .ZN(DP_mult_215_n1688) );
  INV_X1 DP_mult_215_U1896 ( .A(DP_sw1_9_), .ZN(DP_mult_215_n1689) );
  OAI22_X1 DP_mult_215_U1895 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1688), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1689), .ZN(DP_mult_215_n2120)
         );
  AOI221_X1 DP_mult_215_U1894 ( .B1(DP_sw1_11_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_10_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2120), .ZN(
        DP_mult_215_n2119) );
  XNOR2_X1 DP_mult_215_U1893 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2119), 
        .ZN(DP_mult_215_n2118) );
  AOI222_X1 DP_mult_215_U1892 ( .A1(DP_mult_215_n2117), .A2(DP_mult_215_n2118), 
        .B1(DP_mult_215_n2117), .B2(DP_mult_215_n654), .C1(DP_mult_215_n654), 
        .C2(DP_mult_215_n2118), .ZN(DP_mult_215_n2112) );
  INV_X1 DP_mult_215_U1891 ( .A(DP_mult_215_n1386), .ZN(DP_mult_215_n1692) );
  INV_X1 DP_mult_215_U1890 ( .A(DP_sw1_10_), .ZN(DP_mult_215_n1693) );
  OAI22_X1 DP_mult_215_U1889 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1692), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1693), .ZN(DP_mult_215_n2116)
         );
  AOI221_X1 DP_mult_215_U1888 ( .B1(DP_sw1_12_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_11_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2116), .ZN(
        DP_mult_215_n2115) );
  XNOR2_X1 DP_mult_215_U1887 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2115), 
        .ZN(DP_mult_215_n2113) );
  INV_X1 DP_mult_215_U1886 ( .A(DP_mult_215_n646), .ZN(DP_mult_215_n2114) );
  OAI222_X1 DP_mult_215_U1885 ( .A1(DP_mult_215_n2112), .A2(DP_mult_215_n2113), 
        .B1(DP_mult_215_n2112), .B2(DP_mult_215_n2114), .C1(DP_mult_215_n2114), 
        .C2(DP_mult_215_n2113), .ZN(DP_mult_215_n2108) );
  INV_X1 DP_mult_215_U1884 ( .A(DP_mult_215_n1385), .ZN(DP_mult_215_n1696) );
  INV_X1 DP_mult_215_U1883 ( .A(DP_sw1_11_), .ZN(DP_mult_215_n1697) );
  OAI22_X1 DP_mult_215_U1882 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1696), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1697), .ZN(DP_mult_215_n2111)
         );
  AOI221_X1 DP_mult_215_U1881 ( .B1(DP_sw1_13_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_12_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2111), .ZN(
        DP_mult_215_n2110) );
  XNOR2_X1 DP_mult_215_U1880 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2110), 
        .ZN(DP_mult_215_n2109) );
  AOI222_X1 DP_mult_215_U1879 ( .A1(DP_mult_215_n2108), .A2(DP_mult_215_n2109), 
        .B1(DP_mult_215_n2108), .B2(DP_mult_215_n638), .C1(DP_mult_215_n638), 
        .C2(DP_mult_215_n2109), .ZN(DP_mult_215_n2103) );
  INV_X1 DP_mult_215_U1878 ( .A(DP_mult_215_n1384), .ZN(DP_mult_215_n1700) );
  INV_X1 DP_mult_215_U1877 ( .A(DP_sw1_12_), .ZN(DP_mult_215_n1701) );
  OAI22_X1 DP_mult_215_U1876 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1700), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1701), .ZN(DP_mult_215_n2107)
         );
  AOI221_X1 DP_mult_215_U1875 ( .B1(DP_sw1_14_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_13_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2107), .ZN(
        DP_mult_215_n2106) );
  XNOR2_X1 DP_mult_215_U1874 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2106), 
        .ZN(DP_mult_215_n2104) );
  INV_X1 DP_mult_215_U1873 ( .A(DP_mult_215_n630), .ZN(DP_mult_215_n2105) );
  OAI222_X1 DP_mult_215_U1872 ( .A1(DP_mult_215_n2103), .A2(DP_mult_215_n2104), 
        .B1(DP_mult_215_n2103), .B2(DP_mult_215_n2105), .C1(DP_mult_215_n2105), 
        .C2(DP_mult_215_n2104), .ZN(DP_mult_215_n2099) );
  INV_X1 DP_mult_215_U1871 ( .A(DP_mult_215_n1383), .ZN(DP_mult_215_n1704) );
  INV_X1 DP_mult_215_U1870 ( .A(DP_sw1_13_), .ZN(DP_mult_215_n1705) );
  OAI22_X1 DP_mult_215_U1869 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1704), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1705), .ZN(DP_mult_215_n2102)
         );
  AOI221_X1 DP_mult_215_U1868 ( .B1(DP_sw1_15_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_14_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2102), .ZN(
        DP_mult_215_n2101) );
  XNOR2_X1 DP_mult_215_U1867 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2101), 
        .ZN(DP_mult_215_n2100) );
  AOI222_X1 DP_mult_215_U1866 ( .A1(DP_mult_215_n2099), .A2(DP_mult_215_n2100), 
        .B1(DP_mult_215_n2099), .B2(DP_mult_215_n620), .C1(DP_mult_215_n620), 
        .C2(DP_mult_215_n2100), .ZN(DP_mult_215_n2094) );
  INV_X1 DP_mult_215_U1865 ( .A(DP_mult_215_n1382), .ZN(DP_mult_215_n1708) );
  INV_X1 DP_mult_215_U1864 ( .A(DP_sw1_14_), .ZN(DP_mult_215_n1709) );
  OAI22_X1 DP_mult_215_U1863 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1708), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1709), .ZN(DP_mult_215_n2098)
         );
  AOI221_X1 DP_mult_215_U1862 ( .B1(DP_sw1_16_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_15_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2098), .ZN(
        DP_mult_215_n2097) );
  XNOR2_X1 DP_mult_215_U1861 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2097), 
        .ZN(DP_mult_215_n2095) );
  INV_X1 DP_mult_215_U1860 ( .A(DP_mult_215_n610), .ZN(DP_mult_215_n2096) );
  OAI222_X1 DP_mult_215_U1859 ( .A1(DP_mult_215_n2094), .A2(DP_mult_215_n2095), 
        .B1(DP_mult_215_n2094), .B2(DP_mult_215_n2096), .C1(DP_mult_215_n2096), 
        .C2(DP_mult_215_n2095), .ZN(DP_mult_215_n2090) );
  INV_X1 DP_mult_215_U1858 ( .A(DP_mult_215_n1381), .ZN(DP_mult_215_n1712) );
  INV_X1 DP_mult_215_U1857 ( .A(DP_sw1_15_), .ZN(DP_mult_215_n1713) );
  OAI22_X1 DP_mult_215_U1856 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1712), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1713), .ZN(DP_mult_215_n2093)
         );
  AOI221_X1 DP_mult_215_U1855 ( .B1(DP_sw1_17_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_16_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2093), .ZN(
        DP_mult_215_n2092) );
  XNOR2_X1 DP_mult_215_U1854 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2092), 
        .ZN(DP_mult_215_n2091) );
  AOI222_X1 DP_mult_215_U1853 ( .A1(DP_mult_215_n2090), .A2(DP_mult_215_n2091), 
        .B1(DP_mult_215_n2090), .B2(DP_mult_215_n600), .C1(DP_mult_215_n600), 
        .C2(DP_mult_215_n2091), .ZN(DP_mult_215_n2085) );
  INV_X1 DP_mult_215_U1852 ( .A(DP_mult_215_n1380), .ZN(DP_mult_215_n1716) );
  INV_X1 DP_mult_215_U1851 ( .A(DP_sw1_16_), .ZN(DP_mult_215_n1717) );
  OAI22_X1 DP_mult_215_U1850 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1716), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1717), .ZN(DP_mult_215_n2089)
         );
  AOI221_X1 DP_mult_215_U1849 ( .B1(DP_sw1_18_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_17_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2089), .ZN(
        DP_mult_215_n2088) );
  XNOR2_X1 DP_mult_215_U1848 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2088), 
        .ZN(DP_mult_215_n2086) );
  INV_X1 DP_mult_215_U1847 ( .A(DP_mult_215_n588), .ZN(DP_mult_215_n2087) );
  OAI222_X1 DP_mult_215_U1846 ( .A1(DP_mult_215_n2085), .A2(DP_mult_215_n2086), 
        .B1(DP_mult_215_n2085), .B2(DP_mult_215_n2087), .C1(DP_mult_215_n2087), 
        .C2(DP_mult_215_n2086), .ZN(DP_mult_215_n2081) );
  INV_X1 DP_mult_215_U1845 ( .A(DP_mult_215_n1379), .ZN(DP_mult_215_n1720) );
  INV_X1 DP_mult_215_U1844 ( .A(DP_sw1_17_), .ZN(DP_mult_215_n1721) );
  OAI22_X1 DP_mult_215_U1843 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1720), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1721), .ZN(DP_mult_215_n2084)
         );
  AOI221_X1 DP_mult_215_U1842 ( .B1(DP_sw1_19_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_18_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2084), .ZN(
        DP_mult_215_n2083) );
  XNOR2_X1 DP_mult_215_U1841 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2083), 
        .ZN(DP_mult_215_n2082) );
  AOI222_X1 DP_mult_215_U1840 ( .A1(DP_mult_215_n2081), .A2(DP_mult_215_n2082), 
        .B1(DP_mult_215_n2081), .B2(DP_mult_215_n576), .C1(DP_mult_215_n576), 
        .C2(DP_mult_215_n2082), .ZN(DP_mult_215_n2080) );
  INV_X1 DP_mult_215_U1839 ( .A(DP_mult_215_n2080), .ZN(DP_mult_215_n2076) );
  INV_X1 DP_mult_215_U1838 ( .A(DP_mult_215_n1378), .ZN(DP_mult_215_n1724) );
  INV_X1 DP_mult_215_U1837 ( .A(DP_sw1_18_), .ZN(DP_mult_215_n1725) );
  OAI22_X1 DP_mult_215_U1836 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1724), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1725), .ZN(DP_mult_215_n2079)
         );
  AOI221_X1 DP_mult_215_U1835 ( .B1(DP_sw1_20_), .B2(DP_mult_215_n1561), .C1(
        DP_sw1_19_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2079), .ZN(
        DP_mult_215_n2078) );
  XNOR2_X1 DP_mult_215_U1834 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n2078), 
        .ZN(DP_mult_215_n2077) );
  AOI222_X1 DP_mult_215_U1833 ( .A1(DP_mult_215_n2076), .A2(DP_mult_215_n2077), 
        .B1(DP_mult_215_n2076), .B2(DP_mult_215_n564), .C1(DP_mult_215_n564), 
        .C2(DP_mult_215_n2077), .ZN(DP_mult_215_n2071) );
  INV_X1 DP_mult_215_U1832 ( .A(DP_mult_215_n1377), .ZN(DP_mult_215_n1728) );
  INV_X1 DP_mult_215_U1831 ( .A(DP_sw1_19_), .ZN(DP_mult_215_n1729) );
  OAI22_X1 DP_mult_215_U1830 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1728), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1729), .ZN(DP_mult_215_n2075)
         );
  AOI221_X1 DP_mult_215_U1829 ( .B1(DP_mult_215_n1561), .B2(DP_sw1_21_), .C1(
        DP_sw1_20_), .C2(DP_mult_215_n1562), .A(DP_mult_215_n2075), .ZN(
        DP_mult_215_n2074) );
  XNOR2_X1 DP_mult_215_U1828 ( .A(DP_mult_215_n1742), .B(DP_mult_215_n2074), 
        .ZN(DP_mult_215_n2072) );
  INV_X1 DP_mult_215_U1827 ( .A(DP_mult_215_n550), .ZN(DP_mult_215_n2073) );
  OAI222_X1 DP_mult_215_U1826 ( .A1(DP_mult_215_n2071), .A2(DP_mult_215_n2072), 
        .B1(DP_mult_215_n2071), .B2(DP_mult_215_n2073), .C1(DP_mult_215_n2073), 
        .C2(DP_mult_215_n2072), .ZN(DP_mult_215_n326) );
  XNOR2_X1 DP_mult_215_U1825 ( .A(DP_coeff_ret1[21]), .B(DP_mult_215_n1608), 
        .ZN(DP_mult_215_n2067) );
  INV_X1 DP_mult_215_U1824 ( .A(DP_mult_215_n2067), .ZN(DP_mult_215_n2070) );
  XNOR2_X1 DP_mult_215_U1823 ( .A(DP_coeff_ret1[21]), .B(DP_coeff_ret1[22]), 
        .ZN(DP_mult_215_n2069) );
  XNOR2_X1 DP_mult_215_U1822 ( .A(DP_coeff_ret1[22]), .B(DP_mult_215_n1611), 
        .ZN(DP_mult_215_n2068) );
  NAND3_X1 DP_mult_215_U1821 ( .A1(DP_mult_215_n2067), .A2(DP_mult_215_n2068), 
        .A3(DP_mult_215_n2069), .ZN(DP_mult_215_n1629) );
  INV_X1 DP_mult_215_U1820 ( .A(DP_sw1_21_), .ZN(DP_mult_215_n1643) );
  OAI22_X1 DP_mult_215_U1819 ( .A1(DP_mult_215_n1548), .A2(DP_mult_215_n1618), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1643), .ZN(DP_mult_215_n2066)
         );
  AOI221_X1 DP_mult_215_U1818 ( .B1(DP_sw1_22_), .B2(DP_mult_215_n1560), .C1(
        DP_mult_215_n1375), .C2(DP_mult_215_n1549), .A(DP_mult_215_n2066), 
        .ZN(DP_mult_215_n2065) );
  XOR2_X1 DP_mult_215_U1817 ( .A(DP_mult_215_n1611), .B(DP_mult_215_n2065), 
        .Z(DP_mult_215_n1627) );
  INV_X1 DP_mult_215_U1816 ( .A(DP_mult_215_n1627), .ZN(DP_mult_215_n351) );
  INV_X1 DP_mult_215_U1815 ( .A(DP_mult_215_n356), .ZN(DP_mult_215_n360) );
  OAI22_X1 DP_mult_215_U1814 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1712), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1713), .ZN(DP_mult_215_n2064)
         );
  AOI221_X1 DP_mult_215_U1813 ( .B1(DP_sw1_17_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_16_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2064), .ZN(
        DP_mult_215_n2063) );
  XOR2_X1 DP_mult_215_U1812 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2063), 
        .Z(DP_mult_215_n374) );
  INV_X1 DP_mult_215_U1811 ( .A(DP_mult_215_n374), .ZN(DP_mult_215_n368) );
  INV_X1 DP_mult_215_U1810 ( .A(DP_mult_215_n387), .ZN(DP_mult_215_n395) );
  OAI22_X1 DP_mult_215_U1809 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1688), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1689), .ZN(DP_mult_215_n2062)
         );
  AOI221_X1 DP_mult_215_U1808 ( .B1(DP_sw1_11_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_10_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2062), .ZN(
        DP_mult_215_n2061) );
  XOR2_X1 DP_mult_215_U1807 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2061), 
        .Z(DP_mult_215_n421) );
  INV_X1 DP_mult_215_U1806 ( .A(DP_mult_215_n421), .ZN(DP_mult_215_n411) );
  OAI22_X1 DP_mult_215_U1805 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1676), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1677), .ZN(DP_mult_215_n2060)
         );
  AOI221_X1 DP_mult_215_U1804 ( .B1(DP_sw1_8_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_7_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2060), .ZN(
        DP_mult_215_n2059) );
  XOR2_X1 DP_mult_215_U1803 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2059), 
        .Z(DP_mult_215_n454) );
  INV_X1 DP_mult_215_U1802 ( .A(DP_mult_215_n454), .ZN(DP_mult_215_n442) );
  OAI21_X1 DP_mult_215_U1801 ( .B1(DP_mult_215_n1561), .B2(DP_mult_215_n1563), 
        .A(DP_mult_215_n1615), .ZN(DP_mult_215_n2058) );
  OAI221_X1 DP_mult_215_U1800 ( .B1(DP_mult_215_n1618), .B2(DP_mult_215_n1639), 
        .C1(DP_mult_215_n1619), .C2(DP_mult_215_n1564), .A(DP_mult_215_n2058), 
        .ZN(DP_mult_215_n2057) );
  XOR2_X1 DP_mult_215_U1799 ( .A(DP_mult_215_n2057), .B(DP_mult_215_n1742), 
        .Z(DP_mult_215_n2056) );
  NOR2_X1 DP_mult_215_U1798 ( .A1(DP_mult_215_n2056), .A2(DP_mult_215_n519), 
        .ZN(DP_mult_215_n493) );
  INV_X1 DP_mult_215_U1797 ( .A(DP_mult_215_n493), .ZN(DP_mult_215_n479) );
  XNOR2_X1 DP_mult_215_U1796 ( .A(DP_mult_215_n519), .B(DP_mult_215_n2056), 
        .ZN(DP_mult_215_n506) );
  INV_X1 DP_mult_215_U1795 ( .A(DP_sw1_20_), .ZN(DP_mult_215_n1640) );
  OAI22_X1 DP_mult_215_U1794 ( .A1(DP_mult_215_n1556), .A2(DP_mult_215_n1640), 
        .B1(DP_mult_215_n1550), .B2(DP_mult_215_n1643), .ZN(DP_mult_215_n2055)
         );
  AOI221_X1 DP_mult_215_U1793 ( .B1(DP_sw1_22_), .B2(DP_mult_215_n1559), .C1(
        DP_mult_215_n1376), .C2(DP_mult_215_n1549), .A(DP_mult_215_n2055), 
        .ZN(DP_mult_215_n2054) );
  XNOR2_X1 DP_mult_215_U1792 ( .A(DP_coeff_ret1[23]), .B(DP_mult_215_n2054), 
        .ZN(DP_mult_215_n729) );
  OAI22_X1 DP_mult_215_U1791 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1728), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1729), .ZN(DP_mult_215_n2053)
         );
  AOI221_X1 DP_mult_215_U1790 ( .B1(DP_sw1_21_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_20_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2053), .ZN(
        DP_mult_215_n2052) );
  XNOR2_X1 DP_mult_215_U1789 ( .A(DP_coeff_ret1[23]), .B(DP_mult_215_n2052), 
        .ZN(DP_mult_215_n730) );
  OAI22_X1 DP_mult_215_U1788 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1724), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1725), .ZN(DP_mult_215_n2051)
         );
  AOI221_X1 DP_mult_215_U1787 ( .B1(DP_sw1_20_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_19_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2051), .ZN(
        DP_mult_215_n2050) );
  XNOR2_X1 DP_mult_215_U1786 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2050), 
        .ZN(DP_mult_215_n731) );
  OAI22_X1 DP_mult_215_U1785 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1720), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1721), .ZN(DP_mult_215_n2049)
         );
  AOI221_X1 DP_mult_215_U1784 ( .B1(DP_sw1_19_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_18_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2049), .ZN(
        DP_mult_215_n2048) );
  XNOR2_X1 DP_mult_215_U1783 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2048), 
        .ZN(DP_mult_215_n732) );
  OAI22_X1 DP_mult_215_U1782 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1716), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1717), .ZN(DP_mult_215_n2047)
         );
  AOI221_X1 DP_mult_215_U1781 ( .B1(DP_sw1_18_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_17_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2047), .ZN(
        DP_mult_215_n2046) );
  XNOR2_X1 DP_mult_215_U1780 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2046), 
        .ZN(DP_mult_215_n733) );
  OAI22_X1 DP_mult_215_U1779 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1708), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1709), .ZN(DP_mult_215_n2045)
         );
  AOI221_X1 DP_mult_215_U1778 ( .B1(DP_sw1_16_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_15_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2045), .ZN(
        DP_mult_215_n2044) );
  XNOR2_X1 DP_mult_215_U1777 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2044), 
        .ZN(DP_mult_215_n734) );
  OAI22_X1 DP_mult_215_U1776 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1704), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1705), .ZN(DP_mult_215_n2043)
         );
  AOI221_X1 DP_mult_215_U1775 ( .B1(DP_sw1_15_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_14_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2043), .ZN(
        DP_mult_215_n2042) );
  XNOR2_X1 DP_mult_215_U1774 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2042), 
        .ZN(DP_mult_215_n735) );
  OAI22_X1 DP_mult_215_U1773 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1700), 
        .B1(DP_mult_215_n1556), .B2(DP_mult_215_n1701), .ZN(DP_mult_215_n2041)
         );
  AOI221_X1 DP_mult_215_U1772 ( .B1(DP_sw1_14_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_13_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2041), .ZN(
        DP_mult_215_n2040) );
  XNOR2_X1 DP_mult_215_U1771 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2040), 
        .ZN(DP_mult_215_n736) );
  OAI22_X1 DP_mult_215_U1770 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1696), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1697), .ZN(DP_mult_215_n2039)
         );
  AOI221_X1 DP_mult_215_U1769 ( .B1(DP_sw1_13_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_12_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2039), .ZN(
        DP_mult_215_n2038) );
  XNOR2_X1 DP_mult_215_U1768 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2038), 
        .ZN(DP_mult_215_n737) );
  OAI22_X1 DP_mult_215_U1767 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1692), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1693), .ZN(DP_mult_215_n2037)
         );
  AOI221_X1 DP_mult_215_U1766 ( .B1(DP_sw1_12_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_11_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2037), .ZN(
        DP_mult_215_n2036) );
  XNOR2_X1 DP_mult_215_U1765 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2036), 
        .ZN(DP_mult_215_n738) );
  OAI22_X1 DP_mult_215_U1764 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1684), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1685), .ZN(DP_mult_215_n2035)
         );
  AOI221_X1 DP_mult_215_U1763 ( .B1(DP_sw1_10_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_9_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2035), .ZN(
        DP_mult_215_n2034) );
  XNOR2_X1 DP_mult_215_U1762 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2034), 
        .ZN(DP_mult_215_n739) );
  OAI22_X1 DP_mult_215_U1761 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1680), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1681), .ZN(DP_mult_215_n2033)
         );
  AOI221_X1 DP_mult_215_U1760 ( .B1(DP_sw1_9_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_8_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2033), .ZN(
        DP_mult_215_n2032) );
  XNOR2_X1 DP_mult_215_U1759 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2032), 
        .ZN(DP_mult_215_n740) );
  OAI22_X1 DP_mult_215_U1758 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1672), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1673), .ZN(DP_mult_215_n2031)
         );
  AOI221_X1 DP_mult_215_U1757 ( .B1(DP_sw1_7_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_6_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2031), .ZN(
        DP_mult_215_n2030) );
  XNOR2_X1 DP_mult_215_U1756 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2030), 
        .ZN(DP_mult_215_n741) );
  OAI22_X1 DP_mult_215_U1755 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1668), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1669), .ZN(DP_mult_215_n2029)
         );
  AOI221_X1 DP_mult_215_U1754 ( .B1(DP_sw1_6_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_5_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2029), .ZN(
        DP_mult_215_n2028) );
  XNOR2_X1 DP_mult_215_U1753 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2028), 
        .ZN(DP_mult_215_n742) );
  OAI22_X1 DP_mult_215_U1752 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1664), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1665), .ZN(DP_mult_215_n2027)
         );
  AOI221_X1 DP_mult_215_U1751 ( .B1(DP_sw1_5_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_4_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2027), .ZN(
        DP_mult_215_n2026) );
  XNOR2_X1 DP_mult_215_U1750 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2026), 
        .ZN(DP_mult_215_n743) );
  OAI22_X1 DP_mult_215_U1749 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1660), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1661), .ZN(DP_mult_215_n2025)
         );
  AOI221_X1 DP_mult_215_U1748 ( .B1(DP_sw1_4_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_3_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2025), .ZN(
        DP_mult_215_n2024) );
  XNOR2_X1 DP_mult_215_U1747 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2024), 
        .ZN(DP_mult_215_n744) );
  OAI22_X1 DP_mult_215_U1746 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1657), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1649), .ZN(DP_mult_215_n2023)
         );
  AOI221_X1 DP_mult_215_U1745 ( .B1(DP_sw1_3_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_2_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2023), .ZN(
        DP_mult_215_n2022) );
  XNOR2_X1 DP_mult_215_U1744 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2022), 
        .ZN(DP_mult_215_n745) );
  INV_X1 DP_mult_215_U1743 ( .A(DP_mult_215_n1396), .ZN(DP_mult_215_n1653) );
  INV_X1 DP_mult_215_U1742 ( .A(DP_sw1_0_), .ZN(DP_mult_215_n1647) );
  OAI22_X1 DP_mult_215_U1741 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1653), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1567), .ZN(DP_mult_215_n2021)
         );
  AOI221_X1 DP_mult_215_U1740 ( .B1(DP_sw1_2_), .B2(DP_mult_215_n1559), .C1(
        DP_sw1_1_), .C2(DP_mult_215_n1560), .A(DP_mult_215_n2021), .ZN(
        DP_mult_215_n2020) );
  XNOR2_X1 DP_mult_215_U1739 ( .A(DP_mult_215_n1610), .B(DP_mult_215_n2020), 
        .ZN(DP_mult_215_n746) );
  OAI222_X1 DP_mult_215_U1738 ( .A1(DP_mult_215_n1548), .A2(DP_mult_215_n1649), 
        .B1(DP_mult_215_n1550), .B2(DP_mult_215_n1566), .C1(DP_mult_215_n1558), 
        .C2(DP_mult_215_n1650), .ZN(DP_mult_215_n2019) );
  XNOR2_X1 DP_mult_215_U1737 ( .A(DP_mult_215_n2019), .B(DP_mult_215_n1611), 
        .ZN(DP_mult_215_n747) );
  OAI22_X1 DP_mult_215_U1736 ( .A1(DP_mult_215_n1548), .A2(DP_mult_215_n1567), 
        .B1(DP_mult_215_n1558), .B2(DP_mult_215_n1567), .ZN(DP_mult_215_n2018)
         );
  XNOR2_X1 DP_mult_215_U1735 ( .A(DP_mult_215_n2018), .B(DP_mult_215_n1611), 
        .ZN(DP_mult_215_n748) );
  XOR2_X1 DP_mult_215_U1734 ( .A(DP_coeff_ret1[18]), .B(DP_mult_215_n1607), 
        .Z(DP_mult_215_n2017) );
  XOR2_X1 DP_mult_215_U1733 ( .A(DP_coeff_ret1[19]), .B(DP_mult_215_n1608), 
        .Z(DP_mult_215_n2016) );
  XNOR2_X1 DP_mult_215_U1732 ( .A(DP_coeff_ret1[18]), .B(DP_coeff_ret1[19]), 
        .ZN(DP_mult_215_n2015) );
  NAND3_X1 DP_mult_215_U1731 ( .A1(DP_mult_215_n2017), .A2(DP_mult_215_n2016), 
        .A3(DP_mult_215_n2015), .ZN(DP_mult_215_n1967) );
  INV_X1 DP_mult_215_U1730 ( .A(DP_mult_215_n2017), .ZN(DP_mult_215_n2014) );
  OAI21_X1 DP_mult_215_U1729 ( .B1(DP_mult_215_n1594), .B2(DP_mult_215_n1595), 
        .A(DP_mult_215_n1615), .ZN(DP_mult_215_n2013) );
  OAI221_X1 DP_mult_215_U1728 ( .B1(DP_mult_215_n1617), .B2(DP_mult_215_n1597), 
        .C1(DP_mult_215_n1619), .C2(DP_mult_215_n1593), .A(DP_mult_215_n2013), 
        .ZN(DP_mult_215_n2012) );
  XNOR2_X1 DP_mult_215_U1727 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n2012), 
        .ZN(DP_mult_215_n749) );
  INV_X1 DP_mult_215_U1726 ( .A(DP_mult_215_n1374), .ZN(DP_mult_215_n1633) );
  INV_X1 DP_mult_215_U1725 ( .A(DP_sw1_22_), .ZN(DP_mult_215_n1634) );
  OAI22_X1 DP_mult_215_U1724 ( .A1(DP_mult_215_n1633), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1634), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n2011)
         );
  AOI221_X1 DP_mult_215_U1723 ( .B1(DP_mult_215_n1594), .B2(DP_mult_215_n1614), 
        .C1(DP_mult_215_n1595), .C2(DP_mult_215_n1615), .A(DP_mult_215_n2011), 
        .ZN(DP_mult_215_n2010) );
  XNOR2_X1 DP_mult_215_U1722 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n2010), 
        .ZN(DP_mult_215_n750) );
  OAI22_X1 DP_mult_215_U1721 ( .A1(DP_mult_215_n1620), .A2(DP_mult_215_n1541), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n2009)
         );
  AOI221_X1 DP_mult_215_U1720 ( .B1(DP_mult_215_n1595), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1542), .C2(DP_mult_215_n1375), .A(DP_mult_215_n2009), 
        .ZN(DP_mult_215_n2008) );
  XNOR2_X1 DP_mult_215_U1719 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n2008), 
        .ZN(DP_mult_215_n751) );
  OAI22_X1 DP_mult_215_U1718 ( .A1(DP_mult_215_n1640), .A2(DP_mult_215_n1597), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1543), .ZN(DP_mult_215_n2007)
         );
  AOI221_X1 DP_mult_215_U1717 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1542), .C2(DP_mult_215_n1376), .A(DP_mult_215_n2007), 
        .ZN(DP_mult_215_n2006) );
  XNOR2_X1 DP_mult_215_U1716 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n2006), 
        .ZN(DP_mult_215_n752) );
  OAI22_X1 DP_mult_215_U1715 ( .A1(DP_mult_215_n1728), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1729), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n2005)
         );
  AOI221_X1 DP_mult_215_U1714 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_21_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_20_), .A(DP_mult_215_n2005), .ZN(
        DP_mult_215_n2004) );
  XNOR2_X1 DP_mult_215_U1713 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n2004), 
        .ZN(DP_mult_215_n753) );
  OAI22_X1 DP_mult_215_U1712 ( .A1(DP_mult_215_n1724), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1725), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n2003)
         );
  AOI221_X1 DP_mult_215_U1711 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_20_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_19_), .A(DP_mult_215_n2003), .ZN(
        DP_mult_215_n2002) );
  XNOR2_X1 DP_mult_215_U1710 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n2002), 
        .ZN(DP_mult_215_n754) );
  OAI22_X1 DP_mult_215_U1709 ( .A1(DP_mult_215_n1720), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1721), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n2001)
         );
  AOI221_X1 DP_mult_215_U1708 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_19_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_18_), .A(DP_mult_215_n2001), .ZN(
        DP_mult_215_n2000) );
  XNOR2_X1 DP_mult_215_U1707 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n2000), 
        .ZN(DP_mult_215_n755) );
  OAI22_X1 DP_mult_215_U1706 ( .A1(DP_mult_215_n1716), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1717), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n1999)
         );
  AOI221_X1 DP_mult_215_U1705 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_18_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_17_), .A(DP_mult_215_n1999), .ZN(
        DP_mult_215_n1998) );
  XNOR2_X1 DP_mult_215_U1704 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n1998), 
        .ZN(DP_mult_215_n756) );
  OAI22_X1 DP_mult_215_U1703 ( .A1(DP_mult_215_n1712), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1713), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n1997)
         );
  AOI221_X1 DP_mult_215_U1702 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_17_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_16_), .A(DP_mult_215_n1997), .ZN(
        DP_mult_215_n1996) );
  XNOR2_X1 DP_mult_215_U1701 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n1996), 
        .ZN(DP_mult_215_n757) );
  OAI22_X1 DP_mult_215_U1700 ( .A1(DP_mult_215_n1708), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1709), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n1995)
         );
  AOI221_X1 DP_mult_215_U1699 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_16_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_15_), .A(DP_mult_215_n1995), .ZN(
        DP_mult_215_n1994) );
  XNOR2_X1 DP_mult_215_U1698 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n1994), 
        .ZN(DP_mult_215_n758) );
  OAI22_X1 DP_mult_215_U1697 ( .A1(DP_mult_215_n1704), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1705), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n1993)
         );
  AOI221_X1 DP_mult_215_U1696 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_15_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_14_), .A(DP_mult_215_n1993), .ZN(
        DP_mult_215_n1992) );
  XNOR2_X1 DP_mult_215_U1695 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n1992), 
        .ZN(DP_mult_215_n759) );
  OAI22_X1 DP_mult_215_U1694 ( .A1(DP_mult_215_n1700), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1701), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n1991)
         );
  AOI221_X1 DP_mult_215_U1693 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_14_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_13_), .A(DP_mult_215_n1991), .ZN(
        DP_mult_215_n1990) );
  XNOR2_X1 DP_mult_215_U1692 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n1990), 
        .ZN(DP_mult_215_n760) );
  OAI22_X1 DP_mult_215_U1691 ( .A1(DP_mult_215_n1696), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1697), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n1989)
         );
  AOI221_X1 DP_mult_215_U1690 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_13_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_12_), .A(DP_mult_215_n1989), .ZN(
        DP_mult_215_n1988) );
  XNOR2_X1 DP_mult_215_U1689 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n1988), 
        .ZN(DP_mult_215_n761) );
  OAI22_X1 DP_mult_215_U1688 ( .A1(DP_mult_215_n1692), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1693), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1987)
         );
  AOI221_X1 DP_mult_215_U1687 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_12_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_11_), .A(DP_mult_215_n1987), .ZN(
        DP_mult_215_n1986) );
  XNOR2_X1 DP_mult_215_U1686 ( .A(DP_mult_215_n1609), .B(DP_mult_215_n1986), 
        .ZN(DP_mult_215_n762) );
  OAI22_X1 DP_mult_215_U1685 ( .A1(DP_mult_215_n1688), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1689), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1985)
         );
  AOI221_X1 DP_mult_215_U1684 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_11_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_10_), .A(DP_mult_215_n1985), .ZN(
        DP_mult_215_n1984) );
  XNOR2_X1 DP_mult_215_U1683 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1984), 
        .ZN(DP_mult_215_n763) );
  OAI22_X1 DP_mult_215_U1682 ( .A1(DP_mult_215_n1684), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1685), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1983)
         );
  AOI221_X1 DP_mult_215_U1681 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_10_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_9_), .A(DP_mult_215_n1983), .ZN(
        DP_mult_215_n1982) );
  XNOR2_X1 DP_mult_215_U1680 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1982), 
        .ZN(DP_mult_215_n764) );
  OAI22_X1 DP_mult_215_U1679 ( .A1(DP_mult_215_n1680), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1681), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1981)
         );
  AOI221_X1 DP_mult_215_U1678 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_9_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_8_), .A(DP_mult_215_n1981), .ZN(
        DP_mult_215_n1980) );
  XNOR2_X1 DP_mult_215_U1677 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1980), 
        .ZN(DP_mult_215_n765) );
  OAI22_X1 DP_mult_215_U1676 ( .A1(DP_mult_215_n1676), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1677), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1979)
         );
  AOI221_X1 DP_mult_215_U1675 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_8_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_7_), .A(DP_mult_215_n1979), .ZN(
        DP_mult_215_n1978) );
  XNOR2_X1 DP_mult_215_U1674 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1978), 
        .ZN(DP_mult_215_n766) );
  OAI22_X1 DP_mult_215_U1673 ( .A1(DP_mult_215_n1672), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1673), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1977)
         );
  AOI221_X1 DP_mult_215_U1672 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_7_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_6_), .A(DP_mult_215_n1977), .ZN(
        DP_mult_215_n1976) );
  XNOR2_X1 DP_mult_215_U1671 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1976), 
        .ZN(DP_mult_215_n767) );
  OAI22_X1 DP_mult_215_U1670 ( .A1(DP_mult_215_n1668), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1669), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1975)
         );
  AOI221_X1 DP_mult_215_U1669 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_6_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_5_), .A(DP_mult_215_n1975), .ZN(
        DP_mult_215_n1974) );
  XNOR2_X1 DP_mult_215_U1668 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1974), 
        .ZN(DP_mult_215_n768) );
  OAI22_X1 DP_mult_215_U1667 ( .A1(DP_mult_215_n1664), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1665), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1973)
         );
  AOI221_X1 DP_mult_215_U1666 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_5_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_4_), .A(DP_mult_215_n1973), .ZN(
        DP_mult_215_n1972) );
  XNOR2_X1 DP_mult_215_U1665 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1972), 
        .ZN(DP_mult_215_n769) );
  OAI22_X1 DP_mult_215_U1664 ( .A1(DP_mult_215_n1660), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1661), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1971)
         );
  AOI221_X1 DP_mult_215_U1663 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_4_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_3_), .A(DP_mult_215_n1971), .ZN(
        DP_mult_215_n1970) );
  XNOR2_X1 DP_mult_215_U1662 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1970), 
        .ZN(DP_mult_215_n770) );
  OAI22_X1 DP_mult_215_U1661 ( .A1(DP_mult_215_n1657), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1649), .B2(DP_mult_215_n1597), .ZN(DP_mult_215_n1969)
         );
  AOI221_X1 DP_mult_215_U1660 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_3_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_2_), .A(DP_mult_215_n1969), .ZN(
        DP_mult_215_n1968) );
  XNOR2_X1 DP_mult_215_U1659 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1968), 
        .ZN(DP_mult_215_n771) );
  OAI22_X1 DP_mult_215_U1658 ( .A1(DP_mult_215_n1653), .A2(DP_mult_215_n1593), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1596), .ZN(DP_mult_215_n1966)
         );
  AOI221_X1 DP_mult_215_U1657 ( .B1(DP_mult_215_n1594), .B2(DP_sw1_2_), .C1(
        DP_mult_215_n1595), .C2(DP_sw1_1_), .A(DP_mult_215_n1966), .ZN(
        DP_mult_215_n1965) );
  XNOR2_X1 DP_mult_215_U1656 ( .A(DP_mult_215_n1608), .B(DP_mult_215_n1965), 
        .ZN(DP_mult_215_n772) );
  OAI222_X1 DP_mult_215_U1655 ( .A1(DP_mult_215_n1649), .A2(DP_mult_215_n1541), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1543), .C1(DP_mult_215_n1650), 
        .C2(DP_mult_215_n1593), .ZN(DP_mult_215_n1964) );
  XOR2_X1 DP_mult_215_U1654 ( .A(DP_mult_215_n1964), .B(DP_mult_215_n1608), 
        .Z(DP_mult_215_n773) );
  OAI22_X1 DP_mult_215_U1653 ( .A1(DP_mult_215_n1565), .A2(DP_mult_215_n1541), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1593), .ZN(DP_mult_215_n1963)
         );
  XOR2_X1 DP_mult_215_U1652 ( .A(DP_mult_215_n1963), .B(DP_mult_215_n1608), 
        .Z(DP_mult_215_n774) );
  XOR2_X1 DP_mult_215_U1651 ( .A(DP_coeff_ret1[15]), .B(DP_mult_215_n1605), 
        .Z(DP_mult_215_n1962) );
  XNOR2_X1 DP_mult_215_U1650 ( .A(DP_coeff_ret1[16]), .B(DP_mult_215_n1607), 
        .ZN(DP_mult_215_n1961) );
  XNOR2_X1 DP_mult_215_U1649 ( .A(DP_coeff_ret1[15]), .B(DP_coeff_ret1[16]), 
        .ZN(DP_mult_215_n1960) );
  NAND3_X1 DP_mult_215_U1648 ( .A1(DP_mult_215_n1962), .A2(DP_mult_215_n1961), 
        .A3(DP_mult_215_n1960), .ZN(DP_mult_215_n1912) );
  INV_X1 DP_mult_215_U1647 ( .A(DP_mult_215_n1962), .ZN(DP_mult_215_n1959) );
  OAI21_X1 DP_mult_215_U1646 ( .B1(DP_mult_215_n1589), .B2(DP_mult_215_n1590), 
        .A(DP_mult_215_n1615), .ZN(DP_mult_215_n1958) );
  OAI221_X1 DP_mult_215_U1645 ( .B1(DP_mult_215_n1618), .B2(DP_mult_215_n1592), 
        .C1(DP_mult_215_n1617), .C2(DP_mult_215_n1588), .A(DP_mult_215_n1958), 
        .ZN(DP_mult_215_n1957) );
  XNOR2_X1 DP_mult_215_U1644 ( .A(DP_coeff_ret1[17]), .B(DP_mult_215_n1957), 
        .ZN(DP_mult_215_n775) );
  OAI22_X1 DP_mult_215_U1643 ( .A1(DP_mult_215_n1633), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1634), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1956)
         );
  AOI221_X1 DP_mult_215_U1642 ( .B1(DP_mult_215_n1589), .B2(DP_mult_215_n1613), 
        .C1(DP_mult_215_n1590), .C2(DP_mult_215_n1615), .A(DP_mult_215_n1956), 
        .ZN(DP_mult_215_n1955) );
  XNOR2_X1 DP_mult_215_U1641 ( .A(DP_coeff_ret1[17]), .B(DP_mult_215_n1955), 
        .ZN(DP_mult_215_n776) );
  OAI22_X1 DP_mult_215_U1640 ( .A1(DP_mult_215_n1620), .A2(DP_mult_215_n1534), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1954)
         );
  AOI221_X1 DP_mult_215_U1639 ( .B1(DP_mult_215_n1590), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1537), .C2(DP_mult_215_n1375), .A(DP_mult_215_n1954), 
        .ZN(DP_mult_215_n1953) );
  XNOR2_X1 DP_mult_215_U1638 ( .A(DP_coeff_ret1[17]), .B(DP_mult_215_n1953), 
        .ZN(DP_mult_215_n777) );
  OAI22_X1 DP_mult_215_U1637 ( .A1(DP_mult_215_n1640), .A2(DP_mult_215_n1592), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1540), .ZN(DP_mult_215_n1952)
         );
  AOI221_X1 DP_mult_215_U1636 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1537), .C2(DP_mult_215_n1376), .A(DP_mult_215_n1952), 
        .ZN(DP_mult_215_n1951) );
  XNOR2_X1 DP_mult_215_U1635 ( .A(DP_coeff_ret1[17]), .B(DP_mult_215_n1951), 
        .ZN(DP_mult_215_n778) );
  OAI22_X1 DP_mult_215_U1634 ( .A1(DP_mult_215_n1728), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1729), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1950)
         );
  AOI221_X1 DP_mult_215_U1633 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_21_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_20_), .A(DP_mult_215_n1950), .ZN(
        DP_mult_215_n1949) );
  XNOR2_X1 DP_mult_215_U1632 ( .A(DP_coeff_ret1[17]), .B(DP_mult_215_n1949), 
        .ZN(DP_mult_215_n779) );
  OAI22_X1 DP_mult_215_U1631 ( .A1(DP_mult_215_n1724), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1725), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1948)
         );
  AOI221_X1 DP_mult_215_U1630 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_20_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_19_), .A(DP_mult_215_n1948), .ZN(
        DP_mult_215_n1947) );
  XNOR2_X1 DP_mult_215_U1629 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1947), 
        .ZN(DP_mult_215_n780) );
  OAI22_X1 DP_mult_215_U1628 ( .A1(DP_mult_215_n1720), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1721), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1946)
         );
  AOI221_X1 DP_mult_215_U1627 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_19_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_18_), .A(DP_mult_215_n1946), .ZN(
        DP_mult_215_n1945) );
  XNOR2_X1 DP_mult_215_U1626 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1945), 
        .ZN(DP_mult_215_n781) );
  OAI22_X1 DP_mult_215_U1625 ( .A1(DP_mult_215_n1716), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1717), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1944)
         );
  AOI221_X1 DP_mult_215_U1624 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_18_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_17_), .A(DP_mult_215_n1944), .ZN(
        DP_mult_215_n1943) );
  XNOR2_X1 DP_mult_215_U1623 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1943), 
        .ZN(DP_mult_215_n782) );
  OAI22_X1 DP_mult_215_U1622 ( .A1(DP_mult_215_n1712), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1713), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1942)
         );
  AOI221_X1 DP_mult_215_U1621 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_17_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_16_), .A(DP_mult_215_n1942), .ZN(
        DP_mult_215_n1941) );
  XNOR2_X1 DP_mult_215_U1620 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1941), 
        .ZN(DP_mult_215_n783) );
  OAI22_X1 DP_mult_215_U1619 ( .A1(DP_mult_215_n1708), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1709), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1940)
         );
  AOI221_X1 DP_mult_215_U1618 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_16_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_15_), .A(DP_mult_215_n1940), .ZN(
        DP_mult_215_n1939) );
  XNOR2_X1 DP_mult_215_U1617 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1939), 
        .ZN(DP_mult_215_n784) );
  OAI22_X1 DP_mult_215_U1616 ( .A1(DP_mult_215_n1704), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1705), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1938)
         );
  AOI221_X1 DP_mult_215_U1615 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_15_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_14_), .A(DP_mult_215_n1938), .ZN(
        DP_mult_215_n1937) );
  XNOR2_X1 DP_mult_215_U1614 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1937), 
        .ZN(DP_mult_215_n785) );
  OAI22_X1 DP_mult_215_U1613 ( .A1(DP_mult_215_n1700), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1701), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1936)
         );
  AOI221_X1 DP_mult_215_U1612 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_14_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_13_), .A(DP_mult_215_n1936), .ZN(
        DP_mult_215_n1935) );
  XNOR2_X1 DP_mult_215_U1611 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1935), 
        .ZN(DP_mult_215_n786) );
  OAI22_X1 DP_mult_215_U1610 ( .A1(DP_mult_215_n1696), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1697), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1934)
         );
  AOI221_X1 DP_mult_215_U1609 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_13_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_12_), .A(DP_mult_215_n1934), .ZN(
        DP_mult_215_n1933) );
  XNOR2_X1 DP_mult_215_U1608 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1933), 
        .ZN(DP_mult_215_n787) );
  OAI22_X1 DP_mult_215_U1607 ( .A1(DP_mult_215_n1692), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1693), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1932)
         );
  AOI221_X1 DP_mult_215_U1606 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_12_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_11_), .A(DP_mult_215_n1932), .ZN(
        DP_mult_215_n1931) );
  XNOR2_X1 DP_mult_215_U1605 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1931), 
        .ZN(DP_mult_215_n788) );
  OAI22_X1 DP_mult_215_U1604 ( .A1(DP_mult_215_n1688), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1689), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1930)
         );
  AOI221_X1 DP_mult_215_U1603 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_11_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_10_), .A(DP_mult_215_n1930), .ZN(
        DP_mult_215_n1929) );
  XNOR2_X1 DP_mult_215_U1602 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1929), 
        .ZN(DP_mult_215_n789) );
  OAI22_X1 DP_mult_215_U1601 ( .A1(DP_mult_215_n1684), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1685), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1928)
         );
  AOI221_X1 DP_mult_215_U1600 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_10_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_9_), .A(DP_mult_215_n1928), .ZN(
        DP_mult_215_n1927) );
  XNOR2_X1 DP_mult_215_U1599 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1927), 
        .ZN(DP_mult_215_n790) );
  OAI22_X1 DP_mult_215_U1598 ( .A1(DP_mult_215_n1680), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1681), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1926)
         );
  AOI221_X1 DP_mult_215_U1597 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_9_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_8_), .A(DP_mult_215_n1926), .ZN(
        DP_mult_215_n1925) );
  XNOR2_X1 DP_mult_215_U1596 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1925), 
        .ZN(DP_mult_215_n791) );
  OAI22_X1 DP_mult_215_U1595 ( .A1(DP_mult_215_n1676), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1677), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1924)
         );
  AOI221_X1 DP_mult_215_U1594 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_8_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_7_), .A(DP_mult_215_n1924), .ZN(
        DP_mult_215_n1923) );
  XNOR2_X1 DP_mult_215_U1593 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1923), 
        .ZN(DP_mult_215_n792) );
  OAI22_X1 DP_mult_215_U1592 ( .A1(DP_mult_215_n1672), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1673), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1922)
         );
  AOI221_X1 DP_mult_215_U1591 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_7_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_6_), .A(DP_mult_215_n1922), .ZN(
        DP_mult_215_n1921) );
  XNOR2_X1 DP_mult_215_U1590 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1921), 
        .ZN(DP_mult_215_n793) );
  OAI22_X1 DP_mult_215_U1589 ( .A1(DP_mult_215_n1668), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1669), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1920)
         );
  AOI221_X1 DP_mult_215_U1588 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_6_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_5_), .A(DP_mult_215_n1920), .ZN(
        DP_mult_215_n1919) );
  XNOR2_X1 DP_mult_215_U1587 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1919), 
        .ZN(DP_mult_215_n794) );
  OAI22_X1 DP_mult_215_U1586 ( .A1(DP_mult_215_n1664), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1665), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1918)
         );
  AOI221_X1 DP_mult_215_U1585 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_5_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_4_), .A(DP_mult_215_n1918), .ZN(
        DP_mult_215_n1917) );
  XNOR2_X1 DP_mult_215_U1584 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1917), 
        .ZN(DP_mult_215_n795) );
  OAI22_X1 DP_mult_215_U1583 ( .A1(DP_mult_215_n1660), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1661), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1916)
         );
  AOI221_X1 DP_mult_215_U1582 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_4_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_3_), .A(DP_mult_215_n1916), .ZN(
        DP_mult_215_n1915) );
  XNOR2_X1 DP_mult_215_U1581 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1915), 
        .ZN(DP_mult_215_n796) );
  OAI22_X1 DP_mult_215_U1580 ( .A1(DP_mult_215_n1657), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1649), .B2(DP_mult_215_n1592), .ZN(DP_mult_215_n1914)
         );
  AOI221_X1 DP_mult_215_U1579 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_3_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_2_), .A(DP_mult_215_n1914), .ZN(
        DP_mult_215_n1913) );
  XNOR2_X1 DP_mult_215_U1578 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1913), 
        .ZN(DP_mult_215_n797) );
  OAI22_X1 DP_mult_215_U1577 ( .A1(DP_mult_215_n1653), .A2(DP_mult_215_n1588), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1591), .ZN(DP_mult_215_n1911)
         );
  AOI221_X1 DP_mult_215_U1576 ( .B1(DP_mult_215_n1589), .B2(DP_sw1_2_), .C1(
        DP_mult_215_n1590), .C2(DP_sw1_1_), .A(DP_mult_215_n1911), .ZN(
        DP_mult_215_n1910) );
  XNOR2_X1 DP_mult_215_U1575 ( .A(DP_mult_215_n1606), .B(DP_mult_215_n1910), 
        .ZN(DP_mult_215_n798) );
  OAI222_X1 DP_mult_215_U1574 ( .A1(DP_mult_215_n1649), .A2(DP_mult_215_n1534), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1540), .C1(DP_mult_215_n1650), 
        .C2(DP_mult_215_n1588), .ZN(DP_mult_215_n1909) );
  XNOR2_X1 DP_mult_215_U1573 ( .A(DP_mult_215_n1909), .B(DP_mult_215_n1607), 
        .ZN(DP_mult_215_n799) );
  OAI22_X1 DP_mult_215_U1572 ( .A1(DP_mult_215_n1565), .A2(DP_mult_215_n1534), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1588), .ZN(DP_mult_215_n1908)
         );
  XNOR2_X1 DP_mult_215_U1571 ( .A(DP_mult_215_n1908), .B(DP_mult_215_n1607), 
        .ZN(DP_mult_215_n800) );
  XOR2_X1 DP_mult_215_U1570 ( .A(DP_coeff_ret1[12]), .B(DP_mult_215_n1603), 
        .Z(DP_mult_215_n1907) );
  XNOR2_X1 DP_mult_215_U1569 ( .A(DP_coeff_ret1[13]), .B(DP_mult_215_n1605), 
        .ZN(DP_mult_215_n1906) );
  XNOR2_X1 DP_mult_215_U1568 ( .A(DP_coeff_ret1[12]), .B(DP_coeff_ret1[13]), 
        .ZN(DP_mult_215_n1905) );
  NAND3_X1 DP_mult_215_U1567 ( .A1(DP_mult_215_n1907), .A2(DP_mult_215_n1906), 
        .A3(DP_mult_215_n1905), .ZN(DP_mult_215_n1857) );
  INV_X1 DP_mult_215_U1566 ( .A(DP_mult_215_n1907), .ZN(DP_mult_215_n1904) );
  OAI21_X1 DP_mult_215_U1565 ( .B1(DP_mult_215_n1584), .B2(DP_mult_215_n1585), 
        .A(DP_mult_215_n1615), .ZN(DP_mult_215_n1903) );
  OAI221_X1 DP_mult_215_U1564 ( .B1(DP_mult_215_n1620), .B2(DP_mult_215_n1587), 
        .C1(DP_mult_215_n1619), .C2(DP_mult_215_n1583), .A(DP_mult_215_n1903), 
        .ZN(DP_mult_215_n1902) );
  XNOR2_X1 DP_mult_215_U1563 ( .A(DP_coeff_ret1[14]), .B(DP_mult_215_n1902), 
        .ZN(DP_mult_215_n801) );
  OAI22_X1 DP_mult_215_U1562 ( .A1(DP_mult_215_n1633), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1634), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1901)
         );
  AOI221_X1 DP_mult_215_U1561 ( .B1(DP_mult_215_n1584), .B2(DP_mult_215_n1615), 
        .C1(DP_mult_215_n1585), .C2(DP_mult_215_n1615), .A(DP_mult_215_n1901), 
        .ZN(DP_mult_215_n1900) );
  XNOR2_X1 DP_mult_215_U1560 ( .A(DP_coeff_ret1[14]), .B(DP_mult_215_n1900), 
        .ZN(DP_mult_215_n802) );
  OAI22_X1 DP_mult_215_U1559 ( .A1(DP_mult_215_n1617), .A2(DP_mult_215_n1533), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1899)
         );
  AOI221_X1 DP_mult_215_U1558 ( .B1(DP_mult_215_n1585), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1536), .C2(DP_mult_215_n1375), .A(DP_mult_215_n1899), 
        .ZN(DP_mult_215_n1898) );
  XNOR2_X1 DP_mult_215_U1557 ( .A(DP_coeff_ret1[14]), .B(DP_mult_215_n1898), 
        .ZN(DP_mult_215_n803) );
  OAI22_X1 DP_mult_215_U1556 ( .A1(DP_mult_215_n1640), .A2(DP_mult_215_n1587), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1539), .ZN(DP_mult_215_n1897)
         );
  AOI221_X1 DP_mult_215_U1555 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1536), .C2(DP_mult_215_n1376), .A(DP_mult_215_n1897), 
        .ZN(DP_mult_215_n1896) );
  XNOR2_X1 DP_mult_215_U1554 ( .A(DP_coeff_ret1[14]), .B(DP_mult_215_n1896), 
        .ZN(DP_mult_215_n804) );
  OAI22_X1 DP_mult_215_U1553 ( .A1(DP_mult_215_n1728), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1729), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1895)
         );
  AOI221_X1 DP_mult_215_U1552 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_21_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_20_), .A(DP_mult_215_n1895), .ZN(
        DP_mult_215_n1894) );
  XNOR2_X1 DP_mult_215_U1551 ( .A(DP_coeff_ret1[14]), .B(DP_mult_215_n1894), 
        .ZN(DP_mult_215_n805) );
  OAI22_X1 DP_mult_215_U1550 ( .A1(DP_mult_215_n1724), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1725), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1893)
         );
  AOI221_X1 DP_mult_215_U1549 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_20_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_19_), .A(DP_mult_215_n1893), .ZN(
        DP_mult_215_n1892) );
  XNOR2_X1 DP_mult_215_U1548 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1892), 
        .ZN(DP_mult_215_n806) );
  OAI22_X1 DP_mult_215_U1547 ( .A1(DP_mult_215_n1720), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1721), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1891)
         );
  AOI221_X1 DP_mult_215_U1546 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_19_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_18_), .A(DP_mult_215_n1891), .ZN(
        DP_mult_215_n1890) );
  XNOR2_X1 DP_mult_215_U1545 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1890), 
        .ZN(DP_mult_215_n807) );
  OAI22_X1 DP_mult_215_U1544 ( .A1(DP_mult_215_n1716), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1717), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1889)
         );
  AOI221_X1 DP_mult_215_U1543 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_18_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_17_), .A(DP_mult_215_n1889), .ZN(
        DP_mult_215_n1888) );
  XNOR2_X1 DP_mult_215_U1542 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1888), 
        .ZN(DP_mult_215_n808) );
  OAI22_X1 DP_mult_215_U1541 ( .A1(DP_mult_215_n1712), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1713), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1887)
         );
  AOI221_X1 DP_mult_215_U1540 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_17_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_16_), .A(DP_mult_215_n1887), .ZN(
        DP_mult_215_n1886) );
  XNOR2_X1 DP_mult_215_U1539 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1886), 
        .ZN(DP_mult_215_n809) );
  OAI22_X1 DP_mult_215_U1538 ( .A1(DP_mult_215_n1708), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1709), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1885)
         );
  AOI221_X1 DP_mult_215_U1537 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_16_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_15_), .A(DP_mult_215_n1885), .ZN(
        DP_mult_215_n1884) );
  XNOR2_X1 DP_mult_215_U1536 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1884), 
        .ZN(DP_mult_215_n810) );
  OAI22_X1 DP_mult_215_U1535 ( .A1(DP_mult_215_n1704), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1705), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1883)
         );
  AOI221_X1 DP_mult_215_U1534 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_15_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_14_), .A(DP_mult_215_n1883), .ZN(
        DP_mult_215_n1882) );
  XNOR2_X1 DP_mult_215_U1533 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1882), 
        .ZN(DP_mult_215_n811) );
  OAI22_X1 DP_mult_215_U1532 ( .A1(DP_mult_215_n1700), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1701), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1881)
         );
  AOI221_X1 DP_mult_215_U1531 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_14_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_13_), .A(DP_mult_215_n1881), .ZN(
        DP_mult_215_n1880) );
  XNOR2_X1 DP_mult_215_U1530 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1880), 
        .ZN(DP_mult_215_n812) );
  OAI22_X1 DP_mult_215_U1529 ( .A1(DP_mult_215_n1696), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1697), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1879)
         );
  AOI221_X1 DP_mult_215_U1528 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_13_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_12_), .A(DP_mult_215_n1879), .ZN(
        DP_mult_215_n1878) );
  XNOR2_X1 DP_mult_215_U1527 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1878), 
        .ZN(DP_mult_215_n813) );
  OAI22_X1 DP_mult_215_U1526 ( .A1(DP_mult_215_n1692), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1693), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1877)
         );
  AOI221_X1 DP_mult_215_U1525 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_12_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_11_), .A(DP_mult_215_n1877), .ZN(
        DP_mult_215_n1876) );
  XNOR2_X1 DP_mult_215_U1524 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1876), 
        .ZN(DP_mult_215_n814) );
  OAI22_X1 DP_mult_215_U1523 ( .A1(DP_mult_215_n1688), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1689), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1875)
         );
  AOI221_X1 DP_mult_215_U1522 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_11_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_10_), .A(DP_mult_215_n1875), .ZN(
        DP_mult_215_n1874) );
  XNOR2_X1 DP_mult_215_U1521 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1874), 
        .ZN(DP_mult_215_n815) );
  OAI22_X1 DP_mult_215_U1520 ( .A1(DP_mult_215_n1684), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1685), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1873)
         );
  AOI221_X1 DP_mult_215_U1519 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_10_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_9_), .A(DP_mult_215_n1873), .ZN(
        DP_mult_215_n1872) );
  XNOR2_X1 DP_mult_215_U1518 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1872), 
        .ZN(DP_mult_215_n816) );
  OAI22_X1 DP_mult_215_U1517 ( .A1(DP_mult_215_n1680), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1681), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1871)
         );
  AOI221_X1 DP_mult_215_U1516 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_9_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_8_), .A(DP_mult_215_n1871), .ZN(
        DP_mult_215_n1870) );
  XNOR2_X1 DP_mult_215_U1515 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1870), 
        .ZN(DP_mult_215_n817) );
  OAI22_X1 DP_mult_215_U1514 ( .A1(DP_mult_215_n1676), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1677), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1869)
         );
  AOI221_X1 DP_mult_215_U1513 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_8_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_7_), .A(DP_mult_215_n1869), .ZN(
        DP_mult_215_n1868) );
  XNOR2_X1 DP_mult_215_U1512 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1868), 
        .ZN(DP_mult_215_n818) );
  OAI22_X1 DP_mult_215_U1511 ( .A1(DP_mult_215_n1672), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1673), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1867)
         );
  AOI221_X1 DP_mult_215_U1510 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_7_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_6_), .A(DP_mult_215_n1867), .ZN(
        DP_mult_215_n1866) );
  XNOR2_X1 DP_mult_215_U1509 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1866), 
        .ZN(DP_mult_215_n819) );
  OAI22_X1 DP_mult_215_U1508 ( .A1(DP_mult_215_n1668), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1669), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1865)
         );
  AOI221_X1 DP_mult_215_U1507 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_6_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_5_), .A(DP_mult_215_n1865), .ZN(
        DP_mult_215_n1864) );
  XNOR2_X1 DP_mult_215_U1506 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1864), 
        .ZN(DP_mult_215_n820) );
  OAI22_X1 DP_mult_215_U1505 ( .A1(DP_mult_215_n1664), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1665), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1863)
         );
  AOI221_X1 DP_mult_215_U1504 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_5_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_4_), .A(DP_mult_215_n1863), .ZN(
        DP_mult_215_n1862) );
  XNOR2_X1 DP_mult_215_U1503 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1862), 
        .ZN(DP_mult_215_n821) );
  OAI22_X1 DP_mult_215_U1502 ( .A1(DP_mult_215_n1660), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1661), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1861)
         );
  AOI221_X1 DP_mult_215_U1501 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_4_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_3_), .A(DP_mult_215_n1861), .ZN(
        DP_mult_215_n1860) );
  XNOR2_X1 DP_mult_215_U1500 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1860), 
        .ZN(DP_mult_215_n822) );
  OAI22_X1 DP_mult_215_U1499 ( .A1(DP_mult_215_n1657), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1649), .B2(DP_mult_215_n1587), .ZN(DP_mult_215_n1859)
         );
  AOI221_X1 DP_mult_215_U1498 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_3_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_2_), .A(DP_mult_215_n1859), .ZN(
        DP_mult_215_n1858) );
  XNOR2_X1 DP_mult_215_U1497 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1858), 
        .ZN(DP_mult_215_n823) );
  OAI22_X1 DP_mult_215_U1496 ( .A1(DP_mult_215_n1653), .A2(DP_mult_215_n1583), 
        .B1(DP_mult_215_n1565), .B2(DP_mult_215_n1586), .ZN(DP_mult_215_n1856)
         );
  AOI221_X1 DP_mult_215_U1495 ( .B1(DP_mult_215_n1584), .B2(DP_sw1_2_), .C1(
        DP_mult_215_n1585), .C2(DP_sw1_1_), .A(DP_mult_215_n1856), .ZN(
        DP_mult_215_n1855) );
  XNOR2_X1 DP_mult_215_U1494 ( .A(DP_mult_215_n1604), .B(DP_mult_215_n1855), 
        .ZN(DP_mult_215_n824) );
  OAI222_X1 DP_mult_215_U1493 ( .A1(DP_mult_215_n1649), .A2(DP_mult_215_n1533), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1539), .C1(DP_mult_215_n1650), 
        .C2(DP_mult_215_n1583), .ZN(DP_mult_215_n1854) );
  XNOR2_X1 DP_mult_215_U1492 ( .A(DP_mult_215_n1854), .B(DP_mult_215_n1605), 
        .ZN(DP_mult_215_n825) );
  OAI22_X1 DP_mult_215_U1491 ( .A1(DP_mult_215_n1565), .A2(DP_mult_215_n1533), 
        .B1(DP_mult_215_n1565), .B2(DP_mult_215_n1583), .ZN(DP_mult_215_n1853)
         );
  XNOR2_X1 DP_mult_215_U1490 ( .A(DP_mult_215_n1853), .B(DP_mult_215_n1605), 
        .ZN(DP_mult_215_n826) );
  XOR2_X1 DP_mult_215_U1489 ( .A(DP_coeff_ret1[9]), .B(DP_mult_215_n1601), .Z(
        DP_mult_215_n1852) );
  XNOR2_X1 DP_mult_215_U1488 ( .A(DP_coeff_ret1[10]), .B(DP_mult_215_n1603), 
        .ZN(DP_mult_215_n1851) );
  XNOR2_X1 DP_mult_215_U1487 ( .A(DP_coeff_ret1[10]), .B(DP_coeff_ret1[9]), 
        .ZN(DP_mult_215_n1850) );
  NAND3_X1 DP_mult_215_U1486 ( .A1(DP_mult_215_n1852), .A2(DP_mult_215_n1851), 
        .A3(DP_mult_215_n1850), .ZN(DP_mult_215_n1802) );
  INV_X1 DP_mult_215_U1485 ( .A(DP_mult_215_n1852), .ZN(DP_mult_215_n1849) );
  OAI21_X1 DP_mult_215_U1484 ( .B1(DP_mult_215_n1579), .B2(DP_mult_215_n1580), 
        .A(DP_mult_215_n1615), .ZN(DP_mult_215_n1848) );
  OAI221_X1 DP_mult_215_U1483 ( .B1(DP_mult_215_n1617), .B2(DP_mult_215_n1582), 
        .C1(DP_mult_215_n1620), .C2(DP_mult_215_n1578), .A(DP_mult_215_n1848), 
        .ZN(DP_mult_215_n1847) );
  XNOR2_X1 DP_mult_215_U1482 ( .A(DP_coeff_ret1[11]), .B(DP_mult_215_n1847), 
        .ZN(DP_mult_215_n827) );
  OAI22_X1 DP_mult_215_U1481 ( .A1(DP_mult_215_n1633), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1634), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1846)
         );
  AOI221_X1 DP_mult_215_U1480 ( .B1(DP_mult_215_n1579), .B2(DP_mult_215_n1615), 
        .C1(DP_mult_215_n1580), .C2(DP_mult_215_n1615), .A(DP_mult_215_n1846), 
        .ZN(DP_mult_215_n1845) );
  XNOR2_X1 DP_mult_215_U1479 ( .A(DP_coeff_ret1[11]), .B(DP_mult_215_n1845), 
        .ZN(DP_mult_215_n828) );
  OAI22_X1 DP_mult_215_U1478 ( .A1(DP_mult_215_n1617), .A2(DP_mult_215_n1545), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1844)
         );
  AOI221_X1 DP_mult_215_U1477 ( .B1(DP_mult_215_n1580), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1535), .C2(DP_mult_215_n1375), .A(DP_mult_215_n1844), 
        .ZN(DP_mult_215_n1843) );
  XNOR2_X1 DP_mult_215_U1476 ( .A(DP_coeff_ret1[11]), .B(DP_mult_215_n1843), 
        .ZN(DP_mult_215_n829) );
  OAI22_X1 DP_mult_215_U1475 ( .A1(DP_mult_215_n1640), .A2(DP_mult_215_n1582), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1538), .ZN(DP_mult_215_n1842)
         );
  AOI221_X1 DP_mult_215_U1474 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1535), .C2(DP_mult_215_n1376), .A(DP_mult_215_n1842), 
        .ZN(DP_mult_215_n1841) );
  XNOR2_X1 DP_mult_215_U1473 ( .A(DP_coeff_ret1[11]), .B(DP_mult_215_n1841), 
        .ZN(DP_mult_215_n830) );
  OAI22_X1 DP_mult_215_U1472 ( .A1(DP_mult_215_n1728), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1729), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1840)
         );
  AOI221_X1 DP_mult_215_U1471 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_21_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_20_), .A(DP_mult_215_n1840), .ZN(
        DP_mult_215_n1839) );
  XNOR2_X1 DP_mult_215_U1470 ( .A(DP_coeff_ret1[11]), .B(DP_mult_215_n1839), 
        .ZN(DP_mult_215_n831) );
  OAI22_X1 DP_mult_215_U1469 ( .A1(DP_mult_215_n1724), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1725), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1838)
         );
  AOI221_X1 DP_mult_215_U1468 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_20_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_19_), .A(DP_mult_215_n1838), .ZN(
        DP_mult_215_n1837) );
  XNOR2_X1 DP_mult_215_U1467 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1837), 
        .ZN(DP_mult_215_n832) );
  OAI22_X1 DP_mult_215_U1466 ( .A1(DP_mult_215_n1720), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1721), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1836)
         );
  AOI221_X1 DP_mult_215_U1465 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_19_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_18_), .A(DP_mult_215_n1836), .ZN(
        DP_mult_215_n1835) );
  XNOR2_X1 DP_mult_215_U1464 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1835), 
        .ZN(DP_mult_215_n833) );
  OAI22_X1 DP_mult_215_U1463 ( .A1(DP_mult_215_n1716), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1717), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1834)
         );
  AOI221_X1 DP_mult_215_U1462 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_18_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_17_), .A(DP_mult_215_n1834), .ZN(
        DP_mult_215_n1833) );
  XNOR2_X1 DP_mult_215_U1461 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1833), 
        .ZN(DP_mult_215_n834) );
  OAI22_X1 DP_mult_215_U1460 ( .A1(DP_mult_215_n1712), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1713), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1832)
         );
  AOI221_X1 DP_mult_215_U1459 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_17_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_16_), .A(DP_mult_215_n1832), .ZN(
        DP_mult_215_n1831) );
  XNOR2_X1 DP_mult_215_U1458 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1831), 
        .ZN(DP_mult_215_n835) );
  OAI22_X1 DP_mult_215_U1457 ( .A1(DP_mult_215_n1708), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1709), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1830)
         );
  AOI221_X1 DP_mult_215_U1456 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_16_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_15_), .A(DP_mult_215_n1830), .ZN(
        DP_mult_215_n1829) );
  XNOR2_X1 DP_mult_215_U1455 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1829), 
        .ZN(DP_mult_215_n836) );
  OAI22_X1 DP_mult_215_U1454 ( .A1(DP_mult_215_n1704), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1705), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1828)
         );
  AOI221_X1 DP_mult_215_U1453 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_15_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_14_), .A(DP_mult_215_n1828), .ZN(
        DP_mult_215_n1827) );
  XNOR2_X1 DP_mult_215_U1452 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1827), 
        .ZN(DP_mult_215_n837) );
  OAI22_X1 DP_mult_215_U1451 ( .A1(DP_mult_215_n1700), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1701), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1826)
         );
  AOI221_X1 DP_mult_215_U1450 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_14_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_13_), .A(DP_mult_215_n1826), .ZN(
        DP_mult_215_n1825) );
  XNOR2_X1 DP_mult_215_U1449 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1825), 
        .ZN(DP_mult_215_n838) );
  OAI22_X1 DP_mult_215_U1448 ( .A1(DP_mult_215_n1696), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1697), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1824)
         );
  AOI221_X1 DP_mult_215_U1447 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_13_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_12_), .A(DP_mult_215_n1824), .ZN(
        DP_mult_215_n1823) );
  XNOR2_X1 DP_mult_215_U1446 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1823), 
        .ZN(DP_mult_215_n839) );
  OAI22_X1 DP_mult_215_U1445 ( .A1(DP_mult_215_n1692), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1693), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1822)
         );
  AOI221_X1 DP_mult_215_U1444 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_12_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_11_), .A(DP_mult_215_n1822), .ZN(
        DP_mult_215_n1821) );
  XNOR2_X1 DP_mult_215_U1443 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1821), 
        .ZN(DP_mult_215_n840) );
  OAI22_X1 DP_mult_215_U1442 ( .A1(DP_mult_215_n1688), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1689), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1820)
         );
  AOI221_X1 DP_mult_215_U1441 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_11_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_10_), .A(DP_mult_215_n1820), .ZN(
        DP_mult_215_n1819) );
  XNOR2_X1 DP_mult_215_U1440 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1819), 
        .ZN(DP_mult_215_n841) );
  OAI22_X1 DP_mult_215_U1439 ( .A1(DP_mult_215_n1684), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1685), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1818)
         );
  AOI221_X1 DP_mult_215_U1438 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_10_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_9_), .A(DP_mult_215_n1818), .ZN(
        DP_mult_215_n1817) );
  XNOR2_X1 DP_mult_215_U1437 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1817), 
        .ZN(DP_mult_215_n842) );
  OAI22_X1 DP_mult_215_U1436 ( .A1(DP_mult_215_n1680), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1681), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1816)
         );
  AOI221_X1 DP_mult_215_U1435 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_9_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_8_), .A(DP_mult_215_n1816), .ZN(
        DP_mult_215_n1815) );
  XNOR2_X1 DP_mult_215_U1434 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1815), 
        .ZN(DP_mult_215_n843) );
  OAI22_X1 DP_mult_215_U1433 ( .A1(DP_mult_215_n1676), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1677), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1814)
         );
  AOI221_X1 DP_mult_215_U1432 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_8_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_7_), .A(DP_mult_215_n1814), .ZN(
        DP_mult_215_n1813) );
  XNOR2_X1 DP_mult_215_U1431 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1813), 
        .ZN(DP_mult_215_n844) );
  OAI22_X1 DP_mult_215_U1430 ( .A1(DP_mult_215_n1672), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1673), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1812)
         );
  AOI221_X1 DP_mult_215_U1429 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_7_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_6_), .A(DP_mult_215_n1812), .ZN(
        DP_mult_215_n1811) );
  XNOR2_X1 DP_mult_215_U1428 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1811), 
        .ZN(DP_mult_215_n845) );
  OAI22_X1 DP_mult_215_U1427 ( .A1(DP_mult_215_n1668), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1669), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1810)
         );
  AOI221_X1 DP_mult_215_U1426 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_6_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_5_), .A(DP_mult_215_n1810), .ZN(
        DP_mult_215_n1809) );
  XNOR2_X1 DP_mult_215_U1425 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1809), 
        .ZN(DP_mult_215_n846) );
  OAI22_X1 DP_mult_215_U1424 ( .A1(DP_mult_215_n1664), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1665), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1808)
         );
  AOI221_X1 DP_mult_215_U1423 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_5_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_4_), .A(DP_mult_215_n1808), .ZN(
        DP_mult_215_n1807) );
  XNOR2_X1 DP_mult_215_U1422 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1807), 
        .ZN(DP_mult_215_n847) );
  OAI22_X1 DP_mult_215_U1421 ( .A1(DP_mult_215_n1660), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1661), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1806)
         );
  AOI221_X1 DP_mult_215_U1420 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_4_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_3_), .A(DP_mult_215_n1806), .ZN(
        DP_mult_215_n1805) );
  XNOR2_X1 DP_mult_215_U1419 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1805), 
        .ZN(DP_mult_215_n848) );
  OAI22_X1 DP_mult_215_U1418 ( .A1(DP_mult_215_n1657), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1649), .B2(DP_mult_215_n1582), .ZN(DP_mult_215_n1804)
         );
  AOI221_X1 DP_mult_215_U1417 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_3_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_2_), .A(DP_mult_215_n1804), .ZN(
        DP_mult_215_n1803) );
  XNOR2_X1 DP_mult_215_U1416 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1803), 
        .ZN(DP_mult_215_n849) );
  OAI22_X1 DP_mult_215_U1415 ( .A1(DP_mult_215_n1653), .A2(DP_mult_215_n1578), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1581), .ZN(DP_mult_215_n1801)
         );
  AOI221_X1 DP_mult_215_U1414 ( .B1(DP_mult_215_n1579), .B2(DP_sw1_2_), .C1(
        DP_mult_215_n1580), .C2(DP_sw1_1_), .A(DP_mult_215_n1801), .ZN(
        DP_mult_215_n1800) );
  XNOR2_X1 DP_mult_215_U1413 ( .A(DP_mult_215_n1602), .B(DP_mult_215_n1800), 
        .ZN(DP_mult_215_n850) );
  OAI222_X1 DP_mult_215_U1412 ( .A1(DP_mult_215_n1649), .A2(DP_mult_215_n1545), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1538), .C1(DP_mult_215_n1650), 
        .C2(DP_mult_215_n1578), .ZN(DP_mult_215_n1799) );
  XNOR2_X1 DP_mult_215_U1411 ( .A(DP_mult_215_n1799), .B(DP_mult_215_n1603), 
        .ZN(DP_mult_215_n851) );
  OAI22_X1 DP_mult_215_U1410 ( .A1(DP_mult_215_n1565), .A2(DP_mult_215_n1545), 
        .B1(DP_mult_215_n1565), .B2(DP_mult_215_n1578), .ZN(DP_mult_215_n1798)
         );
  XNOR2_X1 DP_mult_215_U1409 ( .A(DP_mult_215_n1798), .B(DP_mult_215_n1603), 
        .ZN(DP_mult_215_n852) );
  XOR2_X1 DP_mult_215_U1408 ( .A(DP_coeff_ret1[6]), .B(DP_mult_215_n1599), .Z(
        DP_mult_215_n1797) );
  XNOR2_X1 DP_mult_215_U1407 ( .A(DP_coeff_ret1[7]), .B(DP_mult_215_n1601), 
        .ZN(DP_mult_215_n1796) );
  XNOR2_X1 DP_mult_215_U1406 ( .A(DP_coeff_ret1[6]), .B(DP_coeff_ret1[7]), 
        .ZN(DP_mult_215_n1795) );
  NAND3_X1 DP_mult_215_U1405 ( .A1(DP_mult_215_n1797), .A2(DP_mult_215_n1796), 
        .A3(DP_mult_215_n1795), .ZN(DP_mult_215_n1747) );
  INV_X1 DP_mult_215_U1404 ( .A(DP_mult_215_n1797), .ZN(DP_mult_215_n1794) );
  OAI21_X1 DP_mult_215_U1403 ( .B1(DP_mult_215_n1574), .B2(DP_mult_215_n1575), 
        .A(DP_mult_215_n1615), .ZN(DP_mult_215_n1793) );
  OAI221_X1 DP_mult_215_U1402 ( .B1(DP_mult_215_n1617), .B2(DP_mult_215_n1577), 
        .C1(DP_mult_215_n1620), .C2(DP_mult_215_n1573), .A(DP_mult_215_n1793), 
        .ZN(DP_mult_215_n1792) );
  XNOR2_X1 DP_mult_215_U1401 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1792), 
        .ZN(DP_mult_215_n853) );
  OAI22_X1 DP_mult_215_U1400 ( .A1(DP_mult_215_n1633), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1634), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1791)
         );
  AOI221_X1 DP_mult_215_U1399 ( .B1(DP_mult_215_n1574), .B2(DP_mult_215_n1614), 
        .C1(DP_mult_215_n1575), .C2(DP_mult_215_n1615), .A(DP_mult_215_n1791), 
        .ZN(DP_mult_215_n1790) );
  XNOR2_X1 DP_mult_215_U1398 ( .A(DP_coeff_ret1[8]), .B(DP_mult_215_n1790), 
        .ZN(DP_mult_215_n854) );
  OAI22_X1 DP_mult_215_U1397 ( .A1(DP_mult_215_n1617), .A2(DP_mult_215_n1544), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1789)
         );
  AOI221_X1 DP_mult_215_U1396 ( .B1(DP_mult_215_n1575), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1546), .C2(DP_mult_215_n1375), .A(DP_mult_215_n1789), 
        .ZN(DP_mult_215_n1788) );
  XNOR2_X1 DP_mult_215_U1395 ( .A(DP_coeff_ret1[8]), .B(DP_mult_215_n1788), 
        .ZN(DP_mult_215_n855) );
  OAI22_X1 DP_mult_215_U1394 ( .A1(DP_mult_215_n1640), .A2(DP_mult_215_n1577), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1547), .ZN(DP_mult_215_n1787)
         );
  AOI221_X1 DP_mult_215_U1393 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1546), .C2(DP_mult_215_n1376), .A(DP_mult_215_n1787), 
        .ZN(DP_mult_215_n1786) );
  XNOR2_X1 DP_mult_215_U1392 ( .A(DP_coeff_ret1[8]), .B(DP_mult_215_n1786), 
        .ZN(DP_mult_215_n856) );
  OAI22_X1 DP_mult_215_U1391 ( .A1(DP_mult_215_n1728), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1729), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1785)
         );
  AOI221_X1 DP_mult_215_U1390 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_21_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_20_), .A(DP_mult_215_n1785), .ZN(
        DP_mult_215_n1784) );
  XNOR2_X1 DP_mult_215_U1389 ( .A(DP_coeff_ret1[8]), .B(DP_mult_215_n1784), 
        .ZN(DP_mult_215_n857) );
  OAI22_X1 DP_mult_215_U1388 ( .A1(DP_mult_215_n1724), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1725), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1783)
         );
  AOI221_X1 DP_mult_215_U1387 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_20_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_19_), .A(DP_mult_215_n1783), .ZN(
        DP_mult_215_n1782) );
  XNOR2_X1 DP_mult_215_U1386 ( .A(DP_coeff_ret1[8]), .B(DP_mult_215_n1782), 
        .ZN(DP_mult_215_n858) );
  OAI22_X1 DP_mult_215_U1385 ( .A1(DP_mult_215_n1720), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1721), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1781)
         );
  AOI221_X1 DP_mult_215_U1384 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_19_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_18_), .A(DP_mult_215_n1781), .ZN(
        DP_mult_215_n1780) );
  XNOR2_X1 DP_mult_215_U1383 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1780), 
        .ZN(DP_mult_215_n859) );
  OAI22_X1 DP_mult_215_U1382 ( .A1(DP_mult_215_n1716), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1717), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1779)
         );
  AOI221_X1 DP_mult_215_U1381 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_18_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_17_), .A(DP_mult_215_n1779), .ZN(
        DP_mult_215_n1778) );
  XNOR2_X1 DP_mult_215_U1380 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1778), 
        .ZN(DP_mult_215_n860) );
  OAI22_X1 DP_mult_215_U1379 ( .A1(DP_mult_215_n1712), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1713), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1777)
         );
  AOI221_X1 DP_mult_215_U1378 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_17_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_16_), .A(DP_mult_215_n1777), .ZN(
        DP_mult_215_n1776) );
  XNOR2_X1 DP_mult_215_U1377 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1776), 
        .ZN(DP_mult_215_n861) );
  OAI22_X1 DP_mult_215_U1376 ( .A1(DP_mult_215_n1708), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1709), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1775)
         );
  AOI221_X1 DP_mult_215_U1375 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_16_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_15_), .A(DP_mult_215_n1775), .ZN(
        DP_mult_215_n1774) );
  XNOR2_X1 DP_mult_215_U1374 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1774), 
        .ZN(DP_mult_215_n862) );
  OAI22_X1 DP_mult_215_U1373 ( .A1(DP_mult_215_n1704), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1705), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1773)
         );
  AOI221_X1 DP_mult_215_U1372 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_15_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_14_), .A(DP_mult_215_n1773), .ZN(
        DP_mult_215_n1772) );
  XNOR2_X1 DP_mult_215_U1371 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1772), 
        .ZN(DP_mult_215_n863) );
  OAI22_X1 DP_mult_215_U1370 ( .A1(DP_mult_215_n1700), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1701), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1771)
         );
  AOI221_X1 DP_mult_215_U1369 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_14_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_13_), .A(DP_mult_215_n1771), .ZN(
        DP_mult_215_n1770) );
  XNOR2_X1 DP_mult_215_U1368 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1770), 
        .ZN(DP_mult_215_n864) );
  OAI22_X1 DP_mult_215_U1367 ( .A1(DP_mult_215_n1696), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1697), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1769)
         );
  AOI221_X1 DP_mult_215_U1366 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_13_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_12_), .A(DP_mult_215_n1769), .ZN(
        DP_mult_215_n1768) );
  XNOR2_X1 DP_mult_215_U1365 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1768), 
        .ZN(DP_mult_215_n865) );
  OAI22_X1 DP_mult_215_U1364 ( .A1(DP_mult_215_n1692), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1693), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1767)
         );
  AOI221_X1 DP_mult_215_U1363 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_12_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_11_), .A(DP_mult_215_n1767), .ZN(
        DP_mult_215_n1766) );
  XNOR2_X1 DP_mult_215_U1362 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1766), 
        .ZN(DP_mult_215_n866) );
  OAI22_X1 DP_mult_215_U1361 ( .A1(DP_mult_215_n1688), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1689), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1765)
         );
  AOI221_X1 DP_mult_215_U1360 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_11_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_10_), .A(DP_mult_215_n1765), .ZN(
        DP_mult_215_n1764) );
  XNOR2_X1 DP_mult_215_U1359 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1764), 
        .ZN(DP_mult_215_n867) );
  OAI22_X1 DP_mult_215_U1358 ( .A1(DP_mult_215_n1684), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1685), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1763)
         );
  AOI221_X1 DP_mult_215_U1357 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_10_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_9_), .A(DP_mult_215_n1763), .ZN(
        DP_mult_215_n1762) );
  XNOR2_X1 DP_mult_215_U1356 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1762), 
        .ZN(DP_mult_215_n868) );
  OAI22_X1 DP_mult_215_U1355 ( .A1(DP_mult_215_n1680), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1681), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1761)
         );
  AOI221_X1 DP_mult_215_U1354 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_9_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_8_), .A(DP_mult_215_n1761), .ZN(
        DP_mult_215_n1760) );
  XNOR2_X1 DP_mult_215_U1353 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1760), 
        .ZN(DP_mult_215_n869) );
  OAI22_X1 DP_mult_215_U1352 ( .A1(DP_mult_215_n1676), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1677), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1759)
         );
  AOI221_X1 DP_mult_215_U1351 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_8_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_7_), .A(DP_mult_215_n1759), .ZN(
        DP_mult_215_n1758) );
  XNOR2_X1 DP_mult_215_U1350 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1758), 
        .ZN(DP_mult_215_n870) );
  OAI22_X1 DP_mult_215_U1349 ( .A1(DP_mult_215_n1672), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1673), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1757)
         );
  AOI221_X1 DP_mult_215_U1348 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_7_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_6_), .A(DP_mult_215_n1757), .ZN(
        DP_mult_215_n1756) );
  XNOR2_X1 DP_mult_215_U1347 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1756), 
        .ZN(DP_mult_215_n871) );
  OAI22_X1 DP_mult_215_U1346 ( .A1(DP_mult_215_n1668), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1669), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1755)
         );
  AOI221_X1 DP_mult_215_U1345 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_6_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_5_), .A(DP_mult_215_n1755), .ZN(
        DP_mult_215_n1754) );
  XNOR2_X1 DP_mult_215_U1344 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1754), 
        .ZN(DP_mult_215_n872) );
  OAI22_X1 DP_mult_215_U1343 ( .A1(DP_mult_215_n1664), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1665), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1753)
         );
  AOI221_X1 DP_mult_215_U1342 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_5_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_4_), .A(DP_mult_215_n1753), .ZN(
        DP_mult_215_n1752) );
  XNOR2_X1 DP_mult_215_U1341 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1752), 
        .ZN(DP_mult_215_n873) );
  OAI22_X1 DP_mult_215_U1340 ( .A1(DP_mult_215_n1660), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1661), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1751)
         );
  AOI221_X1 DP_mult_215_U1339 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_4_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_3_), .A(DP_mult_215_n1751), .ZN(
        DP_mult_215_n1750) );
  XNOR2_X1 DP_mult_215_U1338 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1750), 
        .ZN(DP_mult_215_n874) );
  OAI22_X1 DP_mult_215_U1337 ( .A1(DP_mult_215_n1657), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1649), .B2(DP_mult_215_n1577), .ZN(DP_mult_215_n1749)
         );
  AOI221_X1 DP_mult_215_U1336 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_3_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_2_), .A(DP_mult_215_n1749), .ZN(
        DP_mult_215_n1748) );
  XNOR2_X1 DP_mult_215_U1335 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1748), 
        .ZN(DP_mult_215_n875) );
  OAI22_X1 DP_mult_215_U1334 ( .A1(DP_mult_215_n1653), .A2(DP_mult_215_n1573), 
        .B1(DP_mult_215_n1565), .B2(DP_mult_215_n1576), .ZN(DP_mult_215_n1746)
         );
  AOI221_X1 DP_mult_215_U1333 ( .B1(DP_mult_215_n1574), .B2(DP_sw1_2_), .C1(
        DP_mult_215_n1575), .C2(DP_sw1_1_), .A(DP_mult_215_n1746), .ZN(
        DP_mult_215_n1745) );
  XNOR2_X1 DP_mult_215_U1332 ( .A(DP_mult_215_n1600), .B(DP_mult_215_n1745), 
        .ZN(DP_mult_215_n876) );
  OAI222_X1 DP_mult_215_U1331 ( .A1(DP_mult_215_n1649), .A2(DP_mult_215_n1544), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1547), .C1(DP_mult_215_n1650), 
        .C2(DP_mult_215_n1573), .ZN(DP_mult_215_n1744) );
  XNOR2_X1 DP_mult_215_U1330 ( .A(DP_mult_215_n1744), .B(DP_mult_215_n1601), 
        .ZN(DP_mult_215_n877) );
  OAI22_X1 DP_mult_215_U1329 ( .A1(DP_mult_215_n1565), .A2(DP_mult_215_n1544), 
        .B1(DP_mult_215_n1565), .B2(DP_mult_215_n1573), .ZN(DP_mult_215_n1743)
         );
  XNOR2_X1 DP_mult_215_U1328 ( .A(DP_mult_215_n1743), .B(DP_mult_215_n1601), 
        .ZN(DP_mult_215_n878) );
  XOR2_X1 DP_mult_215_U1327 ( .A(DP_coeff_ret1[3]), .B(DP_mult_215_n1742), .Z(
        DP_mult_215_n1741) );
  XNOR2_X1 DP_mult_215_U1326 ( .A(DP_coeff_ret1[4]), .B(DP_mult_215_n1599), 
        .ZN(DP_mult_215_n1740) );
  XNOR2_X1 DP_mult_215_U1325 ( .A(DP_coeff_ret1[3]), .B(DP_coeff_ret1[4]), 
        .ZN(DP_mult_215_n1739) );
  NAND3_X1 DP_mult_215_U1324 ( .A1(DP_mult_215_n1741), .A2(DP_mult_215_n1740), 
        .A3(DP_mult_215_n1739), .ZN(DP_mult_215_n1654) );
  INV_X1 DP_mult_215_U1323 ( .A(DP_mult_215_n1741), .ZN(DP_mult_215_n1738) );
  OAI21_X1 DP_mult_215_U1322 ( .B1(DP_mult_215_n1569), .B2(DP_mult_215_n1570), 
        .A(DP_mult_215_n1615), .ZN(DP_mult_215_n1737) );
  OAI221_X1 DP_mult_215_U1321 ( .B1(DP_mult_215_n1617), .B2(DP_mult_215_n1572), 
        .C1(DP_mult_215_n1620), .C2(DP_mult_215_n1568), .A(DP_mult_215_n1737), 
        .ZN(DP_mult_215_n1736) );
  XNOR2_X1 DP_mult_215_U1320 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1736), 
        .ZN(DP_mult_215_n879) );
  OAI22_X1 DP_mult_215_U1319 ( .A1(DP_mult_215_n1633), .A2(DP_mult_215_n1568), 
        .B1(DP_mult_215_n1634), .B2(DP_mult_215_n1572), .ZN(DP_mult_215_n1735)
         );
  AOI221_X1 DP_mult_215_U1318 ( .B1(DP_mult_215_n1569), .B2(DP_mult_215_n1614), 
        .C1(DP_mult_215_n1570), .C2(DP_mult_215_n1615), .A(DP_mult_215_n1735), 
        .ZN(DP_mult_215_n1734) );
  XNOR2_X1 DP_mult_215_U1317 ( .A(DP_coeff_ret1[5]), .B(DP_mult_215_n1734), 
        .ZN(DP_mult_215_n880) );
  OAI22_X1 DP_mult_215_U1316 ( .A1(DP_mult_215_n1616), .A2(DP_mult_215_n1552), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1572), .ZN(DP_mult_215_n1733)
         );
  AOI221_X1 DP_mult_215_U1315 ( .B1(DP_mult_215_n1570), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1551), .C2(DP_mult_215_n1375), .A(DP_mult_215_n1733), 
        .ZN(DP_mult_215_n1732) );
  XNOR2_X1 DP_mult_215_U1314 ( .A(DP_coeff_ret1[5]), .B(DP_mult_215_n1732), 
        .ZN(DP_mult_215_n881) );
  OAI22_X1 DP_mult_215_U1313 ( .A1(DP_mult_215_n1640), .A2(DP_mult_215_n1572), 
        .B1(DP_mult_215_n1643), .B2(DP_mult_215_n1553), .ZN(DP_mult_215_n1731)
         );
  AOI221_X1 DP_mult_215_U1312 ( .B1(DP_mult_215_n1569), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1551), .C2(DP_mult_215_n1376), .A(DP_mult_215_n1731), 
        .ZN(DP_mult_215_n1730) );
  XNOR2_X1 DP_mult_215_U1311 ( .A(DP_coeff_ret1[5]), .B(DP_mult_215_n1730), 
        .ZN(DP_mult_215_n882) );
  OAI22_X1 DP_mult_215_U1310 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1728), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1729), .ZN(DP_mult_215_n1727)
         );
  AOI221_X1 DP_mult_215_U1309 ( .B1(DP_mult_215_n1569), .B2(DP_sw1_21_), .C1(
        DP_mult_215_n1570), .C2(DP_sw1_20_), .A(DP_mult_215_n1727), .ZN(
        DP_mult_215_n1726) );
  XNOR2_X1 DP_mult_215_U1308 ( .A(DP_coeff_ret1[5]), .B(DP_mult_215_n1726), 
        .ZN(DP_mult_215_n883) );
  OAI22_X1 DP_mult_215_U1307 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1724), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1725), .ZN(DP_mult_215_n1723)
         );
  AOI221_X1 DP_mult_215_U1306 ( .B1(DP_mult_215_n1569), .B2(DP_sw1_20_), .C1(
        DP_sw1_19_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1723), .ZN(
        DP_mult_215_n1722) );
  XNOR2_X1 DP_mult_215_U1305 ( .A(DP_coeff_ret1[5]), .B(DP_mult_215_n1722), 
        .ZN(DP_mult_215_n884) );
  OAI22_X1 DP_mult_215_U1304 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1720), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1721), .ZN(DP_mult_215_n1719)
         );
  AOI221_X1 DP_mult_215_U1303 ( .B1(DP_sw1_19_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_18_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1719), .ZN(
        DP_mult_215_n1718) );
  XNOR2_X1 DP_mult_215_U1302 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1718), 
        .ZN(DP_mult_215_n885) );
  OAI22_X1 DP_mult_215_U1301 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1716), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1717), .ZN(DP_mult_215_n1715)
         );
  AOI221_X1 DP_mult_215_U1300 ( .B1(DP_sw1_18_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_17_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1715), .ZN(
        DP_mult_215_n1714) );
  XNOR2_X1 DP_mult_215_U1299 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1714), 
        .ZN(DP_mult_215_n886) );
  OAI22_X1 DP_mult_215_U1298 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1712), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1713), .ZN(DP_mult_215_n1711)
         );
  AOI221_X1 DP_mult_215_U1297 ( .B1(DP_sw1_17_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_16_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1711), .ZN(
        DP_mult_215_n1710) );
  XNOR2_X1 DP_mult_215_U1296 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1710), 
        .ZN(DP_mult_215_n887) );
  OAI22_X1 DP_mult_215_U1295 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1708), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1709), .ZN(DP_mult_215_n1707)
         );
  AOI221_X1 DP_mult_215_U1294 ( .B1(DP_sw1_16_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_15_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1707), .ZN(
        DP_mult_215_n1706) );
  XNOR2_X1 DP_mult_215_U1293 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1706), 
        .ZN(DP_mult_215_n888) );
  OAI22_X1 DP_mult_215_U1292 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1704), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1705), .ZN(DP_mult_215_n1703)
         );
  AOI221_X1 DP_mult_215_U1291 ( .B1(DP_sw1_15_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_14_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1703), .ZN(
        DP_mult_215_n1702) );
  XNOR2_X1 DP_mult_215_U1290 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1702), 
        .ZN(DP_mult_215_n889) );
  OAI22_X1 DP_mult_215_U1289 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1700), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1701), .ZN(DP_mult_215_n1699)
         );
  AOI221_X1 DP_mult_215_U1288 ( .B1(DP_sw1_14_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_13_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1699), .ZN(
        DP_mult_215_n1698) );
  XNOR2_X1 DP_mult_215_U1287 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1698), 
        .ZN(DP_mult_215_n890) );
  OAI22_X1 DP_mult_215_U1286 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1696), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1697), .ZN(DP_mult_215_n1695)
         );
  AOI221_X1 DP_mult_215_U1285 ( .B1(DP_sw1_13_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_12_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1695), .ZN(
        DP_mult_215_n1694) );
  XNOR2_X1 DP_mult_215_U1284 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1694), 
        .ZN(DP_mult_215_n891) );
  OAI22_X1 DP_mult_215_U1283 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1692), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1693), .ZN(DP_mult_215_n1691)
         );
  AOI221_X1 DP_mult_215_U1282 ( .B1(DP_sw1_12_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_11_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1691), .ZN(
        DP_mult_215_n1690) );
  XNOR2_X1 DP_mult_215_U1281 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1690), 
        .ZN(DP_mult_215_n892) );
  OAI22_X1 DP_mult_215_U1280 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1688), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1689), .ZN(DP_mult_215_n1687)
         );
  AOI221_X1 DP_mult_215_U1279 ( .B1(DP_sw1_11_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_10_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1687), .ZN(
        DP_mult_215_n1686) );
  XNOR2_X1 DP_mult_215_U1278 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1686), 
        .ZN(DP_mult_215_n893) );
  OAI22_X1 DP_mult_215_U1277 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1684), 
        .B1(DP_mult_215_n1572), .B2(DP_mult_215_n1685), .ZN(DP_mult_215_n1683)
         );
  AOI221_X1 DP_mult_215_U1276 ( .B1(DP_sw1_10_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_9_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1683), .ZN(
        DP_mult_215_n1682) );
  XNOR2_X1 DP_mult_215_U1275 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1682), 
        .ZN(DP_mult_215_n894) );
  OAI22_X1 DP_mult_215_U1274 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1680), 
        .B1(DP_mult_215_n1572), .B2(DP_mult_215_n1681), .ZN(DP_mult_215_n1679)
         );
  AOI221_X1 DP_mult_215_U1273 ( .B1(DP_sw1_9_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_8_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1679), .ZN(
        DP_mult_215_n1678) );
  XNOR2_X1 DP_mult_215_U1272 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1678), 
        .ZN(DP_mult_215_n895) );
  OAI22_X1 DP_mult_215_U1271 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1676), 
        .B1(DP_mult_215_n1571), .B2(DP_mult_215_n1677), .ZN(DP_mult_215_n1675)
         );
  AOI221_X1 DP_mult_215_U1270 ( .B1(DP_sw1_8_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_7_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1675), .ZN(
        DP_mult_215_n1674) );
  XNOR2_X1 DP_mult_215_U1269 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1674), 
        .ZN(DP_mult_215_n896) );
  OAI22_X1 DP_mult_215_U1268 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1672), 
        .B1(DP_mult_215_n1572), .B2(DP_mult_215_n1673), .ZN(DP_mult_215_n1671)
         );
  AOI221_X1 DP_mult_215_U1267 ( .B1(DP_sw1_7_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_6_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1671), .ZN(
        DP_mult_215_n1670) );
  XNOR2_X1 DP_mult_215_U1266 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1670), 
        .ZN(DP_mult_215_n897) );
  OAI22_X1 DP_mult_215_U1265 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1668), 
        .B1(DP_mult_215_n1572), .B2(DP_mult_215_n1669), .ZN(DP_mult_215_n1667)
         );
  AOI221_X1 DP_mult_215_U1264 ( .B1(DP_sw1_6_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_5_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1667), .ZN(
        DP_mult_215_n1666) );
  XNOR2_X1 DP_mult_215_U1263 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1666), 
        .ZN(DP_mult_215_n898) );
  OAI22_X1 DP_mult_215_U1262 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1664), 
        .B1(DP_mult_215_n1572), .B2(DP_mult_215_n1665), .ZN(DP_mult_215_n1663)
         );
  AOI221_X1 DP_mult_215_U1261 ( .B1(DP_sw1_5_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_4_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1663), .ZN(
        DP_mult_215_n1662) );
  XNOR2_X1 DP_mult_215_U1260 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1662), 
        .ZN(DP_mult_215_n899) );
  OAI22_X1 DP_mult_215_U1259 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1660), 
        .B1(DP_mult_215_n1661), .B2(DP_mult_215_n1572), .ZN(DP_mult_215_n1659)
         );
  AOI221_X1 DP_mult_215_U1258 ( .B1(DP_sw1_4_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_3_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1659), .ZN(
        DP_mult_215_n1658) );
  XNOR2_X1 DP_mult_215_U1257 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1658), 
        .ZN(DP_mult_215_n900) );
  OAI22_X1 DP_mult_215_U1256 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1657), 
        .B1(DP_mult_215_n1649), .B2(DP_mult_215_n1572), .ZN(DP_mult_215_n1656)
         );
  AOI221_X1 DP_mult_215_U1255 ( .B1(DP_sw1_3_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_2_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1656), .ZN(
        DP_mult_215_n1655) );
  XNOR2_X1 DP_mult_215_U1254 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1655), 
        .ZN(DP_mult_215_n901) );
  OAI22_X1 DP_mult_215_U1253 ( .A1(DP_mult_215_n1568), .A2(DP_mult_215_n1653), 
        .B1(DP_mult_215_n1565), .B2(DP_mult_215_n1572), .ZN(DP_mult_215_n1652)
         );
  AOI221_X1 DP_mult_215_U1252 ( .B1(DP_sw1_2_), .B2(DP_mult_215_n1569), .C1(
        DP_sw1_1_), .C2(DP_mult_215_n1570), .A(DP_mult_215_n1652), .ZN(
        DP_mult_215_n1651) );
  XNOR2_X1 DP_mult_215_U1251 ( .A(DP_mult_215_n1598), .B(DP_mult_215_n1651), 
        .ZN(DP_mult_215_n902) );
  OAI222_X1 DP_mult_215_U1250 ( .A1(DP_mult_215_n1552), .A2(DP_mult_215_n1649), 
        .B1(DP_mult_215_n1566), .B2(DP_mult_215_n1553), .C1(DP_mult_215_n1568), 
        .C2(DP_mult_215_n1650), .ZN(DP_mult_215_n1648) );
  XNOR2_X1 DP_mult_215_U1249 ( .A(DP_mult_215_n1648), .B(DP_mult_215_n1599), 
        .ZN(DP_mult_215_n903) );
  OAI22_X1 DP_mult_215_U1248 ( .A1(DP_mult_215_n1565), .A2(DP_mult_215_n1552), 
        .B1(DP_mult_215_n1568), .B2(DP_mult_215_n1567), .ZN(DP_mult_215_n1646)
         );
  XNOR2_X1 DP_mult_215_U1247 ( .A(DP_mult_215_n1646), .B(DP_mult_215_n1599), 
        .ZN(DP_mult_215_n904) );
  OAI22_X1 DP_mult_215_U1246 ( .A1(DP_mult_215_n1633), .A2(DP_mult_215_n1564), 
        .B1(DP_mult_215_n1634), .B2(DP_mult_215_n1639), .ZN(DP_mult_215_n1645)
         );
  AOI221_X1 DP_mult_215_U1245 ( .B1(DP_mult_215_n1561), .B2(DP_mult_215_n1614), 
        .C1(DP_mult_215_n1563), .C2(DP_mult_215_n1615), .A(DP_mult_215_n1645), 
        .ZN(DP_mult_215_n1644) );
  XNOR2_X1 DP_mult_215_U1244 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n1644), 
        .ZN(DP_mult_215_n906) );
  OAI22_X1 DP_mult_215_U1243 ( .A1(DP_mult_215_n1643), .A2(DP_mult_215_n1639), 
        .B1(DP_mult_215_n1617), .B2(DP_mult_215_n1554), .ZN(DP_mult_215_n1642)
         );
  AOI221_X1 DP_mult_215_U1242 ( .B1(DP_mult_215_n1563), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1555), .C2(DP_mult_215_n1375), .A(DP_mult_215_n1642), 
        .ZN(DP_mult_215_n1641) );
  XNOR2_X1 DP_mult_215_U1241 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n1641), 
        .ZN(DP_mult_215_n907) );
  INV_X1 DP_mult_215_U1240 ( .A(DP_mult_215_n1376), .ZN(DP_mult_215_n1638) );
  OAI22_X1 DP_mult_215_U1239 ( .A1(DP_mult_215_n1564), .A2(DP_mult_215_n1638), 
        .B1(DP_mult_215_n1639), .B2(DP_mult_215_n1640), .ZN(DP_mult_215_n1637)
         );
  AOI221_X1 DP_mult_215_U1238 ( .B1(DP_mult_215_n1561), .B2(DP_sw1_22_), .C1(
        DP_mult_215_n1563), .C2(DP_sw1_21_), .A(DP_mult_215_n1637), .ZN(
        DP_mult_215_n1635) );
  XNOR2_X1 DP_mult_215_U1237 ( .A(DP_coeff_ret1[2]), .B(DP_mult_215_n1635), 
        .ZN(DP_mult_215_n908) );
  OAI22_X1 DP_mult_215_U1236 ( .A1(DP_mult_215_n1558), .A2(DP_mult_215_n1633), 
        .B1(DP_mult_215_n1557), .B2(DP_mult_215_n1634), .ZN(DP_mult_215_n1632)
         );
  AOI221_X1 DP_mult_215_U1235 ( .B1(DP_mult_215_n1613), .B2(DP_mult_215_n1559), 
        .C1(DP_mult_215_n1560), .C2(DP_mult_215_n1615), .A(DP_mult_215_n1632), 
        .ZN(DP_mult_215_n1631) );
  XOR2_X1 DP_mult_215_U1234 ( .A(DP_coeff_ret1[23]), .B(DP_mult_215_n1631), 
        .Z(DP_mult_215_n1625) );
  INV_X1 DP_mult_215_U1233 ( .A(DP_mult_215_n1625), .ZN(DP_mult_215_n1621) );
  OAI21_X1 DP_mult_215_U1232 ( .B1(DP_mult_215_n1559), .B2(DP_mult_215_n1560), 
        .A(DP_mult_215_n1615), .ZN(DP_mult_215_n1630) );
  OAI221_X1 DP_mult_215_U1231 ( .B1(DP_mult_215_n1617), .B2(DP_mult_215_n1557), 
        .C1(DP_mult_215_n1620), .C2(DP_mult_215_n1558), .A(DP_mult_215_n1630), 
        .ZN(DP_mult_215_n1628) );
  XOR2_X1 DP_mult_215_U1230 ( .A(DP_mult_215_n1628), .B(DP_mult_215_n1611), 
        .Z(DP_mult_215_n1622) );
  AOI222_X1 DP_mult_215_U1229 ( .A1(DP_mult_215_n1627), .A2(DP_mult_215_n303), 
        .B1(DP_mult_215_n1625), .B2(DP_mult_215_n303), .C1(DP_mult_215_n1627), 
        .C2(DP_mult_215_n1625), .ZN(DP_mult_215_n1624) );
  INV_X1 DP_mult_215_U1228 ( .A(DP_mult_215_n1622), .ZN(DP_mult_215_n1626) );
  OAI22_X1 DP_mult_215_U1227 ( .A1(DP_mult_215_n1624), .A2(DP_mult_215_n1625), 
        .B1(DP_mult_215_n1624), .B2(DP_mult_215_n1626), .ZN(DP_mult_215_n1623)
         );
  AOI21_X1 DP_mult_215_U1226 ( .B1(DP_mult_215_n1621), .B2(DP_mult_215_n1622), 
        .A(DP_mult_215_n1623), .ZN(DP_sw1_coeff_ret1[23]) );
  INV_X1 DP_mult_215_U1225 ( .A(DP_mult_215_n1614), .ZN(DP_mult_215_n1620) );
  INV_X1 DP_mult_215_U1224 ( .A(DP_mult_215_n1614), .ZN(DP_mult_215_n1619) );
  INV_X1 DP_mult_215_U1223 ( .A(DP_mult_215_n1613), .ZN(DP_mult_215_n1618) );
  INV_X1 DP_mult_215_U1222 ( .A(DP_mult_215_n1613), .ZN(DP_mult_215_n1617) );
  INV_X1 DP_mult_215_U1221 ( .A(DP_mult_215_n1612), .ZN(DP_mult_215_n1616) );
  CLKBUF_X1 DP_mult_215_U1220 ( .A(DP_sw1_23_), .Z(DP_mult_215_n1614) );
  CLKBUF_X1 DP_mult_215_U1219 ( .A(DP_sw1_23_), .Z(DP_mult_215_n1613) );
  CLKBUF_X1 DP_mult_215_U1218 ( .A(DP_sw1_23_), .Z(DP_mult_215_n1612) );
  BUF_X1 DP_mult_215_U1217 ( .A(DP_mult_215_n1647), .Z(DP_mult_215_n1567) );
  BUF_X1 DP_mult_215_U1216 ( .A(DP_mult_215_n1647), .Z(DP_mult_215_n1566) );
  BUF_X1 DP_mult_215_U1215 ( .A(DP_mult_215_n1647), .Z(DP_mult_215_n1565) );
  INV_X1 DP_mult_215_U1214 ( .A(DP_mult_215_n1616), .ZN(DP_mult_215_n1615) );
  AND2_X1 DP_mult_215_U1213 ( .A1(DP_coeff_ret1[0]), .A2(DP_mult_215_n2157), 
        .ZN(DP_mult_215_n1555) );
  BUF_X1 DP_mult_215_U1212 ( .A(DP_mult_215_n1636), .Z(DP_mult_215_n1562) );
  OR2_X1 DP_mult_215_U1211 ( .A1(DP_mult_215_n2158), .A2(DP_mult_215_n2157), 
        .ZN(DP_mult_215_n1554) );
  BUF_X1 DP_mult_215_U1210 ( .A(DP_mult_215_n1636), .Z(DP_mult_215_n1563) );
  INV_X1 DP_mult_215_U1209 ( .A(DP_mult_215_n1555), .ZN(DP_mult_215_n1564) );
  NAND3_X1 DP_mult_215_U1208 ( .A1(DP_mult_215_n2157), .A2(DP_mult_215_n2158), 
        .A3(DP_mult_215_n2159), .ZN(DP_mult_215_n1639) );
  INV_X1 DP_mult_215_U1207 ( .A(DP_coeff_ret1[23]), .ZN(DP_mult_215_n1611) );
  INV_X1 DP_mult_215_U1206 ( .A(DP_coeff_ret1[8]), .ZN(DP_mult_215_n1601) );
  INV_X1 DP_mult_215_U1205 ( .A(DP_coeff_ret1[5]), .ZN(DP_mult_215_n1599) );
  OR2_X1 DP_mult_215_U1204 ( .A1(DP_mult_215_n1738), .A2(DP_mult_215_n1739), 
        .ZN(DP_mult_215_n1553) );
  OR2_X1 DP_mult_215_U1203 ( .A1(DP_mult_215_n1740), .A2(DP_mult_215_n1741), 
        .ZN(DP_mult_215_n1552) );
  INV_X1 DP_mult_215_U1202 ( .A(DP_mult_215_n1554), .ZN(DP_mult_215_n1561) );
  INV_X1 DP_mult_215_U1201 ( .A(DP_mult_215_n1611), .ZN(DP_mult_215_n1610) );
  BUF_X1 DP_mult_215_U1200 ( .A(DP_coeff_ret1[20]), .Z(DP_mult_215_n1609) );
  AND2_X1 DP_mult_215_U1199 ( .A1(DP_mult_215_n1738), .A2(DP_mult_215_n1740), 
        .ZN(DP_mult_215_n1551) );
  BUF_X1 DP_mult_215_U1198 ( .A(DP_mult_215_n1654), .Z(DP_mult_215_n1572) );
  BUF_X1 DP_mult_215_U1197 ( .A(DP_mult_215_n1654), .Z(DP_mult_215_n1571) );
  INV_X1 DP_mult_215_U1196 ( .A(DP_mult_215_n1552), .ZN(DP_mult_215_n1569) );
  INV_X1 DP_mult_215_U1195 ( .A(DP_mult_215_n1553), .ZN(DP_mult_215_n1570) );
  INV_X1 DP_mult_215_U1194 ( .A(DP_mult_215_n1601), .ZN(DP_mult_215_n1600) );
  INV_X1 DP_mult_215_U1193 ( .A(DP_mult_215_n1599), .ZN(DP_mult_215_n1598) );
  INV_X1 DP_mult_215_U1192 ( .A(DP_coeff_ret1[17]), .ZN(DP_mult_215_n1607) );
  INV_X1 DP_mult_215_U1191 ( .A(DP_coeff_ret1[11]), .ZN(DP_mult_215_n1603) );
  OR2_X1 DP_mult_215_U1190 ( .A1(DP_mult_215_n2070), .A2(DP_mult_215_n2069), 
        .ZN(DP_mult_215_n1550) );
  AND2_X1 DP_mult_215_U1189 ( .A1(DP_mult_215_n2070), .A2(DP_mult_215_n2068), 
        .ZN(DP_mult_215_n1549) );
  OR2_X1 DP_mult_215_U1188 ( .A1(DP_mult_215_n2068), .A2(DP_mult_215_n2067), 
        .ZN(DP_mult_215_n1548) );
  BUF_X1 DP_mult_215_U1187 ( .A(DP_coeff_ret1[20]), .Z(DP_mult_215_n1608) );
  INV_X1 DP_mult_215_U1186 ( .A(DP_coeff_ret1[14]), .ZN(DP_mult_215_n1605) );
  OR2_X1 DP_mult_215_U1185 ( .A1(DP_mult_215_n1794), .A2(DP_mult_215_n1795), 
        .ZN(DP_mult_215_n1547) );
  AND2_X1 DP_mult_215_U1184 ( .A1(DP_mult_215_n1794), .A2(DP_mult_215_n1796), 
        .ZN(DP_mult_215_n1546) );
  OR2_X1 DP_mult_215_U1183 ( .A1(DP_mult_215_n1851), .A2(DP_mult_215_n1852), 
        .ZN(DP_mult_215_n1545) );
  OR2_X1 DP_mult_215_U1182 ( .A1(DP_mult_215_n1796), .A2(DP_mult_215_n1797), 
        .ZN(DP_mult_215_n1544) );
  BUF_X1 DP_mult_215_U1181 ( .A(DP_mult_215_n1629), .Z(DP_mult_215_n1556) );
  INV_X1 DP_mult_215_U1180 ( .A(DP_mult_215_n1551), .ZN(DP_mult_215_n1568) );
  INV_X1 DP_mult_215_U1179 ( .A(DP_mult_215_n1605), .ZN(DP_mult_215_n1604) );
  INV_X1 DP_mult_215_U1178 ( .A(DP_mult_215_n1603), .ZN(DP_mult_215_n1602) );
  OR2_X1 DP_mult_215_U1177 ( .A1(DP_mult_215_n2014), .A2(DP_mult_215_n2015), 
        .ZN(DP_mult_215_n1543) );
  AND2_X1 DP_mult_215_U1176 ( .A1(DP_mult_215_n2014), .A2(DP_mult_215_n2016), 
        .ZN(DP_mult_215_n1542) );
  OR2_X1 DP_mult_215_U1175 ( .A1(DP_mult_215_n2016), .A2(DP_mult_215_n2017), 
        .ZN(DP_mult_215_n1541) );
  BUF_X1 DP_mult_215_U1174 ( .A(DP_mult_215_n1629), .Z(DP_mult_215_n1557) );
  INV_X1 DP_mult_215_U1173 ( .A(DP_mult_215_n1548), .ZN(DP_mult_215_n1559) );
  INV_X1 DP_mult_215_U1172 ( .A(DP_mult_215_n1549), .ZN(DP_mult_215_n1558) );
  INV_X1 DP_mult_215_U1171 ( .A(DP_mult_215_n1550), .ZN(DP_mult_215_n1560) );
  INV_X1 DP_mult_215_U1170 ( .A(DP_mult_215_n1607), .ZN(DP_mult_215_n1606) );
  INV_X1 DP_mult_215_U1169 ( .A(DP_mult_215_n1545), .ZN(DP_mult_215_n1579) );
  INV_X1 DP_mult_215_U1168 ( .A(DP_mult_215_n1544), .ZN(DP_mult_215_n1574) );
  OR2_X1 DP_mult_215_U1167 ( .A1(DP_mult_215_n1959), .A2(DP_mult_215_n1960), 
        .ZN(DP_mult_215_n1540) );
  OR2_X1 DP_mult_215_U1166 ( .A1(DP_mult_215_n1904), .A2(DP_mult_215_n1905), 
        .ZN(DP_mult_215_n1539) );
  OR2_X1 DP_mult_215_U1165 ( .A1(DP_mult_215_n1849), .A2(DP_mult_215_n1850), 
        .ZN(DP_mult_215_n1538) );
  BUF_X1 DP_mult_215_U1164 ( .A(DP_mult_215_n1802), .Z(DP_mult_215_n1582) );
  BUF_X1 DP_mult_215_U1163 ( .A(DP_mult_215_n1747), .Z(DP_mult_215_n1577) );
  BUF_X1 DP_mult_215_U1162 ( .A(DP_mult_215_n1802), .Z(DP_mult_215_n1581) );
  BUF_X1 DP_mult_215_U1161 ( .A(DP_mult_215_n1747), .Z(DP_mult_215_n1576) );
  INV_X1 DP_mult_215_U1160 ( .A(DP_mult_215_n1546), .ZN(DP_mult_215_n1573) );
  INV_X1 DP_mult_215_U1159 ( .A(DP_mult_215_n1541), .ZN(DP_mult_215_n1594) );
  INV_X1 DP_mult_215_U1158 ( .A(DP_mult_215_n1547), .ZN(DP_mult_215_n1575) );
  AND2_X1 DP_mult_215_U1157 ( .A1(DP_mult_215_n1959), .A2(DP_mult_215_n1961), 
        .ZN(DP_mult_215_n1537) );
  AND2_X1 DP_mult_215_U1156 ( .A1(DP_mult_215_n1904), .A2(DP_mult_215_n1906), 
        .ZN(DP_mult_215_n1536) );
  AND2_X1 DP_mult_215_U1155 ( .A1(DP_mult_215_n1849), .A2(DP_mult_215_n1851), 
        .ZN(DP_mult_215_n1535) );
  OR2_X1 DP_mult_215_U1154 ( .A1(DP_mult_215_n1961), .A2(DP_mult_215_n1962), 
        .ZN(DP_mult_215_n1534) );
  OR2_X1 DP_mult_215_U1153 ( .A1(DP_mult_215_n1906), .A2(DP_mult_215_n1907), 
        .ZN(DP_mult_215_n1533) );
  BUF_X1 DP_mult_215_U1152 ( .A(DP_mult_215_n1967), .Z(DP_mult_215_n1597) );
  BUF_X1 DP_mult_215_U1151 ( .A(DP_mult_215_n1967), .Z(DP_mult_215_n1596) );
  INV_X1 DP_mult_215_U1150 ( .A(DP_mult_215_n1542), .ZN(DP_mult_215_n1593) );
  INV_X1 DP_mult_215_U1149 ( .A(DP_mult_215_n1543), .ZN(DP_mult_215_n1595) );
  BUF_X1 DP_mult_215_U1148 ( .A(DP_mult_215_n1857), .Z(DP_mult_215_n1587) );
  INV_X1 DP_mult_215_U1147 ( .A(DP_mult_215_n1534), .ZN(DP_mult_215_n1589) );
  INV_X1 DP_mult_215_U1146 ( .A(DP_mult_215_n1533), .ZN(DP_mult_215_n1584) );
  INV_X1 DP_mult_215_U1145 ( .A(DP_mult_215_n1540), .ZN(DP_mult_215_n1590) );
  INV_X1 DP_mult_215_U1144 ( .A(DP_mult_215_n1539), .ZN(DP_mult_215_n1585) );
  INV_X1 DP_mult_215_U1143 ( .A(DP_mult_215_n1538), .ZN(DP_mult_215_n1580) );
  BUF_X1 DP_mult_215_U1142 ( .A(DP_mult_215_n1912), .Z(DP_mult_215_n1592) );
  BUF_X1 DP_mult_215_U1141 ( .A(DP_mult_215_n1912), .Z(DP_mult_215_n1591) );
  BUF_X1 DP_mult_215_U1140 ( .A(DP_mult_215_n1857), .Z(DP_mult_215_n1586) );
  INV_X1 DP_mult_215_U1139 ( .A(DP_mult_215_n1536), .ZN(DP_mult_215_n1583) );
  INV_X1 DP_mult_215_U1138 ( .A(DP_mult_215_n1537), .ZN(DP_mult_215_n1588) );
  INV_X1 DP_mult_215_U1137 ( .A(DP_mult_215_n1535), .ZN(DP_mult_215_n1578) );
  HA_X1 DP_mult_215_U1134 ( .A(DP_sw1_0_), .B(DP_sw1_1_), .CO(DP_mult_215_n727), .S(DP_mult_215_n1397) );
  FA_X1 DP_mult_215_U1133 ( .A(DP_sw1_1_), .B(DP_sw1_2_), .CI(DP_mult_215_n727), .CO(DP_mult_215_n726), .S(DP_mult_215_n1396) );
  FA_X1 DP_mult_215_U1132 ( .A(DP_sw1_2_), .B(DP_sw1_3_), .CI(DP_mult_215_n726), .CO(DP_mult_215_n725), .S(DP_mult_215_n1395) );
  FA_X1 DP_mult_215_U1131 ( .A(DP_sw1_3_), .B(DP_sw1_4_), .CI(DP_mult_215_n725), .CO(DP_mult_215_n724), .S(DP_mult_215_n1394) );
  FA_X1 DP_mult_215_U1130 ( .A(DP_sw1_4_), .B(DP_sw1_5_), .CI(DP_mult_215_n724), .CO(DP_mult_215_n723), .S(DP_mult_215_n1393) );
  FA_X1 DP_mult_215_U1129 ( .A(DP_sw1_5_), .B(DP_sw1_6_), .CI(DP_mult_215_n723), .CO(DP_mult_215_n722), .S(DP_mult_215_n1392) );
  FA_X1 DP_mult_215_U1128 ( .A(DP_sw1_6_), .B(DP_sw1_7_), .CI(DP_mult_215_n722), .CO(DP_mult_215_n721), .S(DP_mult_215_n1391) );
  FA_X1 DP_mult_215_U1127 ( .A(DP_sw1_7_), .B(DP_sw1_8_), .CI(DP_mult_215_n721), .CO(DP_mult_215_n720), .S(DP_mult_215_n1390) );
  FA_X1 DP_mult_215_U1126 ( .A(DP_sw1_8_), .B(DP_sw1_9_), .CI(DP_mult_215_n720), .CO(DP_mult_215_n719), .S(DP_mult_215_n1389) );
  FA_X1 DP_mult_215_U1125 ( .A(DP_sw1_9_), .B(DP_sw1_10_), .CI(
        DP_mult_215_n719), .CO(DP_mult_215_n718), .S(DP_mult_215_n1388) );
  FA_X1 DP_mult_215_U1124 ( .A(DP_sw1_10_), .B(DP_sw1_11_), .CI(
        DP_mult_215_n718), .CO(DP_mult_215_n717), .S(DP_mult_215_n1387) );
  FA_X1 DP_mult_215_U1123 ( .A(DP_sw1_11_), .B(DP_sw1_12_), .CI(
        DP_mult_215_n717), .CO(DP_mult_215_n716), .S(DP_mult_215_n1386) );
  FA_X1 DP_mult_215_U1122 ( .A(DP_sw1_12_), .B(DP_sw1_13_), .CI(
        DP_mult_215_n716), .CO(DP_mult_215_n715), .S(DP_mult_215_n1385) );
  FA_X1 DP_mult_215_U1121 ( .A(DP_sw1_13_), .B(DP_sw1_14_), .CI(
        DP_mult_215_n715), .CO(DP_mult_215_n714), .S(DP_mult_215_n1384) );
  FA_X1 DP_mult_215_U1120 ( .A(DP_sw1_14_), .B(DP_sw1_15_), .CI(
        DP_mult_215_n714), .CO(DP_mult_215_n713), .S(DP_mult_215_n1383) );
  FA_X1 DP_mult_215_U1119 ( .A(DP_sw1_15_), .B(DP_sw1_16_), .CI(
        DP_mult_215_n713), .CO(DP_mult_215_n712), .S(DP_mult_215_n1382) );
  FA_X1 DP_mult_215_U1118 ( .A(DP_sw1_16_), .B(DP_sw1_17_), .CI(
        DP_mult_215_n712), .CO(DP_mult_215_n711), .S(DP_mult_215_n1381) );
  FA_X1 DP_mult_215_U1117 ( .A(DP_sw1_17_), .B(DP_sw1_18_), .CI(
        DP_mult_215_n711), .CO(DP_mult_215_n710), .S(DP_mult_215_n1380) );
  FA_X1 DP_mult_215_U1116 ( .A(DP_sw1_18_), .B(DP_sw1_19_), .CI(
        DP_mult_215_n710), .CO(DP_mult_215_n709), .S(DP_mult_215_n1379) );
  FA_X1 DP_mult_215_U1115 ( .A(DP_sw1_19_), .B(DP_sw1_20_), .CI(
        DP_mult_215_n709), .CO(DP_mult_215_n708), .S(DP_mult_215_n1378) );
  FA_X1 DP_mult_215_U1114 ( .A(DP_sw1_20_), .B(DP_sw1_21_), .CI(
        DP_mult_215_n708), .CO(DP_mult_215_n707), .S(DP_mult_215_n1377) );
  FA_X1 DP_mult_215_U1113 ( .A(DP_sw1_21_), .B(DP_sw1_22_), .CI(
        DP_mult_215_n707), .CO(DP_mult_215_n706), .S(DP_mult_215_n1376) );
  FA_X1 DP_mult_215_U1112 ( .A(DP_sw1_22_), .B(DP_mult_215_n1615), .CI(
        DP_mult_215_n706), .CO(DP_mult_215_n1374), .S(DP_mult_215_n1375) );
  HA_X1 DP_mult_215_U408 ( .A(DP_mult_215_n904), .B(DP_mult_215_n1598), .CO(
        DP_mult_215_n687), .S(DP_mult_215_n688) );
  HA_X1 DP_mult_215_U407 ( .A(DP_mult_215_n687), .B(DP_mult_215_n903), .CO(
        DP_mult_215_n685), .S(DP_mult_215_n686) );
  HA_X1 DP_mult_215_U406 ( .A(DP_mult_215_n685), .B(DP_mult_215_n902), .CO(
        DP_mult_215_n683), .S(DP_mult_215_n684) );
  HA_X1 DP_mult_215_U405 ( .A(DP_mult_215_n878), .B(DP_mult_215_n1600), .CO(
        DP_mult_215_n681), .S(DP_mult_215_n682) );
  FA_X1 DP_mult_215_U404 ( .A(DP_mult_215_n901), .B(DP_mult_215_n682), .CI(
        DP_mult_215_n683), .CO(DP_mult_215_n679), .S(DP_mult_215_n680) );
  HA_X1 DP_mult_215_U403 ( .A(DP_mult_215_n681), .B(DP_mult_215_n877), .CO(
        DP_mult_215_n677), .S(DP_mult_215_n678) );
  FA_X1 DP_mult_215_U402 ( .A(DP_mult_215_n900), .B(DP_mult_215_n678), .CI(
        DP_mult_215_n679), .CO(DP_mult_215_n675), .S(DP_mult_215_n676) );
  HA_X1 DP_mult_215_U401 ( .A(DP_mult_215_n677), .B(DP_mult_215_n876), .CO(
        DP_mult_215_n673), .S(DP_mult_215_n674) );
  FA_X1 DP_mult_215_U400 ( .A(DP_mult_215_n899), .B(DP_mult_215_n674), .CI(
        DP_mult_215_n675), .CO(DP_mult_215_n671), .S(DP_mult_215_n672) );
  HA_X1 DP_mult_215_U399 ( .A(DP_mult_215_n852), .B(DP_mult_215_n1602), .CO(
        DP_mult_215_n669), .S(DP_mult_215_n670) );
  FA_X1 DP_mult_215_U398 ( .A(DP_mult_215_n875), .B(DP_mult_215_n670), .CI(
        DP_mult_215_n673), .CO(DP_mult_215_n667), .S(DP_mult_215_n668) );
  FA_X1 DP_mult_215_U397 ( .A(DP_mult_215_n898), .B(DP_mult_215_n668), .CI(
        DP_mult_215_n671), .CO(DP_mult_215_n665), .S(DP_mult_215_n666) );
  HA_X1 DP_mult_215_U396 ( .A(DP_mult_215_n669), .B(DP_mult_215_n851), .CO(
        DP_mult_215_n663), .S(DP_mult_215_n664) );
  FA_X1 DP_mult_215_U395 ( .A(DP_mult_215_n874), .B(DP_mult_215_n664), .CI(
        DP_mult_215_n667), .CO(DP_mult_215_n661), .S(DP_mult_215_n662) );
  FA_X1 DP_mult_215_U394 ( .A(DP_mult_215_n897), .B(DP_mult_215_n662), .CI(
        DP_mult_215_n665), .CO(DP_mult_215_n659), .S(DP_mult_215_n660) );
  HA_X1 DP_mult_215_U393 ( .A(DP_mult_215_n663), .B(DP_mult_215_n850), .CO(
        DP_mult_215_n657), .S(DP_mult_215_n658) );
  FA_X1 DP_mult_215_U392 ( .A(DP_mult_215_n873), .B(DP_mult_215_n658), .CI(
        DP_mult_215_n661), .CO(DP_mult_215_n655), .S(DP_mult_215_n656) );
  FA_X1 DP_mult_215_U391 ( .A(DP_mult_215_n896), .B(DP_mult_215_n656), .CI(
        DP_mult_215_n659), .CO(DP_mult_215_n653), .S(DP_mult_215_n654) );
  HA_X1 DP_mult_215_U390 ( .A(DP_mult_215_n826), .B(DP_mult_215_n1604), .CO(
        DP_mult_215_n651), .S(DP_mult_215_n652) );
  FA_X1 DP_mult_215_U389 ( .A(DP_mult_215_n849), .B(DP_mult_215_n652), .CI(
        DP_mult_215_n657), .CO(DP_mult_215_n649), .S(DP_mult_215_n650) );
  FA_X1 DP_mult_215_U388 ( .A(DP_mult_215_n872), .B(DP_mult_215_n650), .CI(
        DP_mult_215_n655), .CO(DP_mult_215_n647), .S(DP_mult_215_n648) );
  FA_X1 DP_mult_215_U387 ( .A(DP_mult_215_n895), .B(DP_mult_215_n648), .CI(
        DP_mult_215_n653), .CO(DP_mult_215_n645), .S(DP_mult_215_n646) );
  HA_X1 DP_mult_215_U386 ( .A(DP_mult_215_n651), .B(DP_mult_215_n825), .CO(
        DP_mult_215_n643), .S(DP_mult_215_n644) );
  FA_X1 DP_mult_215_U385 ( .A(DP_mult_215_n848), .B(DP_mult_215_n644), .CI(
        DP_mult_215_n649), .CO(DP_mult_215_n641), .S(DP_mult_215_n642) );
  FA_X1 DP_mult_215_U384 ( .A(DP_mult_215_n871), .B(DP_mult_215_n642), .CI(
        DP_mult_215_n647), .CO(DP_mult_215_n639), .S(DP_mult_215_n640) );
  FA_X1 DP_mult_215_U383 ( .A(DP_mult_215_n894), .B(DP_mult_215_n640), .CI(
        DP_mult_215_n645), .CO(DP_mult_215_n637), .S(DP_mult_215_n638) );
  HA_X1 DP_mult_215_U382 ( .A(DP_mult_215_n643), .B(DP_mult_215_n824), .CO(
        DP_mult_215_n635), .S(DP_mult_215_n636) );
  FA_X1 DP_mult_215_U381 ( .A(DP_mult_215_n847), .B(DP_mult_215_n636), .CI(
        DP_mult_215_n641), .CO(DP_mult_215_n633), .S(DP_mult_215_n634) );
  FA_X1 DP_mult_215_U380 ( .A(DP_mult_215_n870), .B(DP_mult_215_n634), .CI(
        DP_mult_215_n639), .CO(DP_mult_215_n631), .S(DP_mult_215_n632) );
  FA_X1 DP_mult_215_U379 ( .A(DP_mult_215_n893), .B(DP_mult_215_n632), .CI(
        DP_mult_215_n637), .CO(DP_mult_215_n629), .S(DP_mult_215_n630) );
  HA_X1 DP_mult_215_U378 ( .A(DP_mult_215_n800), .B(DP_mult_215_n1606), .CO(
        DP_mult_215_n627), .S(DP_mult_215_n628) );
  FA_X1 DP_mult_215_U377 ( .A(DP_mult_215_n823), .B(DP_mult_215_n628), .CI(
        DP_mult_215_n635), .CO(DP_mult_215_n625), .S(DP_mult_215_n626) );
  FA_X1 DP_mult_215_U376 ( .A(DP_mult_215_n846), .B(DP_mult_215_n626), .CI(
        DP_mult_215_n633), .CO(DP_mult_215_n623), .S(DP_mult_215_n624) );
  FA_X1 DP_mult_215_U375 ( .A(DP_mult_215_n869), .B(DP_mult_215_n624), .CI(
        DP_mult_215_n631), .CO(DP_mult_215_n621), .S(DP_mult_215_n622) );
  FA_X1 DP_mult_215_U374 ( .A(DP_mult_215_n892), .B(DP_mult_215_n622), .CI(
        DP_mult_215_n629), .CO(DP_mult_215_n619), .S(DP_mult_215_n620) );
  HA_X1 DP_mult_215_U373 ( .A(DP_mult_215_n627), .B(DP_mult_215_n799), .CO(
        DP_mult_215_n617), .S(DP_mult_215_n618) );
  FA_X1 DP_mult_215_U372 ( .A(DP_mult_215_n822), .B(DP_mult_215_n618), .CI(
        DP_mult_215_n625), .CO(DP_mult_215_n615), .S(DP_mult_215_n616) );
  FA_X1 DP_mult_215_U371 ( .A(DP_mult_215_n845), .B(DP_mult_215_n616), .CI(
        DP_mult_215_n623), .CO(DP_mult_215_n613), .S(DP_mult_215_n614) );
  FA_X1 DP_mult_215_U370 ( .A(DP_mult_215_n868), .B(DP_mult_215_n614), .CI(
        DP_mult_215_n621), .CO(DP_mult_215_n611), .S(DP_mult_215_n612) );
  FA_X1 DP_mult_215_U369 ( .A(DP_mult_215_n891), .B(DP_mult_215_n612), .CI(
        DP_mult_215_n619), .CO(DP_mult_215_n609), .S(DP_mult_215_n610) );
  HA_X1 DP_mult_215_U368 ( .A(DP_mult_215_n617), .B(DP_mult_215_n798), .CO(
        DP_mult_215_n607), .S(DP_mult_215_n608) );
  FA_X1 DP_mult_215_U367 ( .A(DP_mult_215_n821), .B(DP_mult_215_n608), .CI(
        DP_mult_215_n615), .CO(DP_mult_215_n605), .S(DP_mult_215_n606) );
  FA_X1 DP_mult_215_U366 ( .A(DP_mult_215_n844), .B(DP_mult_215_n606), .CI(
        DP_mult_215_n613), .CO(DP_mult_215_n603), .S(DP_mult_215_n604) );
  FA_X1 DP_mult_215_U365 ( .A(DP_mult_215_n867), .B(DP_mult_215_n604), .CI(
        DP_mult_215_n611), .CO(DP_mult_215_n601), .S(DP_mult_215_n602) );
  FA_X1 DP_mult_215_U364 ( .A(DP_mult_215_n890), .B(DP_mult_215_n602), .CI(
        DP_mult_215_n609), .CO(DP_mult_215_n599), .S(DP_mult_215_n600) );
  HA_X1 DP_mult_215_U363 ( .A(DP_mult_215_n774), .B(DP_mult_215_n1608), .CO(
        DP_mult_215_n597), .S(DP_mult_215_n598) );
  FA_X1 DP_mult_215_U362 ( .A(DP_mult_215_n797), .B(DP_mult_215_n598), .CI(
        DP_mult_215_n607), .CO(DP_mult_215_n595), .S(DP_mult_215_n596) );
  FA_X1 DP_mult_215_U361 ( .A(DP_mult_215_n820), .B(DP_mult_215_n596), .CI(
        DP_mult_215_n605), .CO(DP_mult_215_n593), .S(DP_mult_215_n594) );
  FA_X1 DP_mult_215_U360 ( .A(DP_mult_215_n843), .B(DP_mult_215_n594), .CI(
        DP_mult_215_n603), .CO(DP_mult_215_n591), .S(DP_mult_215_n592) );
  FA_X1 DP_mult_215_U359 ( .A(DP_mult_215_n866), .B(DP_mult_215_n592), .CI(
        DP_mult_215_n601), .CO(DP_mult_215_n589), .S(DP_mult_215_n590) );
  FA_X1 DP_mult_215_U358 ( .A(DP_mult_215_n889), .B(DP_mult_215_n590), .CI(
        DP_mult_215_n599), .CO(DP_mult_215_n587), .S(DP_mult_215_n588) );
  HA_X1 DP_mult_215_U357 ( .A(DP_mult_215_n597), .B(DP_mult_215_n773), .CO(
        DP_mult_215_n585), .S(DP_mult_215_n586) );
  FA_X1 DP_mult_215_U356 ( .A(DP_mult_215_n796), .B(DP_mult_215_n586), .CI(
        DP_mult_215_n595), .CO(DP_mult_215_n583), .S(DP_mult_215_n584) );
  FA_X1 DP_mult_215_U355 ( .A(DP_mult_215_n819), .B(DP_mult_215_n584), .CI(
        DP_mult_215_n593), .CO(DP_mult_215_n581), .S(DP_mult_215_n582) );
  FA_X1 DP_mult_215_U354 ( .A(DP_mult_215_n842), .B(DP_mult_215_n582), .CI(
        DP_mult_215_n591), .CO(DP_mult_215_n579), .S(DP_mult_215_n580) );
  FA_X1 DP_mult_215_U353 ( .A(DP_mult_215_n865), .B(DP_mult_215_n580), .CI(
        DP_mult_215_n589), .CO(DP_mult_215_n577), .S(DP_mult_215_n578) );
  FA_X1 DP_mult_215_U352 ( .A(DP_mult_215_n888), .B(DP_mult_215_n578), .CI(
        DP_mult_215_n587), .CO(DP_mult_215_n575), .S(DP_mult_215_n576) );
  HA_X1 DP_mult_215_U351 ( .A(DP_mult_215_n585), .B(DP_mult_215_n772), .CO(
        DP_mult_215_n573), .S(DP_mult_215_n574) );
  FA_X1 DP_mult_215_U350 ( .A(DP_mult_215_n795), .B(DP_mult_215_n574), .CI(
        DP_mult_215_n583), .CO(DP_mult_215_n571), .S(DP_mult_215_n572) );
  FA_X1 DP_mult_215_U349 ( .A(DP_mult_215_n818), .B(DP_mult_215_n572), .CI(
        DP_mult_215_n581), .CO(DP_mult_215_n569), .S(DP_mult_215_n570) );
  FA_X1 DP_mult_215_U348 ( .A(DP_mult_215_n841), .B(DP_mult_215_n570), .CI(
        DP_mult_215_n579), .CO(DP_mult_215_n567), .S(DP_mult_215_n568) );
  FA_X1 DP_mult_215_U347 ( .A(DP_mult_215_n864), .B(DP_mult_215_n568), .CI(
        DP_mult_215_n577), .CO(DP_mult_215_n565), .S(DP_mult_215_n566) );
  FA_X1 DP_mult_215_U346 ( .A(DP_mult_215_n887), .B(DP_mult_215_n566), .CI(
        DP_mult_215_n575), .CO(DP_mult_215_n563), .S(DP_mult_215_n564) );
  HA_X1 DP_mult_215_U345 ( .A(DP_mult_215_n748), .B(DP_mult_215_n1610), .CO(
        DP_mult_215_n561), .S(DP_mult_215_n562) );
  FA_X1 DP_mult_215_U344 ( .A(DP_mult_215_n771), .B(DP_mult_215_n562), .CI(
        DP_mult_215_n573), .CO(DP_mult_215_n559), .S(DP_mult_215_n560) );
  FA_X1 DP_mult_215_U343 ( .A(DP_mult_215_n794), .B(DP_mult_215_n560), .CI(
        DP_mult_215_n571), .CO(DP_mult_215_n557), .S(DP_mult_215_n558) );
  FA_X1 DP_mult_215_U342 ( .A(DP_mult_215_n817), .B(DP_mult_215_n558), .CI(
        DP_mult_215_n569), .CO(DP_mult_215_n555), .S(DP_mult_215_n556) );
  FA_X1 DP_mult_215_U341 ( .A(DP_mult_215_n840), .B(DP_mult_215_n556), .CI(
        DP_mult_215_n567), .CO(DP_mult_215_n553), .S(DP_mult_215_n554) );
  FA_X1 DP_mult_215_U340 ( .A(DP_mult_215_n863), .B(DP_mult_215_n554), .CI(
        DP_mult_215_n565), .CO(DP_mult_215_n551), .S(DP_mult_215_n552) );
  FA_X1 DP_mult_215_U339 ( .A(DP_mult_215_n886), .B(DP_mult_215_n552), .CI(
        DP_mult_215_n563), .CO(DP_mult_215_n549), .S(DP_mult_215_n550) );
  HA_X1 DP_mult_215_U338 ( .A(DP_mult_215_n561), .B(DP_mult_215_n747), .CO(
        DP_mult_215_n547), .S(DP_mult_215_n548) );
  FA_X1 DP_mult_215_U337 ( .A(DP_mult_215_n770), .B(DP_mult_215_n548), .CI(
        DP_mult_215_n559), .CO(DP_mult_215_n545), .S(DP_mult_215_n546) );
  FA_X1 DP_mult_215_U336 ( .A(DP_mult_215_n793), .B(DP_mult_215_n546), .CI(
        DP_mult_215_n557), .CO(DP_mult_215_n543), .S(DP_mult_215_n544) );
  FA_X1 DP_mult_215_U335 ( .A(DP_mult_215_n816), .B(DP_mult_215_n544), .CI(
        DP_mult_215_n555), .CO(DP_mult_215_n541), .S(DP_mult_215_n542) );
  FA_X1 DP_mult_215_U334 ( .A(DP_mult_215_n839), .B(DP_mult_215_n542), .CI(
        DP_mult_215_n553), .CO(DP_mult_215_n539), .S(DP_mult_215_n540) );
  FA_X1 DP_mult_215_U333 ( .A(DP_mult_215_n862), .B(DP_mult_215_n540), .CI(
        DP_mult_215_n551), .CO(DP_mult_215_n537), .S(DP_mult_215_n538) );
  FA_X1 DP_mult_215_U332 ( .A(DP_mult_215_n885), .B(DP_mult_215_n538), .CI(
        DP_mult_215_n549), .CO(DP_mult_215_n535), .S(DP_mult_215_n536) );
  HA_X1 DP_mult_215_U331 ( .A(DP_mult_215_n547), .B(DP_mult_215_n746), .CO(
        DP_mult_215_n533), .S(DP_mult_215_n534) );
  FA_X1 DP_mult_215_U330 ( .A(DP_mult_215_n769), .B(DP_mult_215_n534), .CI(
        DP_mult_215_n545), .CO(DP_mult_215_n531), .S(DP_mult_215_n532) );
  FA_X1 DP_mult_215_U329 ( .A(DP_mult_215_n792), .B(DP_mult_215_n532), .CI(
        DP_mult_215_n543), .CO(DP_mult_215_n529), .S(DP_mult_215_n530) );
  FA_X1 DP_mult_215_U328 ( .A(DP_mult_215_n815), .B(DP_mult_215_n530), .CI(
        DP_mult_215_n541), .CO(DP_mult_215_n527), .S(DP_mult_215_n528) );
  FA_X1 DP_mult_215_U327 ( .A(DP_mult_215_n838), .B(DP_mult_215_n528), .CI(
        DP_mult_215_n539), .CO(DP_mult_215_n525), .S(DP_mult_215_n526) );
  FA_X1 DP_mult_215_U326 ( .A(DP_mult_215_n861), .B(DP_mult_215_n526), .CI(
        DP_mult_215_n537), .CO(DP_mult_215_n523), .S(DP_mult_215_n524) );
  FA_X1 DP_mult_215_U325 ( .A(DP_mult_215_n884), .B(DP_mult_215_n524), .CI(
        DP_mult_215_n535), .CO(DP_mult_215_n521), .S(DP_mult_215_n522) );
  HA_X1 DP_mult_215_U324 ( .A(DP_mult_215_n533), .B(DP_mult_215_n745), .CO(
        DP_mult_215_n519), .S(DP_mult_215_n520) );
  FA_X1 DP_mult_215_U323 ( .A(DP_mult_215_n768), .B(DP_mult_215_n520), .CI(
        DP_mult_215_n531), .CO(DP_mult_215_n517), .S(DP_mult_215_n518) );
  FA_X1 DP_mult_215_U322 ( .A(DP_mult_215_n791), .B(DP_mult_215_n518), .CI(
        DP_mult_215_n529), .CO(DP_mult_215_n515), .S(DP_mult_215_n516) );
  FA_X1 DP_mult_215_U321 ( .A(DP_mult_215_n814), .B(DP_mult_215_n516), .CI(
        DP_mult_215_n527), .CO(DP_mult_215_n513), .S(DP_mult_215_n514) );
  FA_X1 DP_mult_215_U320 ( .A(DP_mult_215_n837), .B(DP_mult_215_n514), .CI(
        DP_mult_215_n525), .CO(DP_mult_215_n511), .S(DP_mult_215_n512) );
  FA_X1 DP_mult_215_U319 ( .A(DP_mult_215_n860), .B(DP_mult_215_n512), .CI(
        DP_mult_215_n523), .CO(DP_mult_215_n509), .S(DP_mult_215_n510) );
  FA_X1 DP_mult_215_U318 ( .A(DP_mult_215_n883), .B(DP_mult_215_n510), .CI(
        DP_mult_215_n521), .CO(DP_mult_215_n507), .S(DP_mult_215_n508) );
  FA_X1 DP_mult_215_U315 ( .A(DP_mult_215_n506), .B(DP_mult_215_n744), .CI(
        DP_mult_215_n767), .CO(DP_mult_215_n504), .S(DP_mult_215_n505) );
  FA_X1 DP_mult_215_U314 ( .A(DP_mult_215_n505), .B(DP_mult_215_n517), .CI(
        DP_mult_215_n790), .CO(DP_mult_215_n502), .S(DP_mult_215_n503) );
  FA_X1 DP_mult_215_U313 ( .A(DP_mult_215_n503), .B(DP_mult_215_n515), .CI(
        DP_mult_215_n813), .CO(DP_mult_215_n500), .S(DP_mult_215_n501) );
  FA_X1 DP_mult_215_U312 ( .A(DP_mult_215_n501), .B(DP_mult_215_n513), .CI(
        DP_mult_215_n836), .CO(DP_mult_215_n498), .S(DP_mult_215_n499) );
  FA_X1 DP_mult_215_U311 ( .A(DP_mult_215_n499), .B(DP_mult_215_n511), .CI(
        DP_mult_215_n859), .CO(DP_mult_215_n496), .S(DP_mult_215_n497) );
  FA_X1 DP_mult_215_U310 ( .A(DP_mult_215_n497), .B(DP_mult_215_n509), .CI(
        DP_mult_215_n882), .CO(DP_mult_215_n494), .S(DP_mult_215_n495) );
  FA_X1 DP_mult_215_U308 ( .A(DP_mult_215_n743), .B(DP_mult_215_n493), .CI(
        DP_mult_215_n766), .CO(DP_mult_215_n491), .S(DP_mult_215_n492) );
  FA_X1 DP_mult_215_U307 ( .A(DP_mult_215_n492), .B(DP_mult_215_n504), .CI(
        DP_mult_215_n789), .CO(DP_mult_215_n489), .S(DP_mult_215_n490) );
  FA_X1 DP_mult_215_U306 ( .A(DP_mult_215_n490), .B(DP_mult_215_n502), .CI(
        DP_mult_215_n500), .CO(DP_mult_215_n487), .S(DP_mult_215_n488) );
  FA_X1 DP_mult_215_U305 ( .A(DP_mult_215_n488), .B(DP_mult_215_n812), .CI(
        DP_mult_215_n835), .CO(DP_mult_215_n485), .S(DP_mult_215_n486) );
  FA_X1 DP_mult_215_U304 ( .A(DP_mult_215_n486), .B(DP_mult_215_n498), .CI(
        DP_mult_215_n496), .CO(DP_mult_215_n483), .S(DP_mult_215_n484) );
  FA_X1 DP_mult_215_U303 ( .A(DP_mult_215_n484), .B(DP_mult_215_n858), .CI(
        DP_mult_215_n881), .CO(DP_mult_215_n481), .S(DP_mult_215_n482) );
  FA_X1 DP_mult_215_U301 ( .A(DP_mult_215_n742), .B(DP_mult_215_n493), .CI(
        DP_mult_215_n491), .CO(DP_mult_215_n477), .S(DP_mult_215_n478) );
  FA_X1 DP_mult_215_U300 ( .A(DP_mult_215_n478), .B(DP_mult_215_n765), .CI(
        DP_mult_215_n788), .CO(DP_mult_215_n475), .S(DP_mult_215_n476) );
  FA_X1 DP_mult_215_U299 ( .A(DP_mult_215_n476), .B(DP_mult_215_n489), .CI(
        DP_mult_215_n487), .CO(DP_mult_215_n473), .S(DP_mult_215_n474) );
  FA_X1 DP_mult_215_U298 ( .A(DP_mult_215_n474), .B(DP_mult_215_n811), .CI(
        DP_mult_215_n834), .CO(DP_mult_215_n471), .S(DP_mult_215_n472) );
  FA_X1 DP_mult_215_U297 ( .A(DP_mult_215_n472), .B(DP_mult_215_n485), .CI(
        DP_mult_215_n483), .CO(DP_mult_215_n469), .S(DP_mult_215_n470) );
  FA_X1 DP_mult_215_U296 ( .A(DP_mult_215_n880), .B(DP_mult_215_n857), .CI(
        DP_mult_215_n470), .CO(DP_mult_215_n467), .S(DP_mult_215_n468) );
  FA_X1 DP_mult_215_U295 ( .A(DP_mult_215_n479), .B(DP_mult_215_n879), .CI(
        DP_mult_215_n741), .CO(DP_mult_215_n465), .S(DP_mult_215_n466) );
  FA_X1 DP_mult_215_U294 ( .A(DP_mult_215_n764), .B(DP_mult_215_n466), .CI(
        DP_mult_215_n477), .CO(DP_mult_215_n463), .S(DP_mult_215_n464) );
  FA_X1 DP_mult_215_U293 ( .A(DP_mult_215_n475), .B(DP_mult_215_n464), .CI(
        DP_mult_215_n787), .CO(DP_mult_215_n461), .S(DP_mult_215_n462) );
  FA_X1 DP_mult_215_U292 ( .A(DP_mult_215_n810), .B(DP_mult_215_n462), .CI(
        DP_mult_215_n473), .CO(DP_mult_215_n459), .S(DP_mult_215_n460) );
  FA_X1 DP_mult_215_U291 ( .A(DP_mult_215_n471), .B(DP_mult_215_n460), .CI(
        DP_mult_215_n833), .CO(DP_mult_215_n457), .S(DP_mult_215_n458) );
  FA_X1 DP_mult_215_U290 ( .A(DP_mult_215_n856), .B(DP_mult_215_n458), .CI(
        DP_mult_215_n469), .CO(DP_mult_215_n455), .S(DP_mult_215_n456) );
  FA_X1 DP_mult_215_U288 ( .A(DP_mult_215_n454), .B(DP_mult_215_n465), .CI(
        DP_mult_215_n763), .CO(DP_mult_215_n452), .S(DP_mult_215_n453) );
  FA_X1 DP_mult_215_U287 ( .A(DP_mult_215_n453), .B(DP_mult_215_n463), .CI(
        DP_mult_215_n786), .CO(DP_mult_215_n450), .S(DP_mult_215_n451) );
  FA_X1 DP_mult_215_U286 ( .A(DP_mult_215_n451), .B(DP_mult_215_n461), .CI(
        DP_mult_215_n809), .CO(DP_mult_215_n448), .S(DP_mult_215_n449) );
  FA_X1 DP_mult_215_U285 ( .A(DP_mult_215_n449), .B(DP_mult_215_n459), .CI(
        DP_mult_215_n832), .CO(DP_mult_215_n446), .S(DP_mult_215_n447) );
  FA_X1 DP_mult_215_U284 ( .A(DP_mult_215_n447), .B(DP_mult_215_n457), .CI(
        DP_mult_215_n855), .CO(DP_mult_215_n444), .S(DP_mult_215_n445) );
  FA_X1 DP_mult_215_U282 ( .A(DP_mult_215_n740), .B(DP_mult_215_n454), .CI(
        DP_mult_215_n762), .CO(DP_mult_215_n440), .S(DP_mult_215_n441) );
  FA_X1 DP_mult_215_U281 ( .A(DP_mult_215_n441), .B(DP_mult_215_n452), .CI(
        DP_mult_215_n450), .CO(DP_mult_215_n438), .S(DP_mult_215_n439) );
  FA_X1 DP_mult_215_U280 ( .A(DP_mult_215_n439), .B(DP_mult_215_n785), .CI(
        DP_mult_215_n808), .CO(DP_mult_215_n436), .S(DP_mult_215_n437) );
  FA_X1 DP_mult_215_U279 ( .A(DP_mult_215_n437), .B(DP_mult_215_n448), .CI(
        DP_mult_215_n446), .CO(DP_mult_215_n434), .S(DP_mult_215_n435) );
  FA_X1 DP_mult_215_U278 ( .A(DP_mult_215_n854), .B(DP_mult_215_n831), .CI(
        DP_mult_215_n435), .CO(DP_mult_215_n432), .S(DP_mult_215_n433) );
  FA_X1 DP_mult_215_U277 ( .A(DP_mult_215_n442), .B(DP_mult_215_n853), .CI(
        DP_mult_215_n739), .CO(DP_mult_215_n430), .S(DP_mult_215_n431) );
  FA_X1 DP_mult_215_U276 ( .A(DP_mult_215_n440), .B(DP_mult_215_n431), .CI(
        DP_mult_215_n761), .CO(DP_mult_215_n428), .S(DP_mult_215_n429) );
  FA_X1 DP_mult_215_U275 ( .A(DP_mult_215_n784), .B(DP_mult_215_n429), .CI(
        DP_mult_215_n438), .CO(DP_mult_215_n426), .S(DP_mult_215_n427) );
  FA_X1 DP_mult_215_U274 ( .A(DP_mult_215_n436), .B(DP_mult_215_n427), .CI(
        DP_mult_215_n807), .CO(DP_mult_215_n424), .S(DP_mult_215_n425) );
  FA_X1 DP_mult_215_U273 ( .A(DP_mult_215_n830), .B(DP_mult_215_n425), .CI(
        DP_mult_215_n434), .CO(DP_mult_215_n422), .S(DP_mult_215_n423) );
  FA_X1 DP_mult_215_U271 ( .A(DP_mult_215_n421), .B(DP_mult_215_n430), .CI(
        DP_mult_215_n760), .CO(DP_mult_215_n419), .S(DP_mult_215_n420) );
  FA_X1 DP_mult_215_U270 ( .A(DP_mult_215_n420), .B(DP_mult_215_n428), .CI(
        DP_mult_215_n783), .CO(DP_mult_215_n417), .S(DP_mult_215_n418) );
  FA_X1 DP_mult_215_U269 ( .A(DP_mult_215_n418), .B(DP_mult_215_n426), .CI(
        DP_mult_215_n806), .CO(DP_mult_215_n415), .S(DP_mult_215_n416) );
  FA_X1 DP_mult_215_U268 ( .A(DP_mult_215_n416), .B(DP_mult_215_n424), .CI(
        DP_mult_215_n829), .CO(DP_mult_215_n413), .S(DP_mult_215_n414) );
  FA_X1 DP_mult_215_U266 ( .A(DP_mult_215_n738), .B(DP_mult_215_n421), .CI(
        DP_mult_215_n419), .CO(DP_mult_215_n409), .S(DP_mult_215_n410) );
  FA_X1 DP_mult_215_U265 ( .A(DP_mult_215_n410), .B(DP_mult_215_n759), .CI(
        DP_mult_215_n782), .CO(DP_mult_215_n407), .S(DP_mult_215_n408) );
  FA_X1 DP_mult_215_U264 ( .A(DP_mult_215_n408), .B(DP_mult_215_n417), .CI(
        DP_mult_215_n415), .CO(DP_mult_215_n405), .S(DP_mult_215_n406) );
  FA_X1 DP_mult_215_U263 ( .A(DP_mult_215_n828), .B(DP_mult_215_n805), .CI(
        DP_mult_215_n406), .CO(DP_mult_215_n403), .S(DP_mult_215_n404) );
  FA_X1 DP_mult_215_U262 ( .A(DP_mult_215_n411), .B(DP_mult_215_n827), .CI(
        DP_mult_215_n737), .CO(DP_mult_215_n387), .S(DP_mult_215_n402) );
  FA_X1 DP_mult_215_U261 ( .A(DP_mult_215_n758), .B(DP_mult_215_n402), .CI(
        DP_mult_215_n409), .CO(DP_mult_215_n400), .S(DP_mult_215_n401) );
  FA_X1 DP_mult_215_U260 ( .A(DP_mult_215_n407), .B(DP_mult_215_n401), .CI(
        DP_mult_215_n781), .CO(DP_mult_215_n398), .S(DP_mult_215_n399) );
  FA_X1 DP_mult_215_U259 ( .A(DP_mult_215_n804), .B(DP_mult_215_n399), .CI(
        DP_mult_215_n405), .CO(DP_mult_215_n396), .S(DP_mult_215_n397) );
  FA_X1 DP_mult_215_U257 ( .A(DP_mult_215_n395), .B(DP_mult_215_n736), .CI(
        DP_mult_215_n757), .CO(DP_mult_215_n393), .S(DP_mult_215_n394) );
  FA_X1 DP_mult_215_U256 ( .A(DP_mult_215_n394), .B(DP_mult_215_n400), .CI(
        DP_mult_215_n780), .CO(DP_mult_215_n391), .S(DP_mult_215_n392) );
  FA_X1 DP_mult_215_U255 ( .A(DP_mult_215_n392), .B(DP_mult_215_n398), .CI(
        DP_mult_215_n803), .CO(DP_mult_215_n389), .S(DP_mult_215_n390) );
  FA_X1 DP_mult_215_U253 ( .A(DP_mult_215_n735), .B(DP_mult_215_n395), .CI(
        DP_mult_215_n756), .CO(DP_mult_215_n385), .S(DP_mult_215_n386) );
  FA_X1 DP_mult_215_U252 ( .A(DP_mult_215_n386), .B(DP_mult_215_n393), .CI(
        DP_mult_215_n391), .CO(DP_mult_215_n383), .S(DP_mult_215_n384) );
  FA_X1 DP_mult_215_U251 ( .A(DP_mult_215_n802), .B(DP_mult_215_n779), .CI(
        DP_mult_215_n384), .CO(DP_mult_215_n381), .S(DP_mult_215_n382) );
  FA_X1 DP_mult_215_U250 ( .A(DP_mult_215_n387), .B(DP_mult_215_n801), .CI(
        DP_mult_215_n734), .CO(DP_mult_215_n379), .S(DP_mult_215_n380) );
  FA_X1 DP_mult_215_U249 ( .A(DP_mult_215_n385), .B(DP_mult_215_n380), .CI(
        DP_mult_215_n755), .CO(DP_mult_215_n377), .S(DP_mult_215_n378) );
  FA_X1 DP_mult_215_U248 ( .A(DP_mult_215_n778), .B(DP_mult_215_n378), .CI(
        DP_mult_215_n383), .CO(DP_mult_215_n375), .S(DP_mult_215_n376) );
  FA_X1 DP_mult_215_U246 ( .A(DP_mult_215_n374), .B(DP_mult_215_n379), .CI(
        DP_mult_215_n754), .CO(DP_mult_215_n372), .S(DP_mult_215_n373) );
  FA_X1 DP_mult_215_U245 ( .A(DP_mult_215_n373), .B(DP_mult_215_n377), .CI(
        DP_mult_215_n777), .CO(DP_mult_215_n370), .S(DP_mult_215_n371) );
  FA_X1 DP_mult_215_U243 ( .A(DP_mult_215_n733), .B(DP_mult_215_n374), .CI(
        DP_mult_215_n372), .CO(DP_mult_215_n366), .S(DP_mult_215_n367) );
  FA_X1 DP_mult_215_U242 ( .A(DP_mult_215_n776), .B(DP_mult_215_n753), .CI(
        DP_mult_215_n367), .CO(DP_mult_215_n364), .S(DP_mult_215_n365) );
  FA_X1 DP_mult_215_U241 ( .A(DP_mult_215_n368), .B(DP_mult_215_n775), .CI(
        DP_mult_215_n732), .CO(DP_mult_215_n356), .S(DP_mult_215_n363) );
  FA_X1 DP_mult_215_U240 ( .A(DP_mult_215_n752), .B(DP_mult_215_n363), .CI(
        DP_mult_215_n366), .CO(DP_mult_215_n361), .S(DP_mult_215_n362) );
  FA_X1 DP_mult_215_U238 ( .A(DP_mult_215_n360), .B(DP_mult_215_n731), .CI(
        DP_mult_215_n751), .CO(DP_mult_215_n358), .S(DP_mult_215_n359) );
  FA_X1 DP_mult_215_U236 ( .A(DP_mult_215_n730), .B(DP_mult_215_n360), .CI(
        DP_mult_215_n750), .CO(DP_mult_215_n354), .S(DP_mult_215_n355) );
  FA_X1 DP_mult_215_U235 ( .A(DP_mult_215_n356), .B(DP_mult_215_n749), .CI(
        DP_mult_215_n729), .CO(DP_mult_215_n352), .S(DP_mult_215_n353) );
  FA_X1 DP_mult_215_U204 ( .A(DP_mult_215_n908), .B(DP_mult_215_n536), .CI(
        DP_mult_215_n326), .CO(DP_mult_215_n325), .S(DP_sw1_coeff_ret1[0]) );
  FA_X1 DP_mult_215_U203 ( .A(DP_mult_215_n907), .B(DP_mult_215_n522), .CI(
        DP_mult_215_n325), .CO(DP_mult_215_n324), .S(DP_sw1_coeff_ret1[1]) );
  FA_X1 DP_mult_215_U202 ( .A(DP_mult_215_n508), .B(DP_mult_215_n906), .CI(
        DP_mult_215_n324), .CO(DP_mult_215_n323), .S(DP_sw1_coeff_ret1[2]) );
  FA_X1 DP_mult_215_U201 ( .A(DP_mult_215_n495), .B(DP_mult_215_n507), .CI(
        DP_mult_215_n323), .CO(DP_mult_215_n322), .S(DP_sw1_coeff_ret1[3]) );
  FA_X1 DP_mult_215_U200 ( .A(DP_mult_215_n482), .B(DP_mult_215_n494), .CI(
        DP_mult_215_n322), .CO(DP_mult_215_n321), .S(DP_sw1_coeff_ret1[4]) );
  FA_X1 DP_mult_215_U199 ( .A(DP_mult_215_n468), .B(DP_mult_215_n481), .CI(
        DP_mult_215_n321), .CO(DP_mult_215_n320), .S(DP_sw1_coeff_ret1[5]) );
  FA_X1 DP_mult_215_U198 ( .A(DP_mult_215_n456), .B(DP_mult_215_n467), .CI(
        DP_mult_215_n320), .CO(DP_mult_215_n319), .S(DP_sw1_coeff_ret1[6]) );
  FA_X1 DP_mult_215_U197 ( .A(DP_mult_215_n445), .B(DP_mult_215_n455), .CI(
        DP_mult_215_n319), .CO(DP_mult_215_n318), .S(DP_sw1_coeff_ret1[7]) );
  FA_X1 DP_mult_215_U196 ( .A(DP_mult_215_n433), .B(DP_mult_215_n444), .CI(
        DP_mult_215_n318), .CO(DP_mult_215_n317), .S(DP_sw1_coeff_ret1[8]) );
  FA_X1 DP_mult_215_U195 ( .A(DP_mult_215_n423), .B(DP_mult_215_n432), .CI(
        DP_mult_215_n317), .CO(DP_mult_215_n316), .S(DP_sw1_coeff_ret1[9]) );
  FA_X1 DP_mult_215_U194 ( .A(DP_mult_215_n414), .B(DP_mult_215_n422), .CI(
        DP_mult_215_n316), .CO(DP_mult_215_n315), .S(DP_sw1_coeff_ret1[10]) );
  FA_X1 DP_mult_215_U193 ( .A(DP_mult_215_n404), .B(DP_mult_215_n413), .CI(
        DP_mult_215_n315), .CO(DP_mult_215_n314), .S(DP_sw1_coeff_ret1[11]) );
  FA_X1 DP_mult_215_U192 ( .A(DP_mult_215_n397), .B(DP_mult_215_n403), .CI(
        DP_mult_215_n314), .CO(DP_mult_215_n313), .S(DP_sw1_coeff_ret1[12]) );
  FA_X1 DP_mult_215_U191 ( .A(DP_mult_215_n390), .B(DP_mult_215_n396), .CI(
        DP_mult_215_n313), .CO(DP_mult_215_n312), .S(DP_sw1_coeff_ret1[13]) );
  FA_X1 DP_mult_215_U190 ( .A(DP_mult_215_n382), .B(DP_mult_215_n389), .CI(
        DP_mult_215_n312), .CO(DP_mult_215_n311), .S(DP_sw1_coeff_ret1[14]) );
  FA_X1 DP_mult_215_U189 ( .A(DP_mult_215_n376), .B(DP_mult_215_n381), .CI(
        DP_mult_215_n311), .CO(DP_mult_215_n310), .S(DP_sw1_coeff_ret1[15]) );
  FA_X1 DP_mult_215_U188 ( .A(DP_mult_215_n371), .B(DP_mult_215_n375), .CI(
        DP_mult_215_n310), .CO(DP_mult_215_n309), .S(DP_sw1_coeff_ret1[16]) );
  FA_X1 DP_mult_215_U187 ( .A(DP_mult_215_n365), .B(DP_mult_215_n370), .CI(
        DP_mult_215_n309), .CO(DP_mult_215_n308), .S(DP_sw1_coeff_ret1[17]) );
  FA_X1 DP_mult_215_U186 ( .A(DP_mult_215_n362), .B(DP_mult_215_n364), .CI(
        DP_mult_215_n308), .CO(DP_mult_215_n307), .S(DP_sw1_coeff_ret1[18]) );
  FA_X1 DP_mult_215_U185 ( .A(DP_mult_215_n359), .B(DP_mult_215_n361), .CI(
        DP_mult_215_n307), .CO(DP_mult_215_n306), .S(DP_sw1_coeff_ret1[19]) );
  FA_X1 DP_mult_215_U184 ( .A(DP_mult_215_n355), .B(DP_mult_215_n358), .CI(
        DP_mult_215_n306), .CO(DP_mult_215_n305), .S(DP_sw1_coeff_ret1[20]) );
  FA_X1 DP_mult_215_U183 ( .A(DP_mult_215_n353), .B(DP_mult_215_n354), .CI(
        DP_mult_215_n305), .CO(DP_mult_215_n304), .S(DP_sw1_coeff_ret1[21]) );
  FA_X1 DP_mult_215_U182 ( .A(DP_mult_215_n351), .B(DP_mult_215_n352), .CI(
        DP_mult_215_n304), .CO(DP_mult_215_n303), .S(DP_sw1_coeff_ret1[22]) );
  XNOR2_X1 DP_mult_216_U1130 ( .A(DP_b_int_0__2_), .B(DP_mult_216_n975), .ZN(
        DP_mult_216_n1257) );
  INV_X1 DP_mult_216_U1129 ( .A(DP_b_int_0__0_), .ZN(DP_mult_216_n990) );
  XOR2_X1 DP_mult_216_U1128 ( .A(DP_b_int_0__1_), .B(DP_mult_216_n964), .Z(
        DP_mult_216_n1256) );
  INV_X1 DP_mult_216_U1127 ( .A(DP_mult_216_n992), .ZN(DP_mult_216_n1001) );
  INV_X1 DP_mult_216_U1126 ( .A(DP_mult_216_n1256), .ZN(DP_mult_216_n1263) );
  OAI22_X1 DP_mult_216_U1125 ( .A1(DP_mult_216_n1001), .A2(DP_mult_216_n1056), 
        .B1(DP_mult_216_n967), .B2(DP_mult_216_n1056), .ZN(DP_mult_216_n1266)
         );
  XNOR2_X1 DP_mult_216_U1124 ( .A(DP_mult_216_n1266), .B(DP_mult_216_n975), 
        .ZN(DP_mult_216_n1264) );
  NOR2_X1 DP_mult_216_U1123 ( .A1(DP_mult_216_n964), .A2(DP_pipe00[0]), .ZN(
        DP_mult_216_n1265) );
  AOI222_X1 DP_mult_216_U1122 ( .A1(DP_mult_216_n1264), .A2(DP_mult_216_n363), 
        .B1(DP_mult_216_n1265), .B2(DP_mult_216_n1264), .C1(DP_mult_216_n1265), 
        .C2(DP_mult_216_n363), .ZN(DP_mult_216_n1259) );
  INV_X1 DP_mult_216_U1121 ( .A(DP_pipe00[1]), .ZN(DP_mult_216_n1060) );
  XNOR2_X1 DP_mult_216_U1120 ( .A(DP_b_int_0__1_), .B(DP_b_int_0__2_), .ZN(
        DP_mult_216_n1258) );
  INV_X1 DP_mult_216_U1119 ( .A(DP_mult_216_n825), .ZN(DP_mult_216_n1062) );
  OAI222_X1 DP_mult_216_U1118 ( .A1(DP_mult_216_n1060), .A2(DP_mult_216_n1001), 
        .B1(DP_mult_216_n958), .B2(DP_mult_216_n1056), .C1(DP_mult_216_n967), 
        .C2(DP_mult_216_n1062), .ZN(DP_mult_216_n1262) );
  XNOR2_X1 DP_mult_216_U1117 ( .A(DP_mult_216_n1262), .B(DP_mult_216_n974), 
        .ZN(DP_mult_216_n1260) );
  INV_X1 DP_mult_216_U1116 ( .A(DP_mult_216_n361), .ZN(DP_mult_216_n1261) );
  OAI222_X1 DP_mult_216_U1115 ( .A1(DP_mult_216_n1259), .A2(DP_mult_216_n1260), 
        .B1(DP_mult_216_n1259), .B2(DP_mult_216_n1261), .C1(DP_mult_216_n1261), 
        .C2(DP_mult_216_n1260), .ZN(DP_mult_216_n1252) );
  INV_X1 DP_mult_216_U1114 ( .A(DP_mult_216_n824), .ZN(DP_mult_216_n1067) );
  NAND3_X1 DP_mult_216_U1113 ( .A1(DP_mult_216_n1256), .A2(DP_mult_216_n1257), 
        .A3(DP_mult_216_n1258), .ZN(DP_mult_216_n996) );
  OAI22_X1 DP_mult_216_U1112 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1067), 
        .B1(DP_mult_216_n968), .B2(DP_mult_216_n1056), .ZN(DP_mult_216_n1255)
         );
  AOI221_X1 DP_mult_216_U1111 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[2]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[1]), .A(DP_mult_216_n1255), .ZN(
        DP_mult_216_n1254) );
  XNOR2_X1 DP_mult_216_U1110 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1254), 
        .ZN(DP_mult_216_n1253) );
  AOI222_X1 DP_mult_216_U1109 ( .A1(DP_mult_216_n1252), .A2(DP_mult_216_n1253), 
        .B1(DP_mult_216_n1252), .B2(DP_mult_216_n359), .C1(DP_mult_216_n359), 
        .C2(DP_mult_216_n1253), .ZN(DP_mult_216_n1247) );
  INV_X1 DP_mult_216_U1108 ( .A(DP_mult_216_n355), .ZN(DP_mult_216_n1248) );
  INV_X1 DP_mult_216_U1107 ( .A(DP_mult_216_n823), .ZN(DP_mult_216_n1071) );
  OAI22_X1 DP_mult_216_U1106 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1071), 
        .B1(DP_mult_216_n1060), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1251)
         );
  AOI221_X1 DP_mult_216_U1105 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[3]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[2]), .A(DP_mult_216_n1251), .ZN(
        DP_mult_216_n1250) );
  XNOR2_X1 DP_mult_216_U1104 ( .A(DP_mult_216_n975), .B(DP_mult_216_n1250), 
        .ZN(DP_mult_216_n1249) );
  OAI222_X1 DP_mult_216_U1103 ( .A1(DP_mult_216_n1247), .A2(DP_mult_216_n1248), 
        .B1(DP_mult_216_n1247), .B2(DP_mult_216_n1249), .C1(DP_mult_216_n1249), 
        .C2(DP_mult_216_n1248), .ZN(DP_mult_216_n1243) );
  INV_X1 DP_mult_216_U1102 ( .A(DP_mult_216_n822), .ZN(DP_mult_216_n1074) );
  INV_X1 DP_mult_216_U1101 ( .A(DP_pipe00[2]), .ZN(DP_mult_216_n1075) );
  OAI22_X1 DP_mult_216_U1100 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1074), 
        .B1(DP_mult_216_n1075), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1246)
         );
  AOI221_X1 DP_mult_216_U1099 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[4]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[3]), .A(DP_mult_216_n1246), .ZN(
        DP_mult_216_n1245) );
  XNOR2_X1 DP_mult_216_U1098 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1245), 
        .ZN(DP_mult_216_n1244) );
  AOI222_X1 DP_mult_216_U1097 ( .A1(DP_mult_216_n1243), .A2(DP_mult_216_n351), 
        .B1(DP_mult_216_n1243), .B2(DP_mult_216_n1244), .C1(DP_mult_216_n1244), 
        .C2(DP_mult_216_n351), .ZN(DP_mult_216_n1238) );
  INV_X1 DP_mult_216_U1096 ( .A(DP_mult_216_n347), .ZN(DP_mult_216_n1239) );
  INV_X1 DP_mult_216_U1095 ( .A(DP_mult_216_n821), .ZN(DP_mult_216_n1078) );
  INV_X1 DP_mult_216_U1094 ( .A(DP_pipe00[3]), .ZN(DP_mult_216_n1079) );
  OAI22_X1 DP_mult_216_U1093 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1078), 
        .B1(DP_mult_216_n1079), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1242)
         );
  AOI221_X1 DP_mult_216_U1092 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[5]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[4]), .A(DP_mult_216_n1242), .ZN(
        DP_mult_216_n1241) );
  XNOR2_X1 DP_mult_216_U1091 ( .A(DP_mult_216_n975), .B(DP_mult_216_n1241), 
        .ZN(DP_mult_216_n1240) );
  OAI222_X1 DP_mult_216_U1090 ( .A1(DP_mult_216_n1238), .A2(DP_mult_216_n1239), 
        .B1(DP_mult_216_n1238), .B2(DP_mult_216_n1240), .C1(DP_mult_216_n1240), 
        .C2(DP_mult_216_n1239), .ZN(DP_mult_216_n1234) );
  INV_X1 DP_mult_216_U1089 ( .A(DP_mult_216_n820), .ZN(DP_mult_216_n1082) );
  INV_X1 DP_mult_216_U1088 ( .A(DP_pipe00[4]), .ZN(DP_mult_216_n1083) );
  OAI22_X1 DP_mult_216_U1087 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1082), 
        .B1(DP_mult_216_n1083), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1237)
         );
  AOI221_X1 DP_mult_216_U1086 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[6]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[5]), .A(DP_mult_216_n1237), .ZN(
        DP_mult_216_n1236) );
  XNOR2_X1 DP_mult_216_U1085 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1236), 
        .ZN(DP_mult_216_n1235) );
  AOI222_X1 DP_mult_216_U1084 ( .A1(DP_mult_216_n1234), .A2(DP_mult_216_n341), 
        .B1(DP_mult_216_n1234), .B2(DP_mult_216_n1235), .C1(DP_mult_216_n1235), 
        .C2(DP_mult_216_n341), .ZN(DP_mult_216_n1229) );
  INV_X1 DP_mult_216_U1083 ( .A(DP_mult_216_n335), .ZN(DP_mult_216_n1230) );
  INV_X1 DP_mult_216_U1082 ( .A(DP_mult_216_n819), .ZN(DP_mult_216_n1086) );
  INV_X1 DP_mult_216_U1081 ( .A(DP_pipe00[5]), .ZN(DP_mult_216_n1087) );
  OAI22_X1 DP_mult_216_U1080 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1086), 
        .B1(DP_mult_216_n1087), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1233)
         );
  AOI221_X1 DP_mult_216_U1079 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[7]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[6]), .A(DP_mult_216_n1233), .ZN(
        DP_mult_216_n1232) );
  XNOR2_X1 DP_mult_216_U1078 ( .A(DP_mult_216_n975), .B(DP_mult_216_n1232), 
        .ZN(DP_mult_216_n1231) );
  OAI222_X1 DP_mult_216_U1077 ( .A1(DP_mult_216_n1229), .A2(DP_mult_216_n1230), 
        .B1(DP_mult_216_n1229), .B2(DP_mult_216_n1231), .C1(DP_mult_216_n1231), 
        .C2(DP_mult_216_n1230), .ZN(DP_mult_216_n1225) );
  INV_X1 DP_mult_216_U1076 ( .A(DP_mult_216_n818), .ZN(DP_mult_216_n1090) );
  INV_X1 DP_mult_216_U1075 ( .A(DP_pipe00[6]), .ZN(DP_mult_216_n1091) );
  OAI22_X1 DP_mult_216_U1074 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1090), 
        .B1(DP_mult_216_n1091), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1228)
         );
  AOI221_X1 DP_mult_216_U1073 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[8]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[7]), .A(DP_mult_216_n1228), .ZN(
        DP_mult_216_n1227) );
  XNOR2_X1 DP_mult_216_U1072 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1227), 
        .ZN(DP_mult_216_n1226) );
  AOI222_X1 DP_mult_216_U1071 ( .A1(DP_mult_216_n1225), .A2(DP_mult_216_n329), 
        .B1(DP_mult_216_n1225), .B2(DP_mult_216_n1226), .C1(DP_mult_216_n1226), 
        .C2(DP_mult_216_n329), .ZN(DP_mult_216_n1220) );
  INV_X1 DP_mult_216_U1070 ( .A(DP_mult_216_n321), .ZN(DP_mult_216_n1221) );
  INV_X1 DP_mult_216_U1069 ( .A(DP_mult_216_n817), .ZN(DP_mult_216_n1094) );
  INV_X1 DP_mult_216_U1068 ( .A(DP_pipe00[7]), .ZN(DP_mult_216_n1095) );
  OAI22_X1 DP_mult_216_U1067 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1094), 
        .B1(DP_mult_216_n1095), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1224)
         );
  AOI221_X1 DP_mult_216_U1066 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[9]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[8]), .A(DP_mult_216_n1224), .ZN(
        DP_mult_216_n1223) );
  XNOR2_X1 DP_mult_216_U1065 ( .A(DP_mult_216_n975), .B(DP_mult_216_n1223), 
        .ZN(DP_mult_216_n1222) );
  OAI222_X1 DP_mult_216_U1064 ( .A1(DP_mult_216_n1220), .A2(DP_mult_216_n1221), 
        .B1(DP_mult_216_n1220), .B2(DP_mult_216_n1222), .C1(DP_mult_216_n1222), 
        .C2(DP_mult_216_n1221), .ZN(DP_mult_216_n158) );
  XNOR2_X1 DP_mult_216_U1063 ( .A(DP_b_int_0__10_), .B(DP_mult_216_n979), .ZN(
        DP_mult_216_n988) );
  XNOR2_X1 DP_mult_216_U1062 ( .A(DP_mult_216_n980), .B(DP_b_int_0__10_), .ZN(
        DP_mult_216_n1219) );
  NOR2_X1 DP_mult_216_U1061 ( .A1(DP_mult_216_n959), .A2(DP_mult_216_n1219), 
        .ZN(DP_mult_216_n989) );
  AOI22_X1 DP_mult_216_U1060 ( .A1(DP_pipe00[23]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[22]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1218) );
  XOR2_X1 DP_mult_216_U1059 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1218), .Z(
        DP_mult_216_n172) );
  INV_X1 DP_mult_216_U1058 ( .A(DP_mult_216_n177), .ZN(DP_mult_216_n181) );
  AOI22_X1 DP_mult_216_U1057 ( .A1(DP_pipe00[17]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[16]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1217) );
  XOR2_X1 DP_mult_216_U1056 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1217), .Z(
        DP_mult_216_n195) );
  INV_X1 DP_mult_216_U1055 ( .A(DP_mult_216_n195), .ZN(DP_mult_216_n189) );
  OR2_X1 DP_mult_216_U1054 ( .A1(DP_mult_216_n965), .A2(DP_pipe00[23]), .ZN(
        DP_mult_216_n1216) );
  NOR2_X1 DP_mult_216_U1053 ( .A1(DP_mult_216_n1216), .A2(DP_mult_216_n230), 
        .ZN(DP_mult_216_n216) );
  INV_X1 DP_mult_216_U1052 ( .A(DP_mult_216_n216), .ZN(DP_mult_216_n208) );
  XNOR2_X1 DP_mult_216_U1051 ( .A(DP_mult_216_n230), .B(DP_mult_216_n1216), 
        .ZN(DP_mult_216_n223) );
  AOI22_X1 DP_mult_216_U1050 ( .A1(DP_pipe00[22]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[21]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1215) );
  XNOR2_X1 DP_mult_216_U1049 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1215), 
        .ZN(DP_mult_216_n396) );
  AOI22_X1 DP_mult_216_U1048 ( .A1(DP_pipe00[21]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[20]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1214) );
  XNOR2_X1 DP_mult_216_U1047 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1214), 
        .ZN(DP_mult_216_n397) );
  AOI22_X1 DP_mult_216_U1046 ( .A1(DP_pipe00[20]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[19]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1213) );
  XNOR2_X1 DP_mult_216_U1045 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1213), 
        .ZN(DP_mult_216_n398) );
  AOI22_X1 DP_mult_216_U1044 ( .A1(DP_pipe00[19]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[18]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1212) );
  XNOR2_X1 DP_mult_216_U1043 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1212), 
        .ZN(DP_mult_216_n399) );
  AOI22_X1 DP_mult_216_U1042 ( .A1(DP_pipe00[18]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[17]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1211) );
  XNOR2_X1 DP_mult_216_U1041 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1211), 
        .ZN(DP_mult_216_n400) );
  AOI22_X1 DP_mult_216_U1040 ( .A1(DP_pipe00[16]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[15]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1210) );
  XNOR2_X1 DP_mult_216_U1039 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1210), 
        .ZN(DP_mult_216_n401) );
  AOI22_X1 DP_mult_216_U1038 ( .A1(DP_pipe00[15]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[14]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1209) );
  XNOR2_X1 DP_mult_216_U1037 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1209), 
        .ZN(DP_mult_216_n402) );
  AOI22_X1 DP_mult_216_U1036 ( .A1(DP_pipe00[14]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[13]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1208) );
  XNOR2_X1 DP_mult_216_U1035 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1208), 
        .ZN(DP_mult_216_n403) );
  AOI22_X1 DP_mult_216_U1034 ( .A1(DP_pipe00[13]), .A2(DP_mult_216_n960), .B1(
        DP_pipe00[12]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1207) );
  XNOR2_X1 DP_mult_216_U1033 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1207), 
        .ZN(DP_mult_216_n404) );
  AOI22_X1 DP_mult_216_U1032 ( .A1(DP_pipe00[12]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[11]), .B2(DP_mult_216_n963), .ZN(DP_mult_216_n1206) );
  XNOR2_X1 DP_mult_216_U1031 ( .A(DP_mult_216_n981), .B(DP_mult_216_n1206), 
        .ZN(DP_mult_216_n405) );
  AOI22_X1 DP_mult_216_U1030 ( .A1(DP_pipe00[11]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[10]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1205) );
  XNOR2_X1 DP_mult_216_U1029 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1205), 
        .ZN(DP_mult_216_n406) );
  AOI22_X1 DP_mult_216_U1028 ( .A1(DP_pipe00[9]), .A2(DP_mult_216_n962), .B1(
        DP_pipe00[10]), .B2(DP_mult_216_n961), .ZN(DP_mult_216_n1204) );
  XNOR2_X1 DP_mult_216_U1027 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1204), 
        .ZN(DP_mult_216_n407) );
  AOI22_X1 DP_mult_216_U1026 ( .A1(DP_pipe00[9]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[8]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1203) );
  XNOR2_X1 DP_mult_216_U1025 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1203), 
        .ZN(DP_mult_216_n408) );
  AOI22_X1 DP_mult_216_U1024 ( .A1(DP_pipe00[8]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[7]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1202) );
  XNOR2_X1 DP_mult_216_U1023 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1202), 
        .ZN(DP_mult_216_n409) );
  AOI22_X1 DP_mult_216_U1022 ( .A1(DP_pipe00[7]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[6]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1201) );
  XNOR2_X1 DP_mult_216_U1021 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1201), 
        .ZN(DP_mult_216_n410) );
  AOI22_X1 DP_mult_216_U1020 ( .A1(DP_pipe00[6]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[5]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1200) );
  XNOR2_X1 DP_mult_216_U1019 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1200), 
        .ZN(DP_mult_216_n411) );
  AOI22_X1 DP_mult_216_U1018 ( .A1(DP_pipe00[5]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[4]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1199) );
  XNOR2_X1 DP_mult_216_U1017 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1199), 
        .ZN(DP_mult_216_n412) );
  AOI22_X1 DP_mult_216_U1016 ( .A1(DP_pipe00[4]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[3]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1198) );
  XNOR2_X1 DP_mult_216_U1015 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1198), 
        .ZN(DP_mult_216_n413) );
  AOI22_X1 DP_mult_216_U1014 ( .A1(DP_pipe00[3]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[2]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1197) );
  XNOR2_X1 DP_mult_216_U1013 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1197), 
        .ZN(DP_mult_216_n414) );
  AOI22_X1 DP_mult_216_U1012 ( .A1(DP_pipe00[2]), .A2(DP_mult_216_n959), .B1(
        DP_pipe00[1]), .B2(DP_mult_216_n962), .ZN(DP_mult_216_n1196) );
  XNOR2_X1 DP_mult_216_U1011 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1196), 
        .ZN(DP_mult_216_n415) );
  AOI22_X1 DP_mult_216_U1010 ( .A1(DP_pipe00[0]), .A2(DP_mult_216_n962), .B1(
        DP_pipe00[1]), .B2(DP_mult_216_n961), .ZN(DP_mult_216_n1195) );
  XNOR2_X1 DP_mult_216_U1009 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1195), 
        .ZN(DP_mult_216_n416) );
  NAND2_X1 DP_mult_216_U1008 ( .A1(DP_pipe00[0]), .A2(DP_mult_216_n960), .ZN(
        DP_mult_216_n1194) );
  XNOR2_X1 DP_mult_216_U1007 ( .A(DP_mult_216_n980), .B(DP_mult_216_n1194), 
        .ZN(DP_mult_216_n417) );
  XOR2_X1 DP_mult_216_U1006 ( .A(DP_b_int_0__7_), .B(DP_mult_216_n977), .Z(
        DP_mult_216_n1193) );
  INV_X1 DP_mult_216_U1005 ( .A(DP_mult_216_n1193), .ZN(DP_mult_216_n1190) );
  XNOR2_X1 DP_mult_216_U1004 ( .A(DP_b_int_0__8_), .B(DP_mult_216_n979), .ZN(
        DP_mult_216_n1192) );
  INV_X1 DP_mult_216_U1003 ( .A(DP_mult_216_n1135), .ZN(DP_mult_216_n1158) );
  XNOR2_X1 DP_mult_216_U1002 ( .A(DP_b_int_0__7_), .B(DP_b_int_0__8_), .ZN(
        DP_mult_216_n1191) );
  NAND3_X1 DP_mult_216_U1001 ( .A1(DP_mult_216_n1193), .A2(DP_mult_216_n1192), 
        .A3(DP_mult_216_n1191), .ZN(DP_mult_216_n1142) );
  INV_X1 DP_mult_216_U1000 ( .A(DP_mult_216_n1139), .ZN(DP_mult_216_n1134) );
  INV_X1 DP_mult_216_U999 ( .A(DP_mult_216_n1140), .ZN(DP_mult_216_n1137) );
  NAND3_X1 DP_mult_216_U998 ( .A1(DP_mult_216_n973), .A2(DP_mult_216_n1134), 
        .A3(DP_mult_216_n1137), .ZN(DP_mult_216_n1189) );
  AOI22_X1 DP_mult_216_U997 ( .A1(DP_mult_216_n1158), .A2(DP_pipe00[23]), .B1(
        DP_pipe00[23]), .B2(DP_mult_216_n1189), .ZN(DP_mult_216_n1188) );
  XNOR2_X1 DP_mult_216_U996 ( .A(DP_mult_216_n979), .B(DP_mult_216_n1188), 
        .ZN(DP_mult_216_n418) );
  INV_X1 DP_mult_216_U995 ( .A(DP_pipe00[22]), .ZN(DP_mult_216_n1050) );
  INV_X1 DP_mult_216_U994 ( .A(DP_mult_216_n802), .ZN(DP_mult_216_n1051) );
  OAI21_X1 DP_mult_216_U993 ( .B1(DP_mult_216_n1139), .B2(DP_mult_216_n1140), 
        .A(DP_pipe00[23]), .ZN(DP_mult_216_n1187) );
  OAI221_X1 DP_mult_216_U992 ( .B1(DP_mult_216_n1050), .B2(DP_mult_216_n973), 
        .C1(DP_mult_216_n1051), .C2(DP_mult_216_n1135), .A(DP_mult_216_n1187), 
        .ZN(DP_mult_216_n1186) );
  XNOR2_X1 DP_mult_216_U991 ( .A(DP_mult_216_n1186), .B(DP_mult_216_n979), 
        .ZN(DP_mult_216_n419) );
  INV_X1 DP_mult_216_U990 ( .A(DP_mult_216_n803), .ZN(DP_mult_216_n1047) );
  INV_X1 DP_mult_216_U989 ( .A(DP_pipe00[21]), .ZN(DP_mult_216_n1048) );
  OAI22_X1 DP_mult_216_U988 ( .A1(DP_mult_216_n1047), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1048), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1185)
         );
  AOI221_X1 DP_mult_216_U987 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[23]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[22]), .A(DP_mult_216_n1185), 
        .ZN(DP_mult_216_n1184) );
  XNOR2_X1 DP_mult_216_U986 ( .A(DP_b_int_0__9_), .B(DP_mult_216_n1184), .ZN(
        DP_mult_216_n420) );
  INV_X1 DP_mult_216_U985 ( .A(DP_mult_216_n804), .ZN(DP_mult_216_n1043) );
  INV_X1 DP_mult_216_U984 ( .A(DP_pipe00[20]), .ZN(DP_mult_216_n1044) );
  OAI22_X1 DP_mult_216_U983 ( .A1(DP_mult_216_n1043), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1044), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1183)
         );
  AOI221_X1 DP_mult_216_U982 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[22]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[21]), .A(DP_mult_216_n1183), 
        .ZN(DP_mult_216_n1182) );
  XNOR2_X1 DP_mult_216_U981 ( .A(DP_b_int_0__9_), .B(DP_mult_216_n1182), .ZN(
        DP_mult_216_n421) );
  INV_X1 DP_mult_216_U980 ( .A(DP_mult_216_n805), .ZN(DP_mult_216_n1039) );
  INV_X1 DP_mult_216_U979 ( .A(DP_pipe00[19]), .ZN(DP_mult_216_n1040) );
  OAI22_X1 DP_mult_216_U978 ( .A1(DP_mult_216_n1039), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1040), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1181)
         );
  AOI221_X1 DP_mult_216_U977 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[21]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[20]), .A(DP_mult_216_n1181), 
        .ZN(DP_mult_216_n1180) );
  XNOR2_X1 DP_mult_216_U976 ( .A(DP_b_int_0__9_), .B(DP_mult_216_n1180), .ZN(
        DP_mult_216_n422) );
  INV_X1 DP_mult_216_U975 ( .A(DP_mult_216_n806), .ZN(DP_mult_216_n1035) );
  INV_X1 DP_mult_216_U974 ( .A(DP_pipe00[18]), .ZN(DP_mult_216_n1036) );
  OAI22_X1 DP_mult_216_U973 ( .A1(DP_mult_216_n1035), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1036), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1179)
         );
  AOI221_X1 DP_mult_216_U972 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[20]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[19]), .A(DP_mult_216_n1179), 
        .ZN(DP_mult_216_n1178) );
  XNOR2_X1 DP_mult_216_U971 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1178), 
        .ZN(DP_mult_216_n423) );
  INV_X1 DP_mult_216_U970 ( .A(DP_pipe00[17]), .ZN(DP_mult_216_n1032) );
  OAI22_X1 DP_mult_216_U969 ( .A1(DP_mult_216_n1040), .A2(DP_mult_216_n1134), 
        .B1(DP_mult_216_n1032), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1177)
         );
  AOI221_X1 DP_mult_216_U968 ( .B1(DP_mult_216_n1140), .B2(DP_pipe00[18]), 
        .C1(DP_mult_216_n1158), .C2(DP_mult_216_n807), .A(DP_mult_216_n1177), 
        .ZN(DP_mult_216_n1176) );
  XNOR2_X1 DP_mult_216_U967 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1176), 
        .ZN(DP_mult_216_n424) );
  INV_X1 DP_mult_216_U966 ( .A(DP_pipe00[16]), .ZN(DP_mult_216_n1028) );
  OAI22_X1 DP_mult_216_U965 ( .A1(DP_mult_216_n1028), .A2(DP_mult_216_n973), 
        .B1(DP_mult_216_n1032), .B2(DP_mult_216_n1137), .ZN(DP_mult_216_n1175)
         );
  AOI221_X1 DP_mult_216_U964 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[18]), 
        .C1(DP_mult_216_n1158), .C2(DP_mult_216_n808), .A(DP_mult_216_n1175), 
        .ZN(DP_mult_216_n1174) );
  XNOR2_X1 DP_mult_216_U963 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1174), 
        .ZN(DP_mult_216_n425) );
  INV_X1 DP_mult_216_U962 ( .A(DP_mult_216_n809), .ZN(DP_mult_216_n1023) );
  INV_X1 DP_mult_216_U961 ( .A(DP_pipe00[15]), .ZN(DP_mult_216_n1024) );
  OAI22_X1 DP_mult_216_U960 ( .A1(DP_mult_216_n1023), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1024), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1173)
         );
  AOI221_X1 DP_mult_216_U959 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[17]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[16]), .A(DP_mult_216_n1173), 
        .ZN(DP_mult_216_n1172) );
  XNOR2_X1 DP_mult_216_U958 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1172), 
        .ZN(DP_mult_216_n426) );
  INV_X1 DP_mult_216_U957 ( .A(DP_mult_216_n810), .ZN(DP_mult_216_n1019) );
  INV_X1 DP_mult_216_U956 ( .A(DP_pipe00[14]), .ZN(DP_mult_216_n1020) );
  OAI22_X1 DP_mult_216_U955 ( .A1(DP_mult_216_n1019), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1020), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1171)
         );
  AOI221_X1 DP_mult_216_U954 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[16]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[15]), .A(DP_mult_216_n1171), 
        .ZN(DP_mult_216_n1170) );
  XNOR2_X1 DP_mult_216_U953 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1170), 
        .ZN(DP_mult_216_n427) );
  INV_X1 DP_mult_216_U952 ( .A(DP_mult_216_n811), .ZN(DP_mult_216_n1015) );
  INV_X1 DP_mult_216_U951 ( .A(DP_pipe00[13]), .ZN(DP_mult_216_n1016) );
  OAI22_X1 DP_mult_216_U950 ( .A1(DP_mult_216_n1015), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1016), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1169)
         );
  AOI221_X1 DP_mult_216_U949 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[15]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[14]), .A(DP_mult_216_n1169), 
        .ZN(DP_mult_216_n1168) );
  XNOR2_X1 DP_mult_216_U948 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1168), 
        .ZN(DP_mult_216_n428) );
  INV_X1 DP_mult_216_U947 ( .A(DP_mult_216_n812), .ZN(DP_mult_216_n1011) );
  INV_X1 DP_mult_216_U946 ( .A(DP_pipe00[12]), .ZN(DP_mult_216_n1012) );
  OAI22_X1 DP_mult_216_U945 ( .A1(DP_mult_216_n1011), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1012), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1167)
         );
  AOI221_X1 DP_mult_216_U944 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[14]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[13]), .A(DP_mult_216_n1167), 
        .ZN(DP_mult_216_n1166) );
  XNOR2_X1 DP_mult_216_U943 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1166), 
        .ZN(DP_mult_216_n429) );
  INV_X1 DP_mult_216_U942 ( .A(DP_mult_216_n813), .ZN(DP_mult_216_n1008) );
  INV_X1 DP_mult_216_U941 ( .A(DP_pipe00[11]), .ZN(DP_mult_216_n1000) );
  OAI22_X1 DP_mult_216_U940 ( .A1(DP_mult_216_n1008), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1000), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1165)
         );
  AOI221_X1 DP_mult_216_U939 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[13]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[12]), .A(DP_mult_216_n1165), 
        .ZN(DP_mult_216_n1164) );
  XNOR2_X1 DP_mult_216_U938 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1164), 
        .ZN(DP_mult_216_n430) );
  INV_X1 DP_mult_216_U937 ( .A(DP_mult_216_n814), .ZN(DP_mult_216_n1004) );
  INV_X1 DP_mult_216_U936 ( .A(DP_pipe00[10]), .ZN(DP_mult_216_n1005) );
  OAI22_X1 DP_mult_216_U935 ( .A1(DP_mult_216_n1004), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1005), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1163)
         );
  AOI221_X1 DP_mult_216_U934 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[12]), 
        .C1(DP_mult_216_n1140), .C2(DP_pipe00[11]), .A(DP_mult_216_n1163), 
        .ZN(DP_mult_216_n1162) );
  XNOR2_X1 DP_mult_216_U933 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1162), 
        .ZN(DP_mult_216_n431) );
  INV_X1 DP_mult_216_U932 ( .A(DP_pipe00[9]), .ZN(DP_mult_216_n999) );
  OAI22_X1 DP_mult_216_U931 ( .A1(DP_mult_216_n1000), .A2(DP_mult_216_n1134), 
        .B1(DP_mult_216_n999), .B2(DP_mult_216_n973), .ZN(DP_mult_216_n1161)
         );
  AOI221_X1 DP_mult_216_U930 ( .B1(DP_mult_216_n1140), .B2(DP_pipe00[10]), 
        .C1(DP_mult_216_n1158), .C2(DP_mult_216_n815), .A(DP_mult_216_n1161), 
        .ZN(DP_mult_216_n1160) );
  XNOR2_X1 DP_mult_216_U929 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1160), 
        .ZN(DP_mult_216_n432) );
  INV_X1 DP_mult_216_U928 ( .A(DP_pipe00[8]), .ZN(DP_mult_216_n995) );
  OAI22_X1 DP_mult_216_U927 ( .A1(DP_mult_216_n995), .A2(DP_mult_216_n973), 
        .B1(DP_mult_216_n999), .B2(DP_mult_216_n1137), .ZN(DP_mult_216_n1159)
         );
  AOI221_X1 DP_mult_216_U926 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[10]), 
        .C1(DP_mult_216_n1158), .C2(DP_mult_216_n816), .A(DP_mult_216_n1159), 
        .ZN(DP_mult_216_n1157) );
  XNOR2_X1 DP_mult_216_U925 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1157), 
        .ZN(DP_mult_216_n433) );
  OAI22_X1 DP_mult_216_U924 ( .A1(DP_mult_216_n1094), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1095), .B2(DP_mult_216_n973), .ZN(DP_mult_216_n1156)
         );
  AOI221_X1 DP_mult_216_U923 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[9]), .C1(
        DP_mult_216_n1140), .C2(DP_pipe00[8]), .A(DP_mult_216_n1156), .ZN(
        DP_mult_216_n1155) );
  XNOR2_X1 DP_mult_216_U922 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1155), 
        .ZN(DP_mult_216_n434) );
  OAI22_X1 DP_mult_216_U921 ( .A1(DP_mult_216_n1090), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1091), .B2(DP_mult_216_n973), .ZN(DP_mult_216_n1154)
         );
  AOI221_X1 DP_mult_216_U920 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[8]), .C1(
        DP_mult_216_n1140), .C2(DP_pipe00[7]), .A(DP_mult_216_n1154), .ZN(
        DP_mult_216_n1153) );
  XNOR2_X1 DP_mult_216_U919 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1153), 
        .ZN(DP_mult_216_n435) );
  OAI22_X1 DP_mult_216_U918 ( .A1(DP_mult_216_n1086), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1087), .B2(DP_mult_216_n973), .ZN(DP_mult_216_n1152)
         );
  AOI221_X1 DP_mult_216_U917 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[7]), .C1(
        DP_mult_216_n1140), .C2(DP_pipe00[6]), .A(DP_mult_216_n1152), .ZN(
        DP_mult_216_n1151) );
  XNOR2_X1 DP_mult_216_U916 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1151), 
        .ZN(DP_mult_216_n436) );
  OAI22_X1 DP_mult_216_U915 ( .A1(DP_mult_216_n1082), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1083), .B2(DP_mult_216_n973), .ZN(DP_mult_216_n1150)
         );
  AOI221_X1 DP_mult_216_U914 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[6]), .C1(
        DP_mult_216_n1140), .C2(DP_pipe00[5]), .A(DP_mult_216_n1150), .ZN(
        DP_mult_216_n1149) );
  XNOR2_X1 DP_mult_216_U913 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1149), 
        .ZN(DP_mult_216_n437) );
  OAI22_X1 DP_mult_216_U912 ( .A1(DP_mult_216_n1078), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1079), .B2(DP_mult_216_n973), .ZN(DP_mult_216_n1148)
         );
  AOI221_X1 DP_mult_216_U911 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[5]), .C1(
        DP_mult_216_n1140), .C2(DP_pipe00[4]), .A(DP_mult_216_n1148), .ZN(
        DP_mult_216_n1147) );
  XNOR2_X1 DP_mult_216_U910 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1147), 
        .ZN(DP_mult_216_n438) );
  OAI22_X1 DP_mult_216_U909 ( .A1(DP_mult_216_n1074), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1075), .B2(DP_mult_216_n973), .ZN(DP_mult_216_n1146)
         );
  AOI221_X1 DP_mult_216_U908 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[4]), .C1(
        DP_mult_216_n1140), .C2(DP_pipe00[3]), .A(DP_mult_216_n1146), .ZN(
        DP_mult_216_n1145) );
  XNOR2_X1 DP_mult_216_U907 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1145), 
        .ZN(DP_mult_216_n439) );
  OAI22_X1 DP_mult_216_U906 ( .A1(DP_mult_216_n1071), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1060), .B2(DP_mult_216_n973), .ZN(DP_mult_216_n1144)
         );
  AOI221_X1 DP_mult_216_U905 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[3]), .C1(
        DP_mult_216_n1140), .C2(DP_pipe00[2]), .A(DP_mult_216_n1144), .ZN(
        DP_mult_216_n1143) );
  XNOR2_X1 DP_mult_216_U904 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1143), 
        .ZN(DP_mult_216_n440) );
  OAI22_X1 DP_mult_216_U903 ( .A1(DP_mult_216_n1067), .A2(DP_mult_216_n1135), 
        .B1(DP_mult_216_n1056), .B2(DP_mult_216_n972), .ZN(DP_mult_216_n1141)
         );
  AOI221_X1 DP_mult_216_U902 ( .B1(DP_mult_216_n1139), .B2(DP_pipe00[2]), .C1(
        DP_mult_216_n1140), .C2(DP_pipe00[1]), .A(DP_mult_216_n1141), .ZN(
        DP_mult_216_n1138) );
  XNOR2_X1 DP_mult_216_U901 ( .A(DP_mult_216_n978), .B(DP_mult_216_n1138), 
        .ZN(DP_mult_216_n441) );
  OAI222_X1 DP_mult_216_U900 ( .A1(DP_mult_216_n1060), .A2(DP_mult_216_n1134), 
        .B1(DP_mult_216_n1056), .B2(DP_mult_216_n1137), .C1(DP_mult_216_n1062), 
        .C2(DP_mult_216_n1135), .ZN(DP_mult_216_n1136) );
  XNOR2_X1 DP_mult_216_U899 ( .A(DP_mult_216_n1136), .B(DP_mult_216_n979), 
        .ZN(DP_mult_216_n442) );
  OAI22_X1 DP_mult_216_U898 ( .A1(DP_mult_216_n1056), .A2(DP_mult_216_n1134), 
        .B1(DP_mult_216_n1056), .B2(DP_mult_216_n1135), .ZN(DP_mult_216_n1133)
         );
  XNOR2_X1 DP_mult_216_U897 ( .A(DP_mult_216_n1133), .B(DP_mult_216_n979), 
        .ZN(DP_mult_216_n443) );
  XOR2_X1 DP_mult_216_U896 ( .A(DP_b_int_0__4_), .B(DP_mult_216_n975), .Z(
        DP_mult_216_n1132) );
  INV_X1 DP_mult_216_U895 ( .A(DP_mult_216_n1132), .ZN(DP_mult_216_n1129) );
  XNOR2_X1 DP_mult_216_U894 ( .A(DP_b_int_0__5_), .B(DP_mult_216_n977), .ZN(
        DP_mult_216_n1131) );
  INV_X1 DP_mult_216_U893 ( .A(DP_mult_216_n1058), .ZN(DP_mult_216_n1097) );
  XNOR2_X1 DP_mult_216_U892 ( .A(DP_b_int_0__4_), .B(DP_b_int_0__5_), .ZN(
        DP_mult_216_n1130) );
  NAND3_X1 DP_mult_216_U891 ( .A1(DP_mult_216_n1132), .A2(DP_mult_216_n1131), 
        .A3(DP_mult_216_n1130), .ZN(DP_mult_216_n1068) );
  INV_X1 DP_mult_216_U890 ( .A(DP_mult_216_n1064), .ZN(DP_mult_216_n1057) );
  INV_X1 DP_mult_216_U889 ( .A(DP_mult_216_n1065), .ZN(DP_mult_216_n1061) );
  NAND3_X1 DP_mult_216_U888 ( .A1(DP_mult_216_n971), .A2(DP_mult_216_n1057), 
        .A3(DP_mult_216_n1061), .ZN(DP_mult_216_n1128) );
  AOI22_X1 DP_mult_216_U887 ( .A1(DP_mult_216_n1097), .A2(DP_pipe00[23]), .B1(
        DP_pipe00[23]), .B2(DP_mult_216_n1128), .ZN(DP_mult_216_n1127) );
  XNOR2_X1 DP_mult_216_U886 ( .A(DP_mult_216_n977), .B(DP_mult_216_n1127), 
        .ZN(DP_mult_216_n444) );
  OAI21_X1 DP_mult_216_U885 ( .B1(DP_mult_216_n1064), .B2(DP_mult_216_n1065), 
        .A(DP_pipe00[23]), .ZN(DP_mult_216_n1126) );
  OAI221_X1 DP_mult_216_U884 ( .B1(DP_mult_216_n1050), .B2(DP_mult_216_n971), 
        .C1(DP_mult_216_n1051), .C2(DP_mult_216_n1058), .A(DP_mult_216_n1126), 
        .ZN(DP_mult_216_n1125) );
  XNOR2_X1 DP_mult_216_U883 ( .A(DP_mult_216_n1125), .B(DP_mult_216_n977), 
        .ZN(DP_mult_216_n445) );
  OAI22_X1 DP_mult_216_U882 ( .A1(DP_mult_216_n1047), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1048), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1124)
         );
  AOI221_X1 DP_mult_216_U881 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[23]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[22]), .A(DP_mult_216_n1124), 
        .ZN(DP_mult_216_n1123) );
  XNOR2_X1 DP_mult_216_U880 ( .A(DP_b_int_0__6_), .B(DP_mult_216_n1123), .ZN(
        DP_mult_216_n446) );
  OAI22_X1 DP_mult_216_U879 ( .A1(DP_mult_216_n1043), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1044), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1122)
         );
  AOI221_X1 DP_mult_216_U878 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[22]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[21]), .A(DP_mult_216_n1122), 
        .ZN(DP_mult_216_n1121) );
  XNOR2_X1 DP_mult_216_U877 ( .A(DP_b_int_0__6_), .B(DP_mult_216_n1121), .ZN(
        DP_mult_216_n447) );
  OAI22_X1 DP_mult_216_U876 ( .A1(DP_mult_216_n1039), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1040), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1120)
         );
  AOI221_X1 DP_mult_216_U875 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[21]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[20]), .A(DP_mult_216_n1120), 
        .ZN(DP_mult_216_n1119) );
  XNOR2_X1 DP_mult_216_U874 ( .A(DP_b_int_0__6_), .B(DP_mult_216_n1119), .ZN(
        DP_mult_216_n448) );
  OAI22_X1 DP_mult_216_U873 ( .A1(DP_mult_216_n1035), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1036), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1118)
         );
  AOI221_X1 DP_mult_216_U872 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[20]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[19]), .A(DP_mult_216_n1118), 
        .ZN(DP_mult_216_n1117) );
  XNOR2_X1 DP_mult_216_U871 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1117), 
        .ZN(DP_mult_216_n449) );
  OAI22_X1 DP_mult_216_U870 ( .A1(DP_mult_216_n1040), .A2(DP_mult_216_n1057), 
        .B1(DP_mult_216_n1032), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1116)
         );
  AOI221_X1 DP_mult_216_U869 ( .B1(DP_mult_216_n1065), .B2(DP_pipe00[18]), 
        .C1(DP_mult_216_n1097), .C2(DP_mult_216_n807), .A(DP_mult_216_n1116), 
        .ZN(DP_mult_216_n1115) );
  XNOR2_X1 DP_mult_216_U868 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1115), 
        .ZN(DP_mult_216_n450) );
  OAI22_X1 DP_mult_216_U867 ( .A1(DP_mult_216_n1028), .A2(DP_mult_216_n971), 
        .B1(DP_mult_216_n1032), .B2(DP_mult_216_n1061), .ZN(DP_mult_216_n1114)
         );
  AOI221_X1 DP_mult_216_U866 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[18]), 
        .C1(DP_mult_216_n1097), .C2(DP_mult_216_n808), .A(DP_mult_216_n1114), 
        .ZN(DP_mult_216_n1113) );
  XNOR2_X1 DP_mult_216_U865 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1113), 
        .ZN(DP_mult_216_n451) );
  OAI22_X1 DP_mult_216_U864 ( .A1(DP_mult_216_n1023), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1024), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1112)
         );
  AOI221_X1 DP_mult_216_U863 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[17]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[16]), .A(DP_mult_216_n1112), 
        .ZN(DP_mult_216_n1111) );
  XNOR2_X1 DP_mult_216_U862 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1111), 
        .ZN(DP_mult_216_n452) );
  OAI22_X1 DP_mult_216_U861 ( .A1(DP_mult_216_n1019), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1020), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1110)
         );
  AOI221_X1 DP_mult_216_U860 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[16]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[15]), .A(DP_mult_216_n1110), 
        .ZN(DP_mult_216_n1109) );
  XNOR2_X1 DP_mult_216_U859 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1109), 
        .ZN(DP_mult_216_n453) );
  OAI22_X1 DP_mult_216_U858 ( .A1(DP_mult_216_n1015), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1016), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1108)
         );
  AOI221_X1 DP_mult_216_U857 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[15]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[14]), .A(DP_mult_216_n1108), 
        .ZN(DP_mult_216_n1107) );
  XNOR2_X1 DP_mult_216_U856 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1107), 
        .ZN(DP_mult_216_n454) );
  OAI22_X1 DP_mult_216_U855 ( .A1(DP_mult_216_n1011), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1012), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1106)
         );
  AOI221_X1 DP_mult_216_U854 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[14]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[13]), .A(DP_mult_216_n1106), 
        .ZN(DP_mult_216_n1105) );
  XNOR2_X1 DP_mult_216_U853 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1105), 
        .ZN(DP_mult_216_n455) );
  OAI22_X1 DP_mult_216_U852 ( .A1(DP_mult_216_n1008), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1000), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1104)
         );
  AOI221_X1 DP_mult_216_U851 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[13]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[12]), .A(DP_mult_216_n1104), 
        .ZN(DP_mult_216_n1103) );
  XNOR2_X1 DP_mult_216_U850 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1103), 
        .ZN(DP_mult_216_n456) );
  OAI22_X1 DP_mult_216_U849 ( .A1(DP_mult_216_n1004), .A2(DP_mult_216_n1058), 
        .B1(DP_mult_216_n1005), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1102)
         );
  AOI221_X1 DP_mult_216_U848 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[12]), 
        .C1(DP_mult_216_n1065), .C2(DP_pipe00[11]), .A(DP_mult_216_n1102), 
        .ZN(DP_mult_216_n1101) );
  XNOR2_X1 DP_mult_216_U847 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1101), 
        .ZN(DP_mult_216_n457) );
  OAI22_X1 DP_mult_216_U846 ( .A1(DP_mult_216_n1000), .A2(DP_mult_216_n1057), 
        .B1(DP_mult_216_n999), .B2(DP_mult_216_n971), .ZN(DP_mult_216_n1100)
         );
  AOI221_X1 DP_mult_216_U845 ( .B1(DP_mult_216_n1065), .B2(DP_pipe00[10]), 
        .C1(DP_mult_216_n1097), .C2(DP_mult_216_n815), .A(DP_mult_216_n1100), 
        .ZN(DP_mult_216_n1099) );
  XNOR2_X1 DP_mult_216_U844 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1099), 
        .ZN(DP_mult_216_n458) );
  OAI22_X1 DP_mult_216_U843 ( .A1(DP_mult_216_n995), .A2(DP_mult_216_n971), 
        .B1(DP_mult_216_n999), .B2(DP_mult_216_n1061), .ZN(DP_mult_216_n1098)
         );
  AOI221_X1 DP_mult_216_U842 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[10]), 
        .C1(DP_mult_216_n1097), .C2(DP_mult_216_n816), .A(DP_mult_216_n1098), 
        .ZN(DP_mult_216_n1096) );
  XNOR2_X1 DP_mult_216_U841 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1096), 
        .ZN(DP_mult_216_n459) );
  OAI22_X1 DP_mult_216_U840 ( .A1(DP_mult_216_n1058), .A2(DP_mult_216_n1094), 
        .B1(DP_mult_216_n1095), .B2(DP_mult_216_n971), .ZN(DP_mult_216_n1093)
         );
  AOI221_X1 DP_mult_216_U839 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[9]), .C1(
        DP_mult_216_n1065), .C2(DP_pipe00[8]), .A(DP_mult_216_n1093), .ZN(
        DP_mult_216_n1092) );
  XNOR2_X1 DP_mult_216_U838 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1092), 
        .ZN(DP_mult_216_n460) );
  OAI22_X1 DP_mult_216_U837 ( .A1(DP_mult_216_n1058), .A2(DP_mult_216_n1090), 
        .B1(DP_mult_216_n1091), .B2(DP_mult_216_n971), .ZN(DP_mult_216_n1089)
         );
  AOI221_X1 DP_mult_216_U836 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[8]), .C1(
        DP_mult_216_n1065), .C2(DP_pipe00[7]), .A(DP_mult_216_n1089), .ZN(
        DP_mult_216_n1088) );
  XNOR2_X1 DP_mult_216_U835 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1088), 
        .ZN(DP_mult_216_n461) );
  OAI22_X1 DP_mult_216_U834 ( .A1(DP_mult_216_n1058), .A2(DP_mult_216_n1086), 
        .B1(DP_mult_216_n1087), .B2(DP_mult_216_n971), .ZN(DP_mult_216_n1085)
         );
  AOI221_X1 DP_mult_216_U833 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[7]), .C1(
        DP_mult_216_n1065), .C2(DP_pipe00[6]), .A(DP_mult_216_n1085), .ZN(
        DP_mult_216_n1084) );
  XNOR2_X1 DP_mult_216_U832 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1084), 
        .ZN(DP_mult_216_n462) );
  OAI22_X1 DP_mult_216_U831 ( .A1(DP_mult_216_n1058), .A2(DP_mult_216_n1082), 
        .B1(DP_mult_216_n1083), .B2(DP_mult_216_n971), .ZN(DP_mult_216_n1081)
         );
  AOI221_X1 DP_mult_216_U830 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[6]), .C1(
        DP_mult_216_n1065), .C2(DP_pipe00[5]), .A(DP_mult_216_n1081), .ZN(
        DP_mult_216_n1080) );
  XNOR2_X1 DP_mult_216_U829 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1080), 
        .ZN(DP_mult_216_n463) );
  OAI22_X1 DP_mult_216_U828 ( .A1(DP_mult_216_n1058), .A2(DP_mult_216_n1078), 
        .B1(DP_mult_216_n1079), .B2(DP_mult_216_n971), .ZN(DP_mult_216_n1077)
         );
  AOI221_X1 DP_mult_216_U827 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[5]), .C1(
        DP_mult_216_n1065), .C2(DP_pipe00[4]), .A(DP_mult_216_n1077), .ZN(
        DP_mult_216_n1076) );
  XNOR2_X1 DP_mult_216_U826 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1076), 
        .ZN(DP_mult_216_n464) );
  OAI22_X1 DP_mult_216_U825 ( .A1(DP_mult_216_n1058), .A2(DP_mult_216_n1074), 
        .B1(DP_mult_216_n1075), .B2(DP_mult_216_n971), .ZN(DP_mult_216_n1073)
         );
  AOI221_X1 DP_mult_216_U824 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[4]), .C1(
        DP_mult_216_n1065), .C2(DP_pipe00[3]), .A(DP_mult_216_n1073), .ZN(
        DP_mult_216_n1072) );
  XNOR2_X1 DP_mult_216_U823 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1072), 
        .ZN(DP_mult_216_n465) );
  OAI22_X1 DP_mult_216_U822 ( .A1(DP_mult_216_n1058), .A2(DP_mult_216_n1071), 
        .B1(DP_mult_216_n1060), .B2(DP_mult_216_n971), .ZN(DP_mult_216_n1070)
         );
  AOI221_X1 DP_mult_216_U821 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[3]), .C1(
        DP_mult_216_n1065), .C2(DP_pipe00[2]), .A(DP_mult_216_n1070), .ZN(
        DP_mult_216_n1069) );
  XNOR2_X1 DP_mult_216_U820 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1069), 
        .ZN(DP_mult_216_n466) );
  OAI22_X1 DP_mult_216_U819 ( .A1(DP_mult_216_n1058), .A2(DP_mult_216_n1067), 
        .B1(DP_mult_216_n1056), .B2(DP_mult_216_n970), .ZN(DP_mult_216_n1066)
         );
  AOI221_X1 DP_mult_216_U818 ( .B1(DP_mult_216_n1064), .B2(DP_pipe00[2]), .C1(
        DP_mult_216_n1065), .C2(DP_pipe00[1]), .A(DP_mult_216_n1066), .ZN(
        DP_mult_216_n1063) );
  XNOR2_X1 DP_mult_216_U817 ( .A(DP_mult_216_n976), .B(DP_mult_216_n1063), 
        .ZN(DP_mult_216_n467) );
  OAI222_X1 DP_mult_216_U816 ( .A1(DP_mult_216_n1060), .A2(DP_mult_216_n1057), 
        .B1(DP_mult_216_n1056), .B2(DP_mult_216_n1061), .C1(DP_mult_216_n1058), 
        .C2(DP_mult_216_n1062), .ZN(DP_mult_216_n1059) );
  XNOR2_X1 DP_mult_216_U815 ( .A(DP_mult_216_n1059), .B(DP_mult_216_n977), 
        .ZN(DP_mult_216_n468) );
  OAI22_X1 DP_mult_216_U814 ( .A1(DP_mult_216_n1056), .A2(DP_mult_216_n1057), 
        .B1(DP_mult_216_n1058), .B2(DP_mult_216_n1056), .ZN(DP_mult_216_n1055)
         );
  XNOR2_X1 DP_mult_216_U813 ( .A(DP_mult_216_n1055), .B(DP_mult_216_n977), 
        .ZN(DP_mult_216_n469) );
  NAND3_X1 DP_mult_216_U812 ( .A1(DP_mult_216_n969), .A2(DP_mult_216_n1001), 
        .A3(DP_mult_216_n958), .ZN(DP_mult_216_n1054) );
  AOI22_X1 DP_mult_216_U811 ( .A1(DP_mult_216_n957), .A2(DP_pipe00[23]), .B1(
        DP_pipe00[23]), .B2(DP_mult_216_n1054), .ZN(DP_mult_216_n1053) );
  XNOR2_X1 DP_mult_216_U810 ( .A(DP_mult_216_n975), .B(DP_mult_216_n1053), 
        .ZN(DP_mult_216_n470) );
  OAI21_X1 DP_mult_216_U809 ( .B1(DP_mult_216_n992), .B2(DP_mult_216_n966), 
        .A(DP_pipe00[23]), .ZN(DP_mult_216_n1052) );
  OAI221_X1 DP_mult_216_U808 ( .B1(DP_mult_216_n1050), .B2(DP_mult_216_n969), 
        .C1(DP_mult_216_n967), .C2(DP_mult_216_n1051), .A(DP_mult_216_n1052), 
        .ZN(DP_mult_216_n1049) );
  XNOR2_X1 DP_mult_216_U807 ( .A(DP_mult_216_n1049), .B(DP_mult_216_n975), 
        .ZN(DP_mult_216_n471) );
  OAI22_X1 DP_mult_216_U806 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1047), 
        .B1(DP_mult_216_n1048), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1046)
         );
  AOI221_X1 DP_mult_216_U805 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[23]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[22]), .A(DP_mult_216_n1046), .ZN(
        DP_mult_216_n1045) );
  XNOR2_X1 DP_mult_216_U804 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1045), 
        .ZN(DP_mult_216_n472) );
  OAI22_X1 DP_mult_216_U803 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1043), 
        .B1(DP_mult_216_n1044), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1042)
         );
  AOI221_X1 DP_mult_216_U802 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[22]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[21]), .A(DP_mult_216_n1042), .ZN(
        DP_mult_216_n1041) );
  XNOR2_X1 DP_mult_216_U801 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1041), 
        .ZN(DP_mult_216_n473) );
  OAI22_X1 DP_mult_216_U800 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1039), 
        .B1(DP_mult_216_n1040), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n1038)
         );
  AOI221_X1 DP_mult_216_U799 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[21]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[20]), .A(DP_mult_216_n1038), .ZN(
        DP_mult_216_n1037) );
  XNOR2_X1 DP_mult_216_U798 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1037), 
        .ZN(DP_mult_216_n474) );
  OAI22_X1 DP_mult_216_U797 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1035), 
        .B1(DP_mult_216_n1036), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1034)
         );
  AOI221_X1 DP_mult_216_U796 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[20]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[19]), .A(DP_mult_216_n1034), .ZN(
        DP_mult_216_n1033) );
  XNOR2_X1 DP_mult_216_U795 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1033), 
        .ZN(DP_mult_216_n475) );
  INV_X1 DP_mult_216_U794 ( .A(DP_mult_216_n807), .ZN(DP_mult_216_n1031) );
  OAI22_X1 DP_mult_216_U793 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1031), 
        .B1(DP_mult_216_n1032), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1030)
         );
  AOI221_X1 DP_mult_216_U792 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[19]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[18]), .A(DP_mult_216_n1030), .ZN(
        DP_mult_216_n1029) );
  XNOR2_X1 DP_mult_216_U791 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1029), 
        .ZN(DP_mult_216_n476) );
  INV_X1 DP_mult_216_U790 ( .A(DP_mult_216_n808), .ZN(DP_mult_216_n1027) );
  OAI22_X1 DP_mult_216_U789 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1027), 
        .B1(DP_mult_216_n1028), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1026)
         );
  AOI221_X1 DP_mult_216_U788 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[18]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[17]), .A(DP_mult_216_n1026), .ZN(
        DP_mult_216_n1025) );
  XNOR2_X1 DP_mult_216_U787 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1025), 
        .ZN(DP_mult_216_n477) );
  OAI22_X1 DP_mult_216_U786 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1023), 
        .B1(DP_mult_216_n1024), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1022)
         );
  AOI221_X1 DP_mult_216_U785 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[17]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[16]), .A(DP_mult_216_n1022), .ZN(
        DP_mult_216_n1021) );
  XNOR2_X1 DP_mult_216_U784 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1021), 
        .ZN(DP_mult_216_n478) );
  OAI22_X1 DP_mult_216_U783 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1019), 
        .B1(DP_mult_216_n1020), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1018)
         );
  AOI221_X1 DP_mult_216_U782 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[16]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[15]), .A(DP_mult_216_n1018), .ZN(
        DP_mult_216_n1017) );
  XNOR2_X1 DP_mult_216_U781 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1017), 
        .ZN(DP_mult_216_n479) );
  OAI22_X1 DP_mult_216_U780 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1015), 
        .B1(DP_mult_216_n1016), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1014)
         );
  AOI221_X1 DP_mult_216_U779 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[15]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[14]), .A(DP_mult_216_n1014), .ZN(
        DP_mult_216_n1013) );
  XNOR2_X1 DP_mult_216_U778 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1013), 
        .ZN(DP_mult_216_n480) );
  OAI22_X1 DP_mult_216_U777 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1011), 
        .B1(DP_mult_216_n1012), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1010)
         );
  AOI221_X1 DP_mult_216_U776 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[14]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[13]), .A(DP_mult_216_n1010), .ZN(
        DP_mult_216_n1009) );
  XNOR2_X1 DP_mult_216_U775 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1009), 
        .ZN(DP_mult_216_n481) );
  OAI22_X1 DP_mult_216_U774 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1008), 
        .B1(DP_mult_216_n1000), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1007)
         );
  AOI221_X1 DP_mult_216_U773 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[13]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[12]), .A(DP_mult_216_n1007), .ZN(
        DP_mult_216_n1006) );
  XNOR2_X1 DP_mult_216_U772 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1006), 
        .ZN(DP_mult_216_n482) );
  OAI22_X1 DP_mult_216_U771 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n1004), 
        .B1(DP_mult_216_n1005), .B2(DP_mult_216_n969), .ZN(DP_mult_216_n1003)
         );
  AOI221_X1 DP_mult_216_U770 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[12]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[11]), .A(DP_mult_216_n1003), .ZN(
        DP_mult_216_n1002) );
  XNOR2_X1 DP_mult_216_U769 ( .A(DP_mult_216_n974), .B(DP_mult_216_n1002), 
        .ZN(DP_mult_216_n483) );
  OAI22_X1 DP_mult_216_U768 ( .A1(DP_mult_216_n999), .A2(DP_mult_216_n969), 
        .B1(DP_mult_216_n1000), .B2(DP_mult_216_n1001), .ZN(DP_mult_216_n998)
         );
  AOI221_X1 DP_mult_216_U767 ( .B1(DP_mult_216_n966), .B2(DP_pipe00[10]), .C1(
        DP_mult_216_n815), .C2(DP_mult_216_n957), .A(DP_mult_216_n998), .ZN(
        DP_mult_216_n997) );
  XNOR2_X1 DP_mult_216_U766 ( .A(DP_mult_216_n974), .B(DP_mult_216_n997), .ZN(
        DP_mult_216_n484) );
  INV_X1 DP_mult_216_U765 ( .A(DP_mult_216_n816), .ZN(DP_mult_216_n994) );
  OAI22_X1 DP_mult_216_U764 ( .A1(DP_mult_216_n967), .A2(DP_mult_216_n994), 
        .B1(DP_mult_216_n995), .B2(DP_mult_216_n968), .ZN(DP_mult_216_n993) );
  AOI221_X1 DP_mult_216_U763 ( .B1(DP_mult_216_n992), .B2(DP_pipe00[10]), .C1(
        DP_mult_216_n966), .C2(DP_pipe00[9]), .A(DP_mult_216_n993), .ZN(
        DP_mult_216_n991) );
  XNOR2_X1 DP_mult_216_U762 ( .A(DP_mult_216_n974), .B(DP_mult_216_n991), .ZN(
        DP_mult_216_n485) );
  NOR2_X1 DP_mult_216_U761 ( .A1(DP_pipe00[22]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n497) );
  NOR2_X1 DP_mult_216_U760 ( .A1(DP_pipe00[21]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n498) );
  NOR2_X1 DP_mult_216_U759 ( .A1(DP_pipe00[20]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n499) );
  NOR2_X1 DP_mult_216_U758 ( .A1(DP_pipe00[19]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n500) );
  NOR2_X1 DP_mult_216_U757 ( .A1(DP_pipe00[18]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n501) );
  NOR2_X1 DP_mult_216_U756 ( .A1(DP_pipe00[17]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n502) );
  NOR2_X1 DP_mult_216_U755 ( .A1(DP_pipe00[16]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n503) );
  NOR2_X1 DP_mult_216_U754 ( .A1(DP_pipe00[15]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n504) );
  NOR2_X1 DP_mult_216_U753 ( .A1(DP_pipe00[14]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n505) );
  NOR2_X1 DP_mult_216_U752 ( .A1(DP_pipe00[13]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n506) );
  NOR2_X1 DP_mult_216_U751 ( .A1(DP_pipe00[12]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n507) );
  NOR2_X1 DP_mult_216_U750 ( .A1(DP_pipe00[11]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n508) );
  NOR2_X1 DP_mult_216_U749 ( .A1(DP_pipe00[10]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n509) );
  NOR2_X1 DP_mult_216_U748 ( .A1(DP_pipe00[9]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n510) );
  NOR2_X1 DP_mult_216_U747 ( .A1(DP_pipe00[8]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n511) );
  NOR2_X1 DP_mult_216_U746 ( .A1(DP_pipe00[7]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n512) );
  NOR2_X1 DP_mult_216_U745 ( .A1(DP_pipe00[6]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n513) );
  NOR2_X1 DP_mult_216_U744 ( .A1(DP_pipe00[5]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n514) );
  NOR2_X1 DP_mult_216_U743 ( .A1(DP_pipe00[4]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n515) );
  NOR2_X1 DP_mult_216_U742 ( .A1(DP_pipe00[3]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n516) );
  NOR2_X1 DP_mult_216_U741 ( .A1(DP_pipe00[2]), .A2(DP_mult_216_n965), .ZN(
        DP_mult_216_n517) );
  NOR2_X1 DP_mult_216_U740 ( .A1(DP_pipe00[1]), .A2(DP_mult_216_n964), .ZN(
        DP_mult_216_n518) );
  INV_X1 DP_mult_216_U739 ( .A(DP_mult_216_n135), .ZN(DP_mult_216_n987) );
  OAI21_X1 DP_mult_216_U738 ( .B1(DP_mult_216_n960), .B2(DP_mult_216_n963), 
        .A(DP_pipe00[23]), .ZN(DP_mult_216_n985) );
  XNOR2_X1 DP_mult_216_U737 ( .A(DP_mult_216_n985), .B(DP_mult_216_n980), .ZN(
        DP_mult_216_n984) );
  OAI222_X1 DP_mult_216_U736 ( .A1(DP_mult_216_n172), .A2(DP_mult_216_n987), 
        .B1(DP_mult_216_n984), .B2(DP_mult_216_n987), .C1(DP_mult_216_n172), 
        .C2(DP_mult_216_n984), .ZN(DP_mult_216_n986) );
  XOR2_X1 DP_mult_216_U735 ( .A(DP_mult_216_n986), .B(DP_mult_216_n980), .Z(
        DP_mult_216_n982) );
  XOR2_X1 DP_mult_216_U734 ( .A(DP_mult_216_n984), .B(DP_mult_216_n985), .Z(
        DP_mult_216_n983) );
  XOR2_X1 DP_mult_216_U733 ( .A(DP_mult_216_n982), .B(DP_mult_216_n983), .Z(
        DP_pipe0_b0[23]) );
  INV_X1 DP_mult_216_U732 ( .A(DP_b_int_0__3_), .ZN(DP_mult_216_n975) );
  BUF_X1 DP_mult_216_U731 ( .A(DP_b_int_0__11_), .Z(DP_mult_216_n981) );
  INV_X1 DP_mult_216_U730 ( .A(DP_b_int_0__6_), .ZN(DP_mult_216_n977) );
  INV_X1 DP_mult_216_U729 ( .A(DP_b_int_0__9_), .ZN(DP_mult_216_n979) );
  BUF_X1 DP_mult_216_U728 ( .A(DP_b_int_0__11_), .Z(DP_mult_216_n980) );
  INV_X1 DP_mult_216_U727 ( .A(DP_pipe00[0]), .ZN(DP_mult_216_n1056) );
  BUF_X1 DP_mult_216_U726 ( .A(DP_mult_216_n989), .Z(DP_mult_216_n963) );
  BUF_X1 DP_mult_216_U725 ( .A(DP_mult_216_n988), .Z(DP_mult_216_n961) );
  OR2_X1 DP_mult_216_U724 ( .A1(DP_mult_216_n1263), .A2(DP_mult_216_n1258), 
        .ZN(DP_mult_216_n958) );
  BUF_X1 DP_mult_216_U723 ( .A(DP_mult_216_n990), .Z(DP_mult_216_n965) );
  BUF_X1 DP_mult_216_U722 ( .A(DP_mult_216_n989), .Z(DP_mult_216_n962) );
  BUF_X1 DP_mult_216_U721 ( .A(DP_mult_216_n988), .Z(DP_mult_216_n960) );
  BUF_X1 DP_mult_216_U720 ( .A(DP_mult_216_n988), .Z(DP_mult_216_n959) );
  INV_X1 DP_mult_216_U719 ( .A(DP_mult_216_n979), .ZN(DP_mult_216_n978) );
  INV_X1 DP_mult_216_U718 ( .A(DP_mult_216_n977), .ZN(DP_mult_216_n976) );
  INV_X1 DP_mult_216_U717 ( .A(DP_mult_216_n975), .ZN(DP_mult_216_n974) );
  NAND2_X1 DP_mult_216_U716 ( .A1(DP_mult_216_n1190), .A2(DP_mult_216_n1192), 
        .ZN(DP_mult_216_n1135) );
  NAND2_X1 DP_mult_216_U715 ( .A1(DP_mult_216_n1129), .A2(DP_mult_216_n1131), 
        .ZN(DP_mult_216_n1058) );
  NOR2_X2 DP_mult_216_U714 ( .A1(DP_mult_216_n1192), .A2(DP_mult_216_n1193), 
        .ZN(DP_mult_216_n1139) );
  NOR2_X2 DP_mult_216_U713 ( .A1(DP_mult_216_n1131), .A2(DP_mult_216_n1132), 
        .ZN(DP_mult_216_n1064) );
  NOR2_X2 DP_mult_216_U712 ( .A1(DP_mult_216_n1190), .A2(DP_mult_216_n1191), 
        .ZN(DP_mult_216_n1140) );
  NOR2_X2 DP_mult_216_U711 ( .A1(DP_mult_216_n1129), .A2(DP_mult_216_n1130), 
        .ZN(DP_mult_216_n1065) );
  AND2_X1 DP_mult_216_U710 ( .A1(DP_mult_216_n1263), .A2(DP_mult_216_n1257), 
        .ZN(DP_mult_216_n957) );
  BUF_X1 DP_mult_216_U709 ( .A(DP_mult_216_n990), .Z(DP_mult_216_n964) );
  NOR2_X2 DP_mult_216_U708 ( .A1(DP_mult_216_n1257), .A2(DP_mult_216_n1256), 
        .ZN(DP_mult_216_n992) );
  BUF_X1 DP_mult_216_U707 ( .A(DP_mult_216_n1142), .Z(DP_mult_216_n973) );
  BUF_X1 DP_mult_216_U706 ( .A(DP_mult_216_n1068), .Z(DP_mult_216_n971) );
  BUF_X1 DP_mult_216_U705 ( .A(DP_mult_216_n996), .Z(DP_mult_216_n969) );
  BUF_X1 DP_mult_216_U704 ( .A(DP_mult_216_n1142), .Z(DP_mult_216_n972) );
  BUF_X1 DP_mult_216_U703 ( .A(DP_mult_216_n1068), .Z(DP_mult_216_n970) );
  BUF_X1 DP_mult_216_U702 ( .A(DP_mult_216_n996), .Z(DP_mult_216_n968) );
  INV_X1 DP_mult_216_U701 ( .A(DP_mult_216_n958), .ZN(DP_mult_216_n966) );
  INV_X1 DP_mult_216_U700 ( .A(DP_mult_216_n957), .ZN(DP_mult_216_n967) );
  HA_X1 DP_mult_216_U696 ( .A(DP_pipe00[0]), .B(DP_pipe00[1]), .CO(
        DP_mult_216_n394), .S(DP_mult_216_n825) );
  FA_X1 DP_mult_216_U695 ( .A(DP_pipe00[1]), .B(DP_pipe00[2]), .CI(
        DP_mult_216_n394), .CO(DP_mult_216_n393), .S(DP_mult_216_n824) );
  FA_X1 DP_mult_216_U694 ( .A(DP_pipe00[2]), .B(DP_pipe00[3]), .CI(
        DP_mult_216_n393), .CO(DP_mult_216_n392), .S(DP_mult_216_n823) );
  FA_X1 DP_mult_216_U693 ( .A(DP_pipe00[3]), .B(DP_pipe00[4]), .CI(
        DP_mult_216_n392), .CO(DP_mult_216_n391), .S(DP_mult_216_n822) );
  FA_X1 DP_mult_216_U692 ( .A(DP_pipe00[4]), .B(DP_pipe00[5]), .CI(
        DP_mult_216_n391), .CO(DP_mult_216_n390), .S(DP_mult_216_n821) );
  FA_X1 DP_mult_216_U691 ( .A(DP_pipe00[5]), .B(DP_pipe00[6]), .CI(
        DP_mult_216_n390), .CO(DP_mult_216_n389), .S(DP_mult_216_n820) );
  FA_X1 DP_mult_216_U690 ( .A(DP_pipe00[6]), .B(DP_pipe00[7]), .CI(
        DP_mult_216_n389), .CO(DP_mult_216_n388), .S(DP_mult_216_n819) );
  FA_X1 DP_mult_216_U689 ( .A(DP_pipe00[7]), .B(DP_pipe00[8]), .CI(
        DP_mult_216_n388), .CO(DP_mult_216_n387), .S(DP_mult_216_n818) );
  FA_X1 DP_mult_216_U688 ( .A(DP_pipe00[8]), .B(DP_pipe00[9]), .CI(
        DP_mult_216_n387), .CO(DP_mult_216_n386), .S(DP_mult_216_n817) );
  FA_X1 DP_mult_216_U687 ( .A(DP_pipe00[9]), .B(DP_pipe00[10]), .CI(
        DP_mult_216_n386), .CO(DP_mult_216_n385), .S(DP_mult_216_n816) );
  FA_X1 DP_mult_216_U686 ( .A(DP_pipe00[10]), .B(DP_pipe00[11]), .CI(
        DP_mult_216_n385), .CO(DP_mult_216_n384), .S(DP_mult_216_n815) );
  FA_X1 DP_mult_216_U685 ( .A(DP_pipe00[11]), .B(DP_pipe00[12]), .CI(
        DP_mult_216_n384), .CO(DP_mult_216_n383), .S(DP_mult_216_n814) );
  FA_X1 DP_mult_216_U684 ( .A(DP_pipe00[12]), .B(DP_pipe00[13]), .CI(
        DP_mult_216_n383), .CO(DP_mult_216_n382), .S(DP_mult_216_n813) );
  FA_X1 DP_mult_216_U683 ( .A(DP_pipe00[13]), .B(DP_pipe00[14]), .CI(
        DP_mult_216_n382), .CO(DP_mult_216_n381), .S(DP_mult_216_n812) );
  FA_X1 DP_mult_216_U682 ( .A(DP_pipe00[14]), .B(DP_pipe00[15]), .CI(
        DP_mult_216_n381), .CO(DP_mult_216_n380), .S(DP_mult_216_n811) );
  FA_X1 DP_mult_216_U681 ( .A(DP_pipe00[15]), .B(DP_pipe00[16]), .CI(
        DP_mult_216_n380), .CO(DP_mult_216_n379), .S(DP_mult_216_n810) );
  FA_X1 DP_mult_216_U680 ( .A(DP_pipe00[16]), .B(DP_pipe00[17]), .CI(
        DP_mult_216_n379), .CO(DP_mult_216_n378), .S(DP_mult_216_n809) );
  FA_X1 DP_mult_216_U679 ( .A(DP_pipe00[17]), .B(DP_pipe00[18]), .CI(
        DP_mult_216_n378), .CO(DP_mult_216_n377), .S(DP_mult_216_n808) );
  FA_X1 DP_mult_216_U678 ( .A(DP_pipe00[18]), .B(DP_pipe00[19]), .CI(
        DP_mult_216_n377), .CO(DP_mult_216_n376), .S(DP_mult_216_n807) );
  FA_X1 DP_mult_216_U677 ( .A(DP_pipe00[19]), .B(DP_pipe00[20]), .CI(
        DP_mult_216_n376), .CO(DP_mult_216_n375), .S(DP_mult_216_n806) );
  FA_X1 DP_mult_216_U676 ( .A(DP_pipe00[20]), .B(DP_pipe00[21]), .CI(
        DP_mult_216_n375), .CO(DP_mult_216_n374), .S(DP_mult_216_n805) );
  FA_X1 DP_mult_216_U675 ( .A(DP_pipe00[21]), .B(DP_pipe00[22]), .CI(
        DP_mult_216_n374), .CO(DP_mult_216_n373), .S(DP_mult_216_n804) );
  FA_X1 DP_mult_216_U674 ( .A(DP_pipe00[22]), .B(DP_pipe00[23]), .CI(
        DP_mult_216_n373), .CO(DP_mult_216_n802), .S(DP_mult_216_n803) );
  HA_X1 DP_mult_216_U210 ( .A(DP_mult_216_n518), .B(DP_mult_216_n974), .CO(
        DP_mult_216_n362), .S(DP_mult_216_n363) );
  HA_X1 DP_mult_216_U209 ( .A(DP_mult_216_n362), .B(DP_mult_216_n517), .CO(
        DP_mult_216_n360), .S(DP_mult_216_n361) );
  HA_X1 DP_mult_216_U208 ( .A(DP_mult_216_n360), .B(DP_mult_216_n516), .CO(
        DP_mult_216_n358), .S(DP_mult_216_n359) );
  HA_X1 DP_mult_216_U207 ( .A(DP_mult_216_n515), .B(DP_mult_216_n976), .CO(
        DP_mult_216_n356), .S(DP_mult_216_n357) );
  FA_X1 DP_mult_216_U206 ( .A(DP_mult_216_n358), .B(DP_mult_216_n357), .CI(
        DP_mult_216_n469), .CO(DP_mult_216_n354), .S(DP_mult_216_n355) );
  HA_X1 DP_mult_216_U205 ( .A(DP_mult_216_n356), .B(DP_mult_216_n514), .CO(
        DP_mult_216_n352), .S(DP_mult_216_n353) );
  FA_X1 DP_mult_216_U204 ( .A(DP_mult_216_n468), .B(DP_mult_216_n353), .CI(
        DP_mult_216_n354), .CO(DP_mult_216_n350), .S(DP_mult_216_n351) );
  HA_X1 DP_mult_216_U203 ( .A(DP_mult_216_n352), .B(DP_mult_216_n513), .CO(
        DP_mult_216_n348), .S(DP_mult_216_n349) );
  FA_X1 DP_mult_216_U202 ( .A(DP_mult_216_n467), .B(DP_mult_216_n349), .CI(
        DP_mult_216_n350), .CO(DP_mult_216_n346), .S(DP_mult_216_n347) );
  HA_X1 DP_mult_216_U201 ( .A(DP_mult_216_n512), .B(DP_mult_216_n978), .CO(
        DP_mult_216_n344), .S(DP_mult_216_n345) );
  FA_X1 DP_mult_216_U200 ( .A(DP_mult_216_n348), .B(DP_mult_216_n345), .CI(
        DP_mult_216_n443), .CO(DP_mult_216_n342), .S(DP_mult_216_n343) );
  FA_X1 DP_mult_216_U199 ( .A(DP_mult_216_n343), .B(DP_mult_216_n466), .CI(
        DP_mult_216_n346), .CO(DP_mult_216_n340), .S(DP_mult_216_n341) );
  HA_X1 DP_mult_216_U198 ( .A(DP_mult_216_n344), .B(DP_mult_216_n511), .CO(
        DP_mult_216_n338), .S(DP_mult_216_n339) );
  FA_X1 DP_mult_216_U197 ( .A(DP_mult_216_n442), .B(DP_mult_216_n339), .CI(
        DP_mult_216_n342), .CO(DP_mult_216_n336), .S(DP_mult_216_n337) );
  FA_X1 DP_mult_216_U196 ( .A(DP_mult_216_n337), .B(DP_mult_216_n465), .CI(
        DP_mult_216_n340), .CO(DP_mult_216_n334), .S(DP_mult_216_n335) );
  HA_X1 DP_mult_216_U195 ( .A(DP_mult_216_n338), .B(DP_mult_216_n510), .CO(
        DP_mult_216_n332), .S(DP_mult_216_n333) );
  FA_X1 DP_mult_216_U194 ( .A(DP_mult_216_n441), .B(DP_mult_216_n333), .CI(
        DP_mult_216_n336), .CO(DP_mult_216_n330), .S(DP_mult_216_n331) );
  FA_X1 DP_mult_216_U193 ( .A(DP_mult_216_n331), .B(DP_mult_216_n464), .CI(
        DP_mult_216_n334), .CO(DP_mult_216_n328), .S(DP_mult_216_n329) );
  HA_X1 DP_mult_216_U192 ( .A(DP_mult_216_n509), .B(DP_mult_216_n980), .CO(
        DP_mult_216_n326), .S(DP_mult_216_n327) );
  FA_X1 DP_mult_216_U191 ( .A(DP_mult_216_n332), .B(DP_mult_216_n327), .CI(
        DP_mult_216_n417), .CO(DP_mult_216_n324), .S(DP_mult_216_n325) );
  FA_X1 DP_mult_216_U190 ( .A(DP_mult_216_n325), .B(DP_mult_216_n440), .CI(
        DP_mult_216_n330), .CO(DP_mult_216_n322), .S(DP_mult_216_n323) );
  FA_X1 DP_mult_216_U189 ( .A(DP_mult_216_n323), .B(DP_mult_216_n463), .CI(
        DP_mult_216_n328), .CO(DP_mult_216_n320), .S(DP_mult_216_n321) );
  HA_X1 DP_mult_216_U188 ( .A(DP_mult_216_n326), .B(DP_mult_216_n508), .CO(
        DP_mult_216_n318), .S(DP_mult_216_n319) );
  FA_X1 DP_mult_216_U187 ( .A(DP_mult_216_n416), .B(DP_mult_216_n319), .CI(
        DP_mult_216_n324), .CO(DP_mult_216_n316), .S(DP_mult_216_n317) );
  FA_X1 DP_mult_216_U186 ( .A(DP_mult_216_n317), .B(DP_mult_216_n439), .CI(
        DP_mult_216_n322), .CO(DP_mult_216_n314), .S(DP_mult_216_n315) );
  FA_X1 DP_mult_216_U185 ( .A(DP_mult_216_n315), .B(DP_mult_216_n462), .CI(
        DP_mult_216_n320), .CO(DP_mult_216_n312), .S(DP_mult_216_n313) );
  HA_X1 DP_mult_216_U184 ( .A(DP_mult_216_n318), .B(DP_mult_216_n507), .CO(
        DP_mult_216_n310), .S(DP_mult_216_n311) );
  FA_X1 DP_mult_216_U183 ( .A(DP_mult_216_n415), .B(DP_mult_216_n311), .CI(
        DP_mult_216_n316), .CO(DP_mult_216_n308), .S(DP_mult_216_n309) );
  FA_X1 DP_mult_216_U182 ( .A(DP_mult_216_n309), .B(DP_mult_216_n438), .CI(
        DP_mult_216_n314), .CO(DP_mult_216_n306), .S(DP_mult_216_n307) );
  FA_X1 DP_mult_216_U181 ( .A(DP_mult_216_n307), .B(DP_mult_216_n461), .CI(
        DP_mult_216_n312), .CO(DP_mult_216_n304), .S(DP_mult_216_n305) );
  HA_X1 DP_mult_216_U180 ( .A(DP_mult_216_n310), .B(DP_mult_216_n506), .CO(
        DP_mult_216_n302), .S(DP_mult_216_n303) );
  FA_X1 DP_mult_216_U179 ( .A(DP_mult_216_n414), .B(DP_mult_216_n303), .CI(
        DP_mult_216_n308), .CO(DP_mult_216_n300), .S(DP_mult_216_n301) );
  FA_X1 DP_mult_216_U178 ( .A(DP_mult_216_n301), .B(DP_mult_216_n437), .CI(
        DP_mult_216_n306), .CO(DP_mult_216_n298), .S(DP_mult_216_n299) );
  FA_X1 DP_mult_216_U177 ( .A(DP_mult_216_n299), .B(DP_mult_216_n460), .CI(
        DP_mult_216_n304), .CO(DP_mult_216_n296), .S(DP_mult_216_n297) );
  HA_X1 DP_mult_216_U176 ( .A(DP_mult_216_n302), .B(DP_mult_216_n505), .CO(
        DP_mult_216_n294), .S(DP_mult_216_n295) );
  FA_X1 DP_mult_216_U175 ( .A(DP_mult_216_n413), .B(DP_mult_216_n295), .CI(
        DP_mult_216_n300), .CO(DP_mult_216_n292), .S(DP_mult_216_n293) );
  FA_X1 DP_mult_216_U174 ( .A(DP_mult_216_n293), .B(DP_mult_216_n436), .CI(
        DP_mult_216_n298), .CO(DP_mult_216_n290), .S(DP_mult_216_n291) );
  FA_X1 DP_mult_216_U173 ( .A(DP_mult_216_n291), .B(DP_mult_216_n459), .CI(
        DP_mult_216_n296), .CO(DP_mult_216_n288), .S(DP_mult_216_n289) );
  HA_X1 DP_mult_216_U172 ( .A(DP_mult_216_n294), .B(DP_mult_216_n504), .CO(
        DP_mult_216_n286), .S(DP_mult_216_n287) );
  FA_X1 DP_mult_216_U171 ( .A(DP_mult_216_n412), .B(DP_mult_216_n287), .CI(
        DP_mult_216_n292), .CO(DP_mult_216_n284), .S(DP_mult_216_n285) );
  FA_X1 DP_mult_216_U170 ( .A(DP_mult_216_n285), .B(DP_mult_216_n435), .CI(
        DP_mult_216_n290), .CO(DP_mult_216_n282), .S(DP_mult_216_n283) );
  FA_X1 DP_mult_216_U169 ( .A(DP_mult_216_n283), .B(DP_mult_216_n458), .CI(
        DP_mult_216_n288), .CO(DP_mult_216_n280), .S(DP_mult_216_n281) );
  HA_X1 DP_mult_216_U168 ( .A(DP_mult_216_n286), .B(DP_mult_216_n503), .CO(
        DP_mult_216_n278), .S(DP_mult_216_n279) );
  FA_X1 DP_mult_216_U167 ( .A(DP_mult_216_n411), .B(DP_mult_216_n279), .CI(
        DP_mult_216_n284), .CO(DP_mult_216_n276), .S(DP_mult_216_n277) );
  FA_X1 DP_mult_216_U166 ( .A(DP_mult_216_n277), .B(DP_mult_216_n434), .CI(
        DP_mult_216_n282), .CO(DP_mult_216_n274), .S(DP_mult_216_n275) );
  FA_X1 DP_mult_216_U165 ( .A(DP_mult_216_n275), .B(DP_mult_216_n457), .CI(
        DP_mult_216_n280), .CO(DP_mult_216_n272), .S(DP_mult_216_n273) );
  HA_X1 DP_mult_216_U164 ( .A(DP_mult_216_n278), .B(DP_mult_216_n502), .CO(
        DP_mult_216_n270), .S(DP_mult_216_n271) );
  FA_X1 DP_mult_216_U163 ( .A(DP_mult_216_n410), .B(DP_mult_216_n271), .CI(
        DP_mult_216_n276), .CO(DP_mult_216_n268), .S(DP_mult_216_n269) );
  FA_X1 DP_mult_216_U162 ( .A(DP_mult_216_n269), .B(DP_mult_216_n433), .CI(
        DP_mult_216_n274), .CO(DP_mult_216_n266), .S(DP_mult_216_n267) );
  FA_X1 DP_mult_216_U161 ( .A(DP_mult_216_n267), .B(DP_mult_216_n456), .CI(
        DP_mult_216_n272), .CO(DP_mult_216_n264), .S(DP_mult_216_n265) );
  HA_X1 DP_mult_216_U160 ( .A(DP_mult_216_n270), .B(DP_mult_216_n501), .CO(
        DP_mult_216_n262), .S(DP_mult_216_n263) );
  FA_X1 DP_mult_216_U159 ( .A(DP_mult_216_n409), .B(DP_mult_216_n263), .CI(
        DP_mult_216_n268), .CO(DP_mult_216_n260), .S(DP_mult_216_n261) );
  FA_X1 DP_mult_216_U158 ( .A(DP_mult_216_n261), .B(DP_mult_216_n432), .CI(
        DP_mult_216_n266), .CO(DP_mult_216_n258), .S(DP_mult_216_n259) );
  FA_X1 DP_mult_216_U157 ( .A(DP_mult_216_n259), .B(DP_mult_216_n455), .CI(
        DP_mult_216_n264), .CO(DP_mult_216_n256), .S(DP_mult_216_n257) );
  HA_X1 DP_mult_216_U156 ( .A(DP_mult_216_n262), .B(DP_mult_216_n500), .CO(
        DP_mult_216_n254), .S(DP_mult_216_n255) );
  FA_X1 DP_mult_216_U155 ( .A(DP_mult_216_n408), .B(DP_mult_216_n255), .CI(
        DP_mult_216_n260), .CO(DP_mult_216_n252), .S(DP_mult_216_n253) );
  FA_X1 DP_mult_216_U154 ( .A(DP_mult_216_n253), .B(DP_mult_216_n431), .CI(
        DP_mult_216_n258), .CO(DP_mult_216_n250), .S(DP_mult_216_n251) );
  FA_X1 DP_mult_216_U153 ( .A(DP_mult_216_n251), .B(DP_mult_216_n454), .CI(
        DP_mult_216_n256), .CO(DP_mult_216_n248), .S(DP_mult_216_n249) );
  HA_X1 DP_mult_216_U152 ( .A(DP_mult_216_n254), .B(DP_mult_216_n499), .CO(
        DP_mult_216_n246), .S(DP_mult_216_n247) );
  FA_X1 DP_mult_216_U151 ( .A(DP_mult_216_n407), .B(DP_mult_216_n247), .CI(
        DP_mult_216_n252), .CO(DP_mult_216_n244), .S(DP_mult_216_n245) );
  FA_X1 DP_mult_216_U150 ( .A(DP_mult_216_n245), .B(DP_mult_216_n430), .CI(
        DP_mult_216_n250), .CO(DP_mult_216_n242), .S(DP_mult_216_n243) );
  FA_X1 DP_mult_216_U149 ( .A(DP_mult_216_n243), .B(DP_mult_216_n453), .CI(
        DP_mult_216_n248), .CO(DP_mult_216_n240), .S(DP_mult_216_n241) );
  HA_X1 DP_mult_216_U148 ( .A(DP_mult_216_n246), .B(DP_mult_216_n498), .CO(
        DP_mult_216_n238), .S(DP_mult_216_n239) );
  FA_X1 DP_mult_216_U147 ( .A(DP_mult_216_n406), .B(DP_mult_216_n239), .CI(
        DP_mult_216_n244), .CO(DP_mult_216_n236), .S(DP_mult_216_n237) );
  FA_X1 DP_mult_216_U146 ( .A(DP_mult_216_n237), .B(DP_mult_216_n429), .CI(
        DP_mult_216_n242), .CO(DP_mult_216_n234), .S(DP_mult_216_n235) );
  FA_X1 DP_mult_216_U145 ( .A(DP_mult_216_n235), .B(DP_mult_216_n452), .CI(
        DP_mult_216_n240), .CO(DP_mult_216_n232), .S(DP_mult_216_n233) );
  HA_X1 DP_mult_216_U144 ( .A(DP_mult_216_n238), .B(DP_mult_216_n497), .CO(
        DP_mult_216_n230), .S(DP_mult_216_n231) );
  FA_X1 DP_mult_216_U143 ( .A(DP_mult_216_n405), .B(DP_mult_216_n231), .CI(
        DP_mult_216_n236), .CO(DP_mult_216_n228), .S(DP_mult_216_n229) );
  FA_X1 DP_mult_216_U142 ( .A(DP_mult_216_n229), .B(DP_mult_216_n428), .CI(
        DP_mult_216_n234), .CO(DP_mult_216_n226), .S(DP_mult_216_n227) );
  FA_X1 DP_mult_216_U141 ( .A(DP_mult_216_n227), .B(DP_mult_216_n451), .CI(
        DP_mult_216_n232), .CO(DP_mult_216_n224), .S(DP_mult_216_n225) );
  FA_X1 DP_mult_216_U138 ( .A(DP_mult_216_n404), .B(DP_mult_216_n223), .CI(
        DP_mult_216_n228), .CO(DP_mult_216_n221), .S(DP_mult_216_n222) );
  FA_X1 DP_mult_216_U137 ( .A(DP_mult_216_n222), .B(DP_mult_216_n427), .CI(
        DP_mult_216_n226), .CO(DP_mult_216_n219), .S(DP_mult_216_n220) );
  FA_X1 DP_mult_216_U136 ( .A(DP_mult_216_n220), .B(DP_mult_216_n450), .CI(
        DP_mult_216_n224), .CO(DP_mult_216_n217), .S(DP_mult_216_n218) );
  FA_X1 DP_mult_216_U134 ( .A(DP_mult_216_n403), .B(DP_mult_216_n216), .CI(
        DP_mult_216_n221), .CO(DP_mult_216_n214), .S(DP_mult_216_n215) );
  FA_X1 DP_mult_216_U133 ( .A(DP_mult_216_n215), .B(DP_mult_216_n426), .CI(
        DP_mult_216_n219), .CO(DP_mult_216_n212), .S(DP_mult_216_n213) );
  FA_X1 DP_mult_216_U132 ( .A(DP_mult_216_n213), .B(DP_mult_216_n449), .CI(
        DP_mult_216_n217), .CO(DP_mult_216_n210), .S(DP_mult_216_n211) );
  FA_X1 DP_mult_216_U130 ( .A(DP_mult_216_n402), .B(DP_mult_216_n216), .CI(
        DP_mult_216_n214), .CO(DP_mult_216_n206), .S(DP_mult_216_n207) );
  FA_X1 DP_mult_216_U129 ( .A(DP_mult_216_n207), .B(DP_mult_216_n425), .CI(
        DP_mult_216_n212), .CO(DP_mult_216_n204), .S(DP_mult_216_n205) );
  FA_X1 DP_mult_216_U128 ( .A(DP_mult_216_n205), .B(DP_mult_216_n448), .CI(
        DP_mult_216_n471), .CO(DP_mult_216_n202), .S(DP_mult_216_n203) );
  FA_X1 DP_mult_216_U127 ( .A(DP_mult_216_n208), .B(DP_mult_216_n470), .CI(
        DP_mult_216_n401), .CO(DP_mult_216_n200), .S(DP_mult_216_n201) );
  FA_X1 DP_mult_216_U126 ( .A(DP_mult_216_n206), .B(DP_mult_216_n201), .CI(
        DP_mult_216_n424), .CO(DP_mult_216_n198), .S(DP_mult_216_n199) );
  FA_X1 DP_mult_216_U125 ( .A(DP_mult_216_n204), .B(DP_mult_216_n199), .CI(
        DP_mult_216_n447), .CO(DP_mult_216_n196), .S(DP_mult_216_n197) );
  FA_X1 DP_mult_216_U123 ( .A(DP_mult_216_n195), .B(DP_mult_216_n200), .CI(
        DP_mult_216_n198), .CO(DP_mult_216_n193), .S(DP_mult_216_n194) );
  FA_X1 DP_mult_216_U122 ( .A(DP_mult_216_n194), .B(DP_mult_216_n423), .CI(
        DP_mult_216_n446), .CO(DP_mult_216_n191), .S(DP_mult_216_n192) );
  FA_X1 DP_mult_216_U120 ( .A(DP_mult_216_n400), .B(DP_mult_216_n195), .CI(
        DP_mult_216_n193), .CO(DP_mult_216_n187), .S(DP_mult_216_n188) );
  FA_X1 DP_mult_216_U119 ( .A(DP_mult_216_n445), .B(DP_mult_216_n422), .CI(
        DP_mult_216_n188), .CO(DP_mult_216_n185), .S(DP_mult_216_n186) );
  FA_X1 DP_mult_216_U118 ( .A(DP_mult_216_n189), .B(DP_mult_216_n444), .CI(
        DP_mult_216_n399), .CO(DP_mult_216_n177), .S(DP_mult_216_n184) );
  FA_X1 DP_mult_216_U117 ( .A(DP_mult_216_n421), .B(DP_mult_216_n184), .CI(
        DP_mult_216_n187), .CO(DP_mult_216_n182), .S(DP_mult_216_n183) );
  FA_X1 DP_mult_216_U115 ( .A(DP_mult_216_n181), .B(DP_mult_216_n398), .CI(
        DP_mult_216_n420), .CO(DP_mult_216_n179), .S(DP_mult_216_n180) );
  FA_X1 DP_mult_216_U113 ( .A(DP_mult_216_n397), .B(DP_mult_216_n181), .CI(
        DP_mult_216_n419), .CO(DP_mult_216_n175), .S(DP_mult_216_n176) );
  FA_X1 DP_mult_216_U112 ( .A(DP_mult_216_n177), .B(DP_mult_216_n418), .CI(
        DP_mult_216_n396), .CO(DP_mult_216_n173), .S(DP_mult_216_n174) );
  FA_X1 DP_mult_216_U96 ( .A(DP_mult_216_n313), .B(DP_mult_216_n485), .CI(
        DP_mult_216_n158), .CO(DP_mult_216_n157), .S(DP_pipe0_b0[0]) );
  FA_X1 DP_mult_216_U95 ( .A(DP_mult_216_n305), .B(DP_mult_216_n484), .CI(
        DP_mult_216_n157), .CO(DP_mult_216_n156), .S(DP_pipe0_b0[1]) );
  FA_X1 DP_mult_216_U94 ( .A(DP_mult_216_n297), .B(DP_mult_216_n483), .CI(
        DP_mult_216_n156), .CO(DP_mult_216_n155), .S(DP_pipe0_b0[2]) );
  FA_X1 DP_mult_216_U93 ( .A(DP_mult_216_n289), .B(DP_mult_216_n482), .CI(
        DP_mult_216_n155), .CO(DP_mult_216_n154), .S(DP_pipe0_b0[3]) );
  FA_X1 DP_mult_216_U92 ( .A(DP_mult_216_n281), .B(DP_mult_216_n481), .CI(
        DP_mult_216_n154), .CO(DP_mult_216_n153), .S(DP_pipe0_b0[4]) );
  FA_X1 DP_mult_216_U91 ( .A(DP_mult_216_n273), .B(DP_mult_216_n480), .CI(
        DP_mult_216_n153), .CO(DP_mult_216_n152), .S(DP_pipe0_b0[5]) );
  FA_X1 DP_mult_216_U90 ( .A(DP_mult_216_n265), .B(DP_mult_216_n479), .CI(
        DP_mult_216_n152), .CO(DP_mult_216_n151), .S(DP_pipe0_b0[6]) );
  FA_X1 DP_mult_216_U89 ( .A(DP_mult_216_n257), .B(DP_mult_216_n478), .CI(
        DP_mult_216_n151), .CO(DP_mult_216_n150), .S(DP_pipe0_b0[7]) );
  FA_X1 DP_mult_216_U88 ( .A(DP_mult_216_n249), .B(DP_mult_216_n477), .CI(
        DP_mult_216_n150), .CO(DP_mult_216_n149), .S(DP_pipe0_b0[8]) );
  FA_X1 DP_mult_216_U87 ( .A(DP_mult_216_n241), .B(DP_mult_216_n476), .CI(
        DP_mult_216_n149), .CO(DP_mult_216_n148), .S(DP_pipe0_b0[9]) );
  FA_X1 DP_mult_216_U86 ( .A(DP_mult_216_n233), .B(DP_mult_216_n475), .CI(
        DP_mult_216_n148), .CO(DP_mult_216_n147), .S(DP_pipe0_b0[10]) );
  FA_X1 DP_mult_216_U85 ( .A(DP_mult_216_n225), .B(DP_mult_216_n474), .CI(
        DP_mult_216_n147), .CO(DP_mult_216_n146), .S(DP_pipe0_b0[11]) );
  FA_X1 DP_mult_216_U84 ( .A(DP_mult_216_n218), .B(DP_mult_216_n473), .CI(
        DP_mult_216_n146), .CO(DP_mult_216_n145), .S(DP_pipe0_b0[12]) );
  FA_X1 DP_mult_216_U83 ( .A(DP_mult_216_n211), .B(DP_mult_216_n472), .CI(
        DP_mult_216_n145), .CO(DP_mult_216_n144), .S(DP_pipe0_b0[13]) );
  FA_X1 DP_mult_216_U82 ( .A(DP_mult_216_n203), .B(DP_mult_216_n210), .CI(
        DP_mult_216_n144), .CO(DP_mult_216_n143), .S(DP_pipe0_b0[14]) );
  FA_X1 DP_mult_216_U81 ( .A(DP_mult_216_n197), .B(DP_mult_216_n202), .CI(
        DP_mult_216_n143), .CO(DP_mult_216_n142), .S(DP_pipe0_b0[15]) );
  FA_X1 DP_mult_216_U80 ( .A(DP_mult_216_n192), .B(DP_mult_216_n196), .CI(
        DP_mult_216_n142), .CO(DP_mult_216_n141), .S(DP_pipe0_b0[16]) );
  FA_X1 DP_mult_216_U79 ( .A(DP_mult_216_n186), .B(DP_mult_216_n191), .CI(
        DP_mult_216_n141), .CO(DP_mult_216_n140), .S(DP_pipe0_b0[17]) );
  FA_X1 DP_mult_216_U78 ( .A(DP_mult_216_n183), .B(DP_mult_216_n185), .CI(
        DP_mult_216_n140), .CO(DP_mult_216_n139), .S(DP_pipe0_b0[18]) );
  FA_X1 DP_mult_216_U77 ( .A(DP_mult_216_n180), .B(DP_mult_216_n182), .CI(
        DP_mult_216_n139), .CO(DP_mult_216_n138), .S(DP_pipe0_b0[19]) );
  FA_X1 DP_mult_216_U76 ( .A(DP_mult_216_n176), .B(DP_mult_216_n179), .CI(
        DP_mult_216_n138), .CO(DP_mult_216_n137), .S(DP_pipe0_b0[20]) );
  FA_X1 DP_mult_216_U75 ( .A(DP_mult_216_n174), .B(DP_mult_216_n175), .CI(
        DP_mult_216_n137), .CO(DP_mult_216_n136), .S(DP_pipe0_b0[21]) );
  FA_X1 DP_mult_216_U74 ( .A(DP_mult_216_n172), .B(DP_mult_216_n173), .CI(
        DP_mult_216_n136), .CO(DP_mult_216_n135), .S(DP_pipe0_b0[22]) );
  INV_X1 DP_mult_214_U1958 ( .A(DP_coeff_ret0[1]), .ZN(DP_mult_214_n2158) );
  NOR2_X1 DP_mult_214_U1957 ( .A1(DP_mult_214_n2158), .A2(DP_coeff_ret0[1]), 
        .ZN(DP_mult_214_n1636) );
  INV_X1 DP_mult_214_U1956 ( .A(DP_coeff_ret0[2]), .ZN(DP_mult_214_n1742) );
  XNOR2_X1 DP_mult_214_U1955 ( .A(DP_coeff_ret0[1]), .B(DP_mult_214_n1742), 
        .ZN(DP_mult_214_n2157) );
  AOI221_X1 DP_mult_214_U1954 ( .B1(DP_sw0_1_), .B2(DP_mult_214_n1563), .C1(
        DP_mult_214_n1396), .C2(DP_mult_214_n1550), .A(DP_mult_214_n1742), 
        .ZN(DP_mult_214_n2159) );
  INV_X1 DP_mult_214_U1953 ( .A(DP_sw0_2_), .ZN(DP_mult_214_n1661) );
  INV_X1 DP_mult_214_U1952 ( .A(DP_mult_214_n1397), .ZN(DP_mult_214_n1650) );
  OAI22_X1 DP_mult_214_U1951 ( .A1(DP_mult_214_n1541), .A2(DP_mult_214_n1661), 
        .B1(DP_mult_214_n1564), .B2(DP_mult_214_n1650), .ZN(DP_mult_214_n2161)
         );
  AOI211_X1 DP_mult_214_U1950 ( .C1(DP_sw0_1_), .C2(DP_mult_214_n1561), .A(
        DP_mult_214_n2161), .B(DP_sw0_0_), .ZN(DP_mult_214_n2160) );
  AND2_X1 DP_mult_214_U1949 ( .A1(DP_mult_214_n2159), .A2(DP_mult_214_n2160), 
        .ZN(DP_mult_214_n2153) );
  INV_X1 DP_mult_214_U1948 ( .A(DP_mult_214_n1395), .ZN(DP_mult_214_n1657) );
  INV_X1 DP_mult_214_U1947 ( .A(DP_sw0_1_), .ZN(DP_mult_214_n1649) );
  OAI22_X1 DP_mult_214_U1946 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1657), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1649), .ZN(DP_mult_214_n2156)
         );
  AOI221_X1 DP_mult_214_U1945 ( .B1(DP_sw0_3_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_2_), .C2(DP_mult_214_n1563), .A(DP_mult_214_n2156), .ZN(
        DP_mult_214_n2155) );
  XNOR2_X1 DP_mult_214_U1944 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2155), 
        .ZN(DP_mult_214_n2154) );
  AOI222_X1 DP_mult_214_U1943 ( .A1(DP_mult_214_n2153), .A2(DP_mult_214_n2154), 
        .B1(DP_mult_214_n2153), .B2(DP_mult_214_n688), .C1(DP_mult_214_n688), 
        .C2(DP_mult_214_n2154), .ZN(DP_mult_214_n2148) );
  INV_X1 DP_mult_214_U1942 ( .A(DP_mult_214_n1394), .ZN(DP_mult_214_n1660) );
  OAI22_X1 DP_mult_214_U1941 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1660), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1661), .ZN(DP_mult_214_n2152)
         );
  AOI221_X1 DP_mult_214_U1940 ( .B1(DP_sw0_4_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_3_), .C2(DP_mult_214_n1563), .A(DP_mult_214_n2152), .ZN(
        DP_mult_214_n2151) );
  XNOR2_X1 DP_mult_214_U1939 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2151), 
        .ZN(DP_mult_214_n2149) );
  INV_X1 DP_mult_214_U1938 ( .A(DP_mult_214_n686), .ZN(DP_mult_214_n2150) );
  OAI222_X1 DP_mult_214_U1937 ( .A1(DP_mult_214_n2148), .A2(DP_mult_214_n2149), 
        .B1(DP_mult_214_n2148), .B2(DP_mult_214_n2150), .C1(DP_mult_214_n2150), 
        .C2(DP_mult_214_n2149), .ZN(DP_mult_214_n2144) );
  INV_X1 DP_mult_214_U1936 ( .A(DP_mult_214_n1393), .ZN(DP_mult_214_n1664) );
  INV_X1 DP_mult_214_U1935 ( .A(DP_sw0_3_), .ZN(DP_mult_214_n1665) );
  OAI22_X1 DP_mult_214_U1934 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1664), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1665), .ZN(DP_mult_214_n2147)
         );
  AOI221_X1 DP_mult_214_U1933 ( .B1(DP_sw0_5_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_4_), .C2(DP_mult_214_n1563), .A(DP_mult_214_n2147), .ZN(
        DP_mult_214_n2146) );
  XNOR2_X1 DP_mult_214_U1932 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2146), 
        .ZN(DP_mult_214_n2145) );
  AOI222_X1 DP_mult_214_U1931 ( .A1(DP_mult_214_n2144), .A2(DP_mult_214_n2145), 
        .B1(DP_mult_214_n2144), .B2(DP_mult_214_n684), .C1(DP_mult_214_n684), 
        .C2(DP_mult_214_n2145), .ZN(DP_mult_214_n2139) );
  INV_X1 DP_mult_214_U1930 ( .A(DP_mult_214_n1392), .ZN(DP_mult_214_n1668) );
  INV_X1 DP_mult_214_U1929 ( .A(DP_sw0_4_), .ZN(DP_mult_214_n1669) );
  OAI22_X1 DP_mult_214_U1928 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1668), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1669), .ZN(DP_mult_214_n2143)
         );
  AOI221_X1 DP_mult_214_U1927 ( .B1(DP_sw0_6_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_5_), .C2(DP_mult_214_n1563), .A(DP_mult_214_n2143), .ZN(
        DP_mult_214_n2142) );
  XNOR2_X1 DP_mult_214_U1926 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2142), 
        .ZN(DP_mult_214_n2140) );
  INV_X1 DP_mult_214_U1925 ( .A(DP_mult_214_n680), .ZN(DP_mult_214_n2141) );
  OAI222_X1 DP_mult_214_U1924 ( .A1(DP_mult_214_n2139), .A2(DP_mult_214_n2140), 
        .B1(DP_mult_214_n2139), .B2(DP_mult_214_n2141), .C1(DP_mult_214_n2141), 
        .C2(DP_mult_214_n2140), .ZN(DP_mult_214_n2135) );
  INV_X1 DP_mult_214_U1923 ( .A(DP_mult_214_n1391), .ZN(DP_mult_214_n1672) );
  INV_X1 DP_mult_214_U1922 ( .A(DP_sw0_5_), .ZN(DP_mult_214_n1673) );
  OAI22_X1 DP_mult_214_U1921 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1672), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1673), .ZN(DP_mult_214_n2138)
         );
  AOI221_X1 DP_mult_214_U1920 ( .B1(DP_sw0_7_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_6_), .C2(DP_mult_214_n1563), .A(DP_mult_214_n2138), .ZN(
        DP_mult_214_n2137) );
  XNOR2_X1 DP_mult_214_U1919 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2137), 
        .ZN(DP_mult_214_n2136) );
  AOI222_X1 DP_mult_214_U1918 ( .A1(DP_mult_214_n2135), .A2(DP_mult_214_n2136), 
        .B1(DP_mult_214_n2135), .B2(DP_mult_214_n676), .C1(DP_mult_214_n676), 
        .C2(DP_mult_214_n2136), .ZN(DP_mult_214_n2130) );
  INV_X1 DP_mult_214_U1917 ( .A(DP_mult_214_n1390), .ZN(DP_mult_214_n1676) );
  INV_X1 DP_mult_214_U1916 ( .A(DP_sw0_6_), .ZN(DP_mult_214_n1677) );
  OAI22_X1 DP_mult_214_U1915 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1676), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1677), .ZN(DP_mult_214_n2134)
         );
  AOI221_X1 DP_mult_214_U1914 ( .B1(DP_sw0_8_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_7_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2134), .ZN(
        DP_mult_214_n2133) );
  XNOR2_X1 DP_mult_214_U1913 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2133), 
        .ZN(DP_mult_214_n2131) );
  INV_X1 DP_mult_214_U1912 ( .A(DP_mult_214_n672), .ZN(DP_mult_214_n2132) );
  OAI222_X1 DP_mult_214_U1911 ( .A1(DP_mult_214_n2130), .A2(DP_mult_214_n2131), 
        .B1(DP_mult_214_n2130), .B2(DP_mult_214_n2132), .C1(DP_mult_214_n2132), 
        .C2(DP_mult_214_n2131), .ZN(DP_mult_214_n2126) );
  INV_X1 DP_mult_214_U1910 ( .A(DP_mult_214_n1389), .ZN(DP_mult_214_n1680) );
  INV_X1 DP_mult_214_U1909 ( .A(DP_sw0_7_), .ZN(DP_mult_214_n1681) );
  OAI22_X1 DP_mult_214_U1908 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1680), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1681), .ZN(DP_mult_214_n2129)
         );
  AOI221_X1 DP_mult_214_U1907 ( .B1(DP_sw0_9_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_8_), .C2(DP_mult_214_n1563), .A(DP_mult_214_n2129), .ZN(
        DP_mult_214_n2128) );
  XNOR2_X1 DP_mult_214_U1906 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2128), 
        .ZN(DP_mult_214_n2127) );
  AOI222_X1 DP_mult_214_U1905 ( .A1(DP_mult_214_n2126), .A2(DP_mult_214_n2127), 
        .B1(DP_mult_214_n2126), .B2(DP_mult_214_n666), .C1(DP_mult_214_n666), 
        .C2(DP_mult_214_n2127), .ZN(DP_mult_214_n2121) );
  INV_X1 DP_mult_214_U1904 ( .A(DP_mult_214_n1388), .ZN(DP_mult_214_n1684) );
  INV_X1 DP_mult_214_U1903 ( .A(DP_sw0_8_), .ZN(DP_mult_214_n1685) );
  OAI22_X1 DP_mult_214_U1902 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1684), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1685), .ZN(DP_mult_214_n2125)
         );
  AOI221_X1 DP_mult_214_U1901 ( .B1(DP_sw0_10_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_9_), .C2(DP_mult_214_n1563), .A(DP_mult_214_n2125), .ZN(
        DP_mult_214_n2124) );
  XNOR2_X1 DP_mult_214_U1900 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2124), 
        .ZN(DP_mult_214_n2122) );
  INV_X1 DP_mult_214_U1899 ( .A(DP_mult_214_n660), .ZN(DP_mult_214_n2123) );
  OAI222_X1 DP_mult_214_U1898 ( .A1(DP_mult_214_n2121), .A2(DP_mult_214_n2122), 
        .B1(DP_mult_214_n2121), .B2(DP_mult_214_n2123), .C1(DP_mult_214_n2123), 
        .C2(DP_mult_214_n2122), .ZN(DP_mult_214_n2117) );
  INV_X1 DP_mult_214_U1897 ( .A(DP_mult_214_n1387), .ZN(DP_mult_214_n1688) );
  INV_X1 DP_mult_214_U1896 ( .A(DP_sw0_9_), .ZN(DP_mult_214_n1689) );
  OAI22_X1 DP_mult_214_U1895 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1688), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1689), .ZN(DP_mult_214_n2120)
         );
  AOI221_X1 DP_mult_214_U1894 ( .B1(DP_sw0_11_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_10_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2120), .ZN(
        DP_mult_214_n2119) );
  XNOR2_X1 DP_mult_214_U1893 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2119), 
        .ZN(DP_mult_214_n2118) );
  AOI222_X1 DP_mult_214_U1892 ( .A1(DP_mult_214_n2117), .A2(DP_mult_214_n2118), 
        .B1(DP_mult_214_n2117), .B2(DP_mult_214_n654), .C1(DP_mult_214_n654), 
        .C2(DP_mult_214_n2118), .ZN(DP_mult_214_n2112) );
  INV_X1 DP_mult_214_U1891 ( .A(DP_mult_214_n1386), .ZN(DP_mult_214_n1692) );
  INV_X1 DP_mult_214_U1890 ( .A(DP_sw0_10_), .ZN(DP_mult_214_n1693) );
  OAI22_X1 DP_mult_214_U1889 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1692), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1693), .ZN(DP_mult_214_n2116)
         );
  AOI221_X1 DP_mult_214_U1888 ( .B1(DP_sw0_12_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_11_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2116), .ZN(
        DP_mult_214_n2115) );
  XNOR2_X1 DP_mult_214_U1887 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2115), 
        .ZN(DP_mult_214_n2113) );
  INV_X1 DP_mult_214_U1886 ( .A(DP_mult_214_n646), .ZN(DP_mult_214_n2114) );
  OAI222_X1 DP_mult_214_U1885 ( .A1(DP_mult_214_n2112), .A2(DP_mult_214_n2113), 
        .B1(DP_mult_214_n2112), .B2(DP_mult_214_n2114), .C1(DP_mult_214_n2114), 
        .C2(DP_mult_214_n2113), .ZN(DP_mult_214_n2108) );
  INV_X1 DP_mult_214_U1884 ( .A(DP_mult_214_n1385), .ZN(DP_mult_214_n1696) );
  INV_X1 DP_mult_214_U1883 ( .A(DP_sw0_11_), .ZN(DP_mult_214_n1697) );
  OAI22_X1 DP_mult_214_U1882 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1696), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1697), .ZN(DP_mult_214_n2111)
         );
  AOI221_X1 DP_mult_214_U1881 ( .B1(DP_sw0_13_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_12_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2111), .ZN(
        DP_mult_214_n2110) );
  XNOR2_X1 DP_mult_214_U1880 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2110), 
        .ZN(DP_mult_214_n2109) );
  AOI222_X1 DP_mult_214_U1879 ( .A1(DP_mult_214_n2108), .A2(DP_mult_214_n2109), 
        .B1(DP_mult_214_n2108), .B2(DP_mult_214_n638), .C1(DP_mult_214_n638), 
        .C2(DP_mult_214_n2109), .ZN(DP_mult_214_n2103) );
  INV_X1 DP_mult_214_U1878 ( .A(DP_mult_214_n1384), .ZN(DP_mult_214_n1700) );
  INV_X1 DP_mult_214_U1877 ( .A(DP_sw0_12_), .ZN(DP_mult_214_n1701) );
  OAI22_X1 DP_mult_214_U1876 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1700), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1701), .ZN(DP_mult_214_n2107)
         );
  AOI221_X1 DP_mult_214_U1875 ( .B1(DP_sw0_14_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_13_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2107), .ZN(
        DP_mult_214_n2106) );
  XNOR2_X1 DP_mult_214_U1874 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2106), 
        .ZN(DP_mult_214_n2104) );
  INV_X1 DP_mult_214_U1873 ( .A(DP_mult_214_n630), .ZN(DP_mult_214_n2105) );
  OAI222_X1 DP_mult_214_U1872 ( .A1(DP_mult_214_n2103), .A2(DP_mult_214_n2104), 
        .B1(DP_mult_214_n2103), .B2(DP_mult_214_n2105), .C1(DP_mult_214_n2105), 
        .C2(DP_mult_214_n2104), .ZN(DP_mult_214_n2099) );
  INV_X1 DP_mult_214_U1871 ( .A(DP_mult_214_n1383), .ZN(DP_mult_214_n1704) );
  INV_X1 DP_mult_214_U1870 ( .A(DP_sw0_13_), .ZN(DP_mult_214_n1705) );
  OAI22_X1 DP_mult_214_U1869 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1704), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1705), .ZN(DP_mult_214_n2102)
         );
  AOI221_X1 DP_mult_214_U1868 ( .B1(DP_sw0_15_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_14_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2102), .ZN(
        DP_mult_214_n2101) );
  XNOR2_X1 DP_mult_214_U1867 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2101), 
        .ZN(DP_mult_214_n2100) );
  AOI222_X1 DP_mult_214_U1866 ( .A1(DP_mult_214_n2099), .A2(DP_mult_214_n2100), 
        .B1(DP_mult_214_n2099), .B2(DP_mult_214_n620), .C1(DP_mult_214_n620), 
        .C2(DP_mult_214_n2100), .ZN(DP_mult_214_n2094) );
  INV_X1 DP_mult_214_U1865 ( .A(DP_mult_214_n1382), .ZN(DP_mult_214_n1708) );
  INV_X1 DP_mult_214_U1864 ( .A(DP_sw0_14_), .ZN(DP_mult_214_n1709) );
  OAI22_X1 DP_mult_214_U1863 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1708), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1709), .ZN(DP_mult_214_n2098)
         );
  AOI221_X1 DP_mult_214_U1862 ( .B1(DP_sw0_16_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_15_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2098), .ZN(
        DP_mult_214_n2097) );
  XNOR2_X1 DP_mult_214_U1861 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2097), 
        .ZN(DP_mult_214_n2095) );
  INV_X1 DP_mult_214_U1860 ( .A(DP_mult_214_n610), .ZN(DP_mult_214_n2096) );
  OAI222_X1 DP_mult_214_U1859 ( .A1(DP_mult_214_n2094), .A2(DP_mult_214_n2095), 
        .B1(DP_mult_214_n2094), .B2(DP_mult_214_n2096), .C1(DP_mult_214_n2096), 
        .C2(DP_mult_214_n2095), .ZN(DP_mult_214_n2090) );
  INV_X1 DP_mult_214_U1858 ( .A(DP_mult_214_n1381), .ZN(DP_mult_214_n1712) );
  INV_X1 DP_mult_214_U1857 ( .A(DP_sw0_15_), .ZN(DP_mult_214_n1713) );
  OAI22_X1 DP_mult_214_U1856 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1712), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1713), .ZN(DP_mult_214_n2093)
         );
  AOI221_X1 DP_mult_214_U1855 ( .B1(DP_sw0_17_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_16_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2093), .ZN(
        DP_mult_214_n2092) );
  XNOR2_X1 DP_mult_214_U1854 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2092), 
        .ZN(DP_mult_214_n2091) );
  AOI222_X1 DP_mult_214_U1853 ( .A1(DP_mult_214_n2090), .A2(DP_mult_214_n2091), 
        .B1(DP_mult_214_n2090), .B2(DP_mult_214_n600), .C1(DP_mult_214_n600), 
        .C2(DP_mult_214_n2091), .ZN(DP_mult_214_n2085) );
  INV_X1 DP_mult_214_U1852 ( .A(DP_mult_214_n1380), .ZN(DP_mult_214_n1716) );
  INV_X1 DP_mult_214_U1851 ( .A(DP_sw0_16_), .ZN(DP_mult_214_n1717) );
  OAI22_X1 DP_mult_214_U1850 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1716), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1717), .ZN(DP_mult_214_n2089)
         );
  AOI221_X1 DP_mult_214_U1849 ( .B1(DP_sw0_18_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_17_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2089), .ZN(
        DP_mult_214_n2088) );
  XNOR2_X1 DP_mult_214_U1848 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2088), 
        .ZN(DP_mult_214_n2086) );
  INV_X1 DP_mult_214_U1847 ( .A(DP_mult_214_n588), .ZN(DP_mult_214_n2087) );
  OAI222_X1 DP_mult_214_U1846 ( .A1(DP_mult_214_n2085), .A2(DP_mult_214_n2086), 
        .B1(DP_mult_214_n2085), .B2(DP_mult_214_n2087), .C1(DP_mult_214_n2087), 
        .C2(DP_mult_214_n2086), .ZN(DP_mult_214_n2081) );
  INV_X1 DP_mult_214_U1845 ( .A(DP_mult_214_n1379), .ZN(DP_mult_214_n1720) );
  INV_X1 DP_mult_214_U1844 ( .A(DP_sw0_17_), .ZN(DP_mult_214_n1721) );
  OAI22_X1 DP_mult_214_U1843 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1720), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1721), .ZN(DP_mult_214_n2084)
         );
  AOI221_X1 DP_mult_214_U1842 ( .B1(DP_sw0_19_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_18_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2084), .ZN(
        DP_mult_214_n2083) );
  XNOR2_X1 DP_mult_214_U1841 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2083), 
        .ZN(DP_mult_214_n2082) );
  AOI222_X1 DP_mult_214_U1840 ( .A1(DP_mult_214_n2081), .A2(DP_mult_214_n2082), 
        .B1(DP_mult_214_n2081), .B2(DP_mult_214_n576), .C1(DP_mult_214_n576), 
        .C2(DP_mult_214_n2082), .ZN(DP_mult_214_n2080) );
  INV_X1 DP_mult_214_U1839 ( .A(DP_mult_214_n2080), .ZN(DP_mult_214_n2076) );
  INV_X1 DP_mult_214_U1838 ( .A(DP_mult_214_n1378), .ZN(DP_mult_214_n1724) );
  INV_X1 DP_mult_214_U1837 ( .A(DP_sw0_18_), .ZN(DP_mult_214_n1725) );
  OAI22_X1 DP_mult_214_U1836 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1724), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1725), .ZN(DP_mult_214_n2079)
         );
  AOI221_X1 DP_mult_214_U1835 ( .B1(DP_sw0_20_), .B2(DP_mult_214_n1561), .C1(
        DP_sw0_19_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2079), .ZN(
        DP_mult_214_n2078) );
  XNOR2_X1 DP_mult_214_U1834 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n2078), 
        .ZN(DP_mult_214_n2077) );
  AOI222_X1 DP_mult_214_U1833 ( .A1(DP_mult_214_n2076), .A2(DP_mult_214_n2077), 
        .B1(DP_mult_214_n2076), .B2(DP_mult_214_n564), .C1(DP_mult_214_n564), 
        .C2(DP_mult_214_n2077), .ZN(DP_mult_214_n2071) );
  INV_X1 DP_mult_214_U1832 ( .A(DP_mult_214_n1377), .ZN(DP_mult_214_n1728) );
  INV_X1 DP_mult_214_U1831 ( .A(DP_sw0_19_), .ZN(DP_mult_214_n1729) );
  OAI22_X1 DP_mult_214_U1830 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1728), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1729), .ZN(DP_mult_214_n2075)
         );
  AOI221_X1 DP_mult_214_U1829 ( .B1(DP_mult_214_n1561), .B2(DP_sw0_21_), .C1(
        DP_sw0_20_), .C2(DP_mult_214_n1562), .A(DP_mult_214_n2075), .ZN(
        DP_mult_214_n2074) );
  XNOR2_X1 DP_mult_214_U1828 ( .A(DP_mult_214_n1742), .B(DP_mult_214_n2074), 
        .ZN(DP_mult_214_n2072) );
  INV_X1 DP_mult_214_U1827 ( .A(DP_mult_214_n550), .ZN(DP_mult_214_n2073) );
  OAI222_X1 DP_mult_214_U1826 ( .A1(DP_mult_214_n2071), .A2(DP_mult_214_n2072), 
        .B1(DP_mult_214_n2071), .B2(DP_mult_214_n2073), .C1(DP_mult_214_n2073), 
        .C2(DP_mult_214_n2072), .ZN(DP_mult_214_n326) );
  XNOR2_X1 DP_mult_214_U1825 ( .A(DP_coeff_ret0[21]), .B(DP_mult_214_n1608), 
        .ZN(DP_mult_214_n2067) );
  INV_X1 DP_mult_214_U1824 ( .A(DP_mult_214_n2067), .ZN(DP_mult_214_n2070) );
  XNOR2_X1 DP_mult_214_U1823 ( .A(DP_coeff_ret0[21]), .B(DP_coeff_ret0[22]), 
        .ZN(DP_mult_214_n2069) );
  XNOR2_X1 DP_mult_214_U1822 ( .A(DP_coeff_ret0[22]), .B(DP_mult_214_n1611), 
        .ZN(DP_mult_214_n2068) );
  NAND3_X1 DP_mult_214_U1821 ( .A1(DP_mult_214_n2067), .A2(DP_mult_214_n2068), 
        .A3(DP_mult_214_n2069), .ZN(DP_mult_214_n1629) );
  INV_X1 DP_mult_214_U1820 ( .A(DP_sw0_21_), .ZN(DP_mult_214_n1643) );
  OAI22_X1 DP_mult_214_U1819 ( .A1(DP_mult_214_n1544), .A2(DP_mult_214_n1618), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1643), .ZN(DP_mult_214_n2066)
         );
  AOI221_X1 DP_mult_214_U1818 ( .B1(DP_sw0_22_), .B2(DP_mult_214_n1560), .C1(
        DP_mult_214_n1375), .C2(DP_mult_214_n1547), .A(DP_mult_214_n2066), 
        .ZN(DP_mult_214_n2065) );
  XOR2_X1 DP_mult_214_U1817 ( .A(DP_mult_214_n1611), .B(DP_mult_214_n2065), 
        .Z(DP_mult_214_n1627) );
  INV_X1 DP_mult_214_U1816 ( .A(DP_mult_214_n1627), .ZN(DP_mult_214_n351) );
  INV_X1 DP_mult_214_U1815 ( .A(DP_mult_214_n356), .ZN(DP_mult_214_n360) );
  OAI22_X1 DP_mult_214_U1814 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1712), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1713), .ZN(DP_mult_214_n2064)
         );
  AOI221_X1 DP_mult_214_U1813 ( .B1(DP_sw0_17_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_16_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2064), .ZN(
        DP_mult_214_n2063) );
  XOR2_X1 DP_mult_214_U1812 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2063), 
        .Z(DP_mult_214_n374) );
  INV_X1 DP_mult_214_U1811 ( .A(DP_mult_214_n374), .ZN(DP_mult_214_n368) );
  INV_X1 DP_mult_214_U1810 ( .A(DP_mult_214_n387), .ZN(DP_mult_214_n395) );
  OAI22_X1 DP_mult_214_U1809 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1688), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1689), .ZN(DP_mult_214_n2062)
         );
  AOI221_X1 DP_mult_214_U1808 ( .B1(DP_sw0_11_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_10_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2062), .ZN(
        DP_mult_214_n2061) );
  XOR2_X1 DP_mult_214_U1807 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2061), 
        .Z(DP_mult_214_n421) );
  INV_X1 DP_mult_214_U1806 ( .A(DP_mult_214_n421), .ZN(DP_mult_214_n411) );
  OAI22_X1 DP_mult_214_U1805 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1676), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1677), .ZN(DP_mult_214_n2060)
         );
  AOI221_X1 DP_mult_214_U1804 ( .B1(DP_sw0_8_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_7_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2060), .ZN(
        DP_mult_214_n2059) );
  XOR2_X1 DP_mult_214_U1803 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2059), 
        .Z(DP_mult_214_n454) );
  INV_X1 DP_mult_214_U1802 ( .A(DP_mult_214_n454), .ZN(DP_mult_214_n442) );
  OAI21_X1 DP_mult_214_U1801 ( .B1(DP_mult_214_n1561), .B2(DP_mult_214_n1563), 
        .A(DP_mult_214_n1615), .ZN(DP_mult_214_n2058) );
  OAI221_X1 DP_mult_214_U1800 ( .B1(DP_mult_214_n1618), .B2(DP_mult_214_n1639), 
        .C1(DP_mult_214_n1619), .C2(DP_mult_214_n1564), .A(DP_mult_214_n2058), 
        .ZN(DP_mult_214_n2057) );
  XOR2_X1 DP_mult_214_U1799 ( .A(DP_mult_214_n2057), .B(DP_mult_214_n1742), 
        .Z(DP_mult_214_n2056) );
  NOR2_X1 DP_mult_214_U1798 ( .A1(DP_mult_214_n2056), .A2(DP_mult_214_n519), 
        .ZN(DP_mult_214_n493) );
  INV_X1 DP_mult_214_U1797 ( .A(DP_mult_214_n493), .ZN(DP_mult_214_n479) );
  XNOR2_X1 DP_mult_214_U1796 ( .A(DP_mult_214_n519), .B(DP_mult_214_n2056), 
        .ZN(DP_mult_214_n506) );
  INV_X1 DP_mult_214_U1795 ( .A(DP_sw0_20_), .ZN(DP_mult_214_n1640) );
  OAI22_X1 DP_mult_214_U1794 ( .A1(DP_mult_214_n1556), .A2(DP_mult_214_n1640), 
        .B1(DP_mult_214_n1552), .B2(DP_mult_214_n1643), .ZN(DP_mult_214_n2055)
         );
  AOI221_X1 DP_mult_214_U1793 ( .B1(DP_sw0_22_), .B2(DP_mult_214_n1559), .C1(
        DP_mult_214_n1376), .C2(DP_mult_214_n1547), .A(DP_mult_214_n2055), 
        .ZN(DP_mult_214_n2054) );
  XNOR2_X1 DP_mult_214_U1792 ( .A(DP_coeff_ret0[23]), .B(DP_mult_214_n2054), 
        .ZN(DP_mult_214_n729) );
  OAI22_X1 DP_mult_214_U1791 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1728), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1729), .ZN(DP_mult_214_n2053)
         );
  AOI221_X1 DP_mult_214_U1790 ( .B1(DP_sw0_21_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_20_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2053), .ZN(
        DP_mult_214_n2052) );
  XNOR2_X1 DP_mult_214_U1789 ( .A(DP_coeff_ret0[23]), .B(DP_mult_214_n2052), 
        .ZN(DP_mult_214_n730) );
  OAI22_X1 DP_mult_214_U1788 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1724), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1725), .ZN(DP_mult_214_n2051)
         );
  AOI221_X1 DP_mult_214_U1787 ( .B1(DP_sw0_20_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_19_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2051), .ZN(
        DP_mult_214_n2050) );
  XNOR2_X1 DP_mult_214_U1786 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2050), 
        .ZN(DP_mult_214_n731) );
  OAI22_X1 DP_mult_214_U1785 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1720), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1721), .ZN(DP_mult_214_n2049)
         );
  AOI221_X1 DP_mult_214_U1784 ( .B1(DP_sw0_19_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_18_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2049), .ZN(
        DP_mult_214_n2048) );
  XNOR2_X1 DP_mult_214_U1783 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2048), 
        .ZN(DP_mult_214_n732) );
  OAI22_X1 DP_mult_214_U1782 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1716), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1717), .ZN(DP_mult_214_n2047)
         );
  AOI221_X1 DP_mult_214_U1781 ( .B1(DP_sw0_18_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_17_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2047), .ZN(
        DP_mult_214_n2046) );
  XNOR2_X1 DP_mult_214_U1780 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2046), 
        .ZN(DP_mult_214_n733) );
  OAI22_X1 DP_mult_214_U1779 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1708), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1709), .ZN(DP_mult_214_n2045)
         );
  AOI221_X1 DP_mult_214_U1778 ( .B1(DP_sw0_16_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_15_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2045), .ZN(
        DP_mult_214_n2044) );
  XNOR2_X1 DP_mult_214_U1777 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2044), 
        .ZN(DP_mult_214_n734) );
  OAI22_X1 DP_mult_214_U1776 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1704), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1705), .ZN(DP_mult_214_n2043)
         );
  AOI221_X1 DP_mult_214_U1775 ( .B1(DP_sw0_15_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_14_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2043), .ZN(
        DP_mult_214_n2042) );
  XNOR2_X1 DP_mult_214_U1774 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2042), 
        .ZN(DP_mult_214_n735) );
  OAI22_X1 DP_mult_214_U1773 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1700), 
        .B1(DP_mult_214_n1556), .B2(DP_mult_214_n1701), .ZN(DP_mult_214_n2041)
         );
  AOI221_X1 DP_mult_214_U1772 ( .B1(DP_sw0_14_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_13_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2041), .ZN(
        DP_mult_214_n2040) );
  XNOR2_X1 DP_mult_214_U1771 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2040), 
        .ZN(DP_mult_214_n736) );
  OAI22_X1 DP_mult_214_U1770 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1696), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1697), .ZN(DP_mult_214_n2039)
         );
  AOI221_X1 DP_mult_214_U1769 ( .B1(DP_sw0_13_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_12_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2039), .ZN(
        DP_mult_214_n2038) );
  XNOR2_X1 DP_mult_214_U1768 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2038), 
        .ZN(DP_mult_214_n737) );
  OAI22_X1 DP_mult_214_U1767 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1692), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1693), .ZN(DP_mult_214_n2037)
         );
  AOI221_X1 DP_mult_214_U1766 ( .B1(DP_sw0_12_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_11_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2037), .ZN(
        DP_mult_214_n2036) );
  XNOR2_X1 DP_mult_214_U1765 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2036), 
        .ZN(DP_mult_214_n738) );
  OAI22_X1 DP_mult_214_U1764 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1684), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1685), .ZN(DP_mult_214_n2035)
         );
  AOI221_X1 DP_mult_214_U1763 ( .B1(DP_sw0_10_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_9_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2035), .ZN(
        DP_mult_214_n2034) );
  XNOR2_X1 DP_mult_214_U1762 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2034), 
        .ZN(DP_mult_214_n739) );
  OAI22_X1 DP_mult_214_U1761 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1680), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1681), .ZN(DP_mult_214_n2033)
         );
  AOI221_X1 DP_mult_214_U1760 ( .B1(DP_sw0_9_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_8_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2033), .ZN(
        DP_mult_214_n2032) );
  XNOR2_X1 DP_mult_214_U1759 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2032), 
        .ZN(DP_mult_214_n740) );
  OAI22_X1 DP_mult_214_U1758 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1672), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1673), .ZN(DP_mult_214_n2031)
         );
  AOI221_X1 DP_mult_214_U1757 ( .B1(DP_sw0_7_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_6_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2031), .ZN(
        DP_mult_214_n2030) );
  XNOR2_X1 DP_mult_214_U1756 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2030), 
        .ZN(DP_mult_214_n741) );
  OAI22_X1 DP_mult_214_U1755 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1668), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1669), .ZN(DP_mult_214_n2029)
         );
  AOI221_X1 DP_mult_214_U1754 ( .B1(DP_sw0_6_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_5_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2029), .ZN(
        DP_mult_214_n2028) );
  XNOR2_X1 DP_mult_214_U1753 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2028), 
        .ZN(DP_mult_214_n742) );
  OAI22_X1 DP_mult_214_U1752 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1664), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1665), .ZN(DP_mult_214_n2027)
         );
  AOI221_X1 DP_mult_214_U1751 ( .B1(DP_sw0_5_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_4_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2027), .ZN(
        DP_mult_214_n2026) );
  XNOR2_X1 DP_mult_214_U1750 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2026), 
        .ZN(DP_mult_214_n743) );
  OAI22_X1 DP_mult_214_U1749 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1660), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1661), .ZN(DP_mult_214_n2025)
         );
  AOI221_X1 DP_mult_214_U1748 ( .B1(DP_sw0_4_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_3_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2025), .ZN(
        DP_mult_214_n2024) );
  XNOR2_X1 DP_mult_214_U1747 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2024), 
        .ZN(DP_mult_214_n744) );
  OAI22_X1 DP_mult_214_U1746 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1657), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1649), .ZN(DP_mult_214_n2023)
         );
  AOI221_X1 DP_mult_214_U1745 ( .B1(DP_sw0_3_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_2_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2023), .ZN(
        DP_mult_214_n2022) );
  XNOR2_X1 DP_mult_214_U1744 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2022), 
        .ZN(DP_mult_214_n745) );
  INV_X1 DP_mult_214_U1743 ( .A(DP_mult_214_n1396), .ZN(DP_mult_214_n1653) );
  INV_X1 DP_mult_214_U1742 ( .A(DP_sw0_0_), .ZN(DP_mult_214_n1647) );
  OAI22_X1 DP_mult_214_U1741 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1653), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1567), .ZN(DP_mult_214_n2021)
         );
  AOI221_X1 DP_mult_214_U1740 ( .B1(DP_sw0_2_), .B2(DP_mult_214_n1559), .C1(
        DP_sw0_1_), .C2(DP_mult_214_n1560), .A(DP_mult_214_n2021), .ZN(
        DP_mult_214_n2020) );
  XNOR2_X1 DP_mult_214_U1739 ( .A(DP_mult_214_n1610), .B(DP_mult_214_n2020), 
        .ZN(DP_mult_214_n746) );
  OAI222_X1 DP_mult_214_U1738 ( .A1(DP_mult_214_n1544), .A2(DP_mult_214_n1649), 
        .B1(DP_mult_214_n1552), .B2(DP_mult_214_n1566), .C1(DP_mult_214_n1558), 
        .C2(DP_mult_214_n1650), .ZN(DP_mult_214_n2019) );
  XNOR2_X1 DP_mult_214_U1737 ( .A(DP_mult_214_n2019), .B(DP_mult_214_n1611), 
        .ZN(DP_mult_214_n747) );
  OAI22_X1 DP_mult_214_U1736 ( .A1(DP_mult_214_n1544), .A2(DP_mult_214_n1567), 
        .B1(DP_mult_214_n1558), .B2(DP_mult_214_n1567), .ZN(DP_mult_214_n2018)
         );
  XNOR2_X1 DP_mult_214_U1735 ( .A(DP_mult_214_n2018), .B(DP_mult_214_n1611), 
        .ZN(DP_mult_214_n748) );
  XOR2_X1 DP_mult_214_U1734 ( .A(DP_coeff_ret0[18]), .B(DP_mult_214_n1607), 
        .Z(DP_mult_214_n2017) );
  XOR2_X1 DP_mult_214_U1733 ( .A(DP_coeff_ret0[19]), .B(DP_mult_214_n1608), 
        .Z(DP_mult_214_n2016) );
  XNOR2_X1 DP_mult_214_U1732 ( .A(DP_coeff_ret0[18]), .B(DP_coeff_ret0[19]), 
        .ZN(DP_mult_214_n2015) );
  NAND3_X1 DP_mult_214_U1731 ( .A1(DP_mult_214_n2017), .A2(DP_mult_214_n2016), 
        .A3(DP_mult_214_n2015), .ZN(DP_mult_214_n1967) );
  INV_X1 DP_mult_214_U1730 ( .A(DP_mult_214_n2017), .ZN(DP_mult_214_n2014) );
  OAI21_X1 DP_mult_214_U1729 ( .B1(DP_mult_214_n1594), .B2(DP_mult_214_n1595), 
        .A(DP_mult_214_n1615), .ZN(DP_mult_214_n2013) );
  OAI221_X1 DP_mult_214_U1728 ( .B1(DP_mult_214_n1617), .B2(DP_mult_214_n1597), 
        .C1(DP_mult_214_n1619), .C2(DP_mult_214_n1593), .A(DP_mult_214_n2013), 
        .ZN(DP_mult_214_n2012) );
  XNOR2_X1 DP_mult_214_U1727 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n2012), 
        .ZN(DP_mult_214_n749) );
  INV_X1 DP_mult_214_U1726 ( .A(DP_mult_214_n1374), .ZN(DP_mult_214_n1633) );
  INV_X1 DP_mult_214_U1725 ( .A(DP_sw0_22_), .ZN(DP_mult_214_n1634) );
  OAI22_X1 DP_mult_214_U1724 ( .A1(DP_mult_214_n1633), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1634), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n2011)
         );
  AOI221_X1 DP_mult_214_U1723 ( .B1(DP_mult_214_n1594), .B2(DP_mult_214_n1614), 
        .C1(DP_mult_214_n1595), .C2(DP_mult_214_n1615), .A(DP_mult_214_n2011), 
        .ZN(DP_mult_214_n2010) );
  XNOR2_X1 DP_mult_214_U1722 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n2010), 
        .ZN(DP_mult_214_n750) );
  OAI22_X1 DP_mult_214_U1721 ( .A1(DP_mult_214_n1620), .A2(DP_mult_214_n1543), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n2009)
         );
  AOI221_X1 DP_mult_214_U1720 ( .B1(DP_mult_214_n1595), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1545), .C2(DP_mult_214_n1375), .A(DP_mult_214_n2009), 
        .ZN(DP_mult_214_n2008) );
  XNOR2_X1 DP_mult_214_U1719 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n2008), 
        .ZN(DP_mult_214_n751) );
  OAI22_X1 DP_mult_214_U1718 ( .A1(DP_mult_214_n1640), .A2(DP_mult_214_n1597), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1555), .ZN(DP_mult_214_n2007)
         );
  AOI221_X1 DP_mult_214_U1717 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1545), .C2(DP_mult_214_n1376), .A(DP_mult_214_n2007), 
        .ZN(DP_mult_214_n2006) );
  XNOR2_X1 DP_mult_214_U1716 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n2006), 
        .ZN(DP_mult_214_n752) );
  OAI22_X1 DP_mult_214_U1715 ( .A1(DP_mult_214_n1728), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1729), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n2005)
         );
  AOI221_X1 DP_mult_214_U1714 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_21_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_20_), .A(DP_mult_214_n2005), .ZN(
        DP_mult_214_n2004) );
  XNOR2_X1 DP_mult_214_U1713 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n2004), 
        .ZN(DP_mult_214_n753) );
  OAI22_X1 DP_mult_214_U1712 ( .A1(DP_mult_214_n1724), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1725), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n2003)
         );
  AOI221_X1 DP_mult_214_U1711 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_20_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_19_), .A(DP_mult_214_n2003), .ZN(
        DP_mult_214_n2002) );
  XNOR2_X1 DP_mult_214_U1710 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n2002), 
        .ZN(DP_mult_214_n754) );
  OAI22_X1 DP_mult_214_U1709 ( .A1(DP_mult_214_n1720), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1721), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n2001)
         );
  AOI221_X1 DP_mult_214_U1708 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_19_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_18_), .A(DP_mult_214_n2001), .ZN(
        DP_mult_214_n2000) );
  XNOR2_X1 DP_mult_214_U1707 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n2000), 
        .ZN(DP_mult_214_n755) );
  OAI22_X1 DP_mult_214_U1706 ( .A1(DP_mult_214_n1716), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1717), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n1999)
         );
  AOI221_X1 DP_mult_214_U1705 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_18_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_17_), .A(DP_mult_214_n1999), .ZN(
        DP_mult_214_n1998) );
  XNOR2_X1 DP_mult_214_U1704 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n1998), 
        .ZN(DP_mult_214_n756) );
  OAI22_X1 DP_mult_214_U1703 ( .A1(DP_mult_214_n1712), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1713), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n1997)
         );
  AOI221_X1 DP_mult_214_U1702 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_17_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_16_), .A(DP_mult_214_n1997), .ZN(
        DP_mult_214_n1996) );
  XNOR2_X1 DP_mult_214_U1701 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n1996), 
        .ZN(DP_mult_214_n757) );
  OAI22_X1 DP_mult_214_U1700 ( .A1(DP_mult_214_n1708), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1709), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n1995)
         );
  AOI221_X1 DP_mult_214_U1699 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_16_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_15_), .A(DP_mult_214_n1995), .ZN(
        DP_mult_214_n1994) );
  XNOR2_X1 DP_mult_214_U1698 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n1994), 
        .ZN(DP_mult_214_n758) );
  OAI22_X1 DP_mult_214_U1697 ( .A1(DP_mult_214_n1704), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1705), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n1993)
         );
  AOI221_X1 DP_mult_214_U1696 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_15_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_14_), .A(DP_mult_214_n1993), .ZN(
        DP_mult_214_n1992) );
  XNOR2_X1 DP_mult_214_U1695 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n1992), 
        .ZN(DP_mult_214_n759) );
  OAI22_X1 DP_mult_214_U1694 ( .A1(DP_mult_214_n1700), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1701), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n1991)
         );
  AOI221_X1 DP_mult_214_U1693 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_14_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_13_), .A(DP_mult_214_n1991), .ZN(
        DP_mult_214_n1990) );
  XNOR2_X1 DP_mult_214_U1692 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n1990), 
        .ZN(DP_mult_214_n760) );
  OAI22_X1 DP_mult_214_U1691 ( .A1(DP_mult_214_n1696), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1697), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n1989)
         );
  AOI221_X1 DP_mult_214_U1690 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_13_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_12_), .A(DP_mult_214_n1989), .ZN(
        DP_mult_214_n1988) );
  XNOR2_X1 DP_mult_214_U1689 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n1988), 
        .ZN(DP_mult_214_n761) );
  OAI22_X1 DP_mult_214_U1688 ( .A1(DP_mult_214_n1692), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1693), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1987)
         );
  AOI221_X1 DP_mult_214_U1687 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_12_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_11_), .A(DP_mult_214_n1987), .ZN(
        DP_mult_214_n1986) );
  XNOR2_X1 DP_mult_214_U1686 ( .A(DP_mult_214_n1609), .B(DP_mult_214_n1986), 
        .ZN(DP_mult_214_n762) );
  OAI22_X1 DP_mult_214_U1685 ( .A1(DP_mult_214_n1688), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1689), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1985)
         );
  AOI221_X1 DP_mult_214_U1684 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_11_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_10_), .A(DP_mult_214_n1985), .ZN(
        DP_mult_214_n1984) );
  XNOR2_X1 DP_mult_214_U1683 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1984), 
        .ZN(DP_mult_214_n763) );
  OAI22_X1 DP_mult_214_U1682 ( .A1(DP_mult_214_n1684), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1685), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1983)
         );
  AOI221_X1 DP_mult_214_U1681 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_10_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_9_), .A(DP_mult_214_n1983), .ZN(
        DP_mult_214_n1982) );
  XNOR2_X1 DP_mult_214_U1680 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1982), 
        .ZN(DP_mult_214_n764) );
  OAI22_X1 DP_mult_214_U1679 ( .A1(DP_mult_214_n1680), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1681), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1981)
         );
  AOI221_X1 DP_mult_214_U1678 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_9_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_8_), .A(DP_mult_214_n1981), .ZN(
        DP_mult_214_n1980) );
  XNOR2_X1 DP_mult_214_U1677 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1980), 
        .ZN(DP_mult_214_n765) );
  OAI22_X1 DP_mult_214_U1676 ( .A1(DP_mult_214_n1676), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1677), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1979)
         );
  AOI221_X1 DP_mult_214_U1675 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_8_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_7_), .A(DP_mult_214_n1979), .ZN(
        DP_mult_214_n1978) );
  XNOR2_X1 DP_mult_214_U1674 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1978), 
        .ZN(DP_mult_214_n766) );
  OAI22_X1 DP_mult_214_U1673 ( .A1(DP_mult_214_n1672), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1673), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1977)
         );
  AOI221_X1 DP_mult_214_U1672 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_7_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_6_), .A(DP_mult_214_n1977), .ZN(
        DP_mult_214_n1976) );
  XNOR2_X1 DP_mult_214_U1671 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1976), 
        .ZN(DP_mult_214_n767) );
  OAI22_X1 DP_mult_214_U1670 ( .A1(DP_mult_214_n1668), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1669), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1975)
         );
  AOI221_X1 DP_mult_214_U1669 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_6_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_5_), .A(DP_mult_214_n1975), .ZN(
        DP_mult_214_n1974) );
  XNOR2_X1 DP_mult_214_U1668 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1974), 
        .ZN(DP_mult_214_n768) );
  OAI22_X1 DP_mult_214_U1667 ( .A1(DP_mult_214_n1664), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1665), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1973)
         );
  AOI221_X1 DP_mult_214_U1666 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_5_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_4_), .A(DP_mult_214_n1973), .ZN(
        DP_mult_214_n1972) );
  XNOR2_X1 DP_mult_214_U1665 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1972), 
        .ZN(DP_mult_214_n769) );
  OAI22_X1 DP_mult_214_U1664 ( .A1(DP_mult_214_n1660), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1661), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1971)
         );
  AOI221_X1 DP_mult_214_U1663 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_4_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_3_), .A(DP_mult_214_n1971), .ZN(
        DP_mult_214_n1970) );
  XNOR2_X1 DP_mult_214_U1662 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1970), 
        .ZN(DP_mult_214_n770) );
  OAI22_X1 DP_mult_214_U1661 ( .A1(DP_mult_214_n1657), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1649), .B2(DP_mult_214_n1597), .ZN(DP_mult_214_n1969)
         );
  AOI221_X1 DP_mult_214_U1660 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_3_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_2_), .A(DP_mult_214_n1969), .ZN(
        DP_mult_214_n1968) );
  XNOR2_X1 DP_mult_214_U1659 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1968), 
        .ZN(DP_mult_214_n771) );
  OAI22_X1 DP_mult_214_U1658 ( .A1(DP_mult_214_n1653), .A2(DP_mult_214_n1593), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1596), .ZN(DP_mult_214_n1966)
         );
  AOI221_X1 DP_mult_214_U1657 ( .B1(DP_mult_214_n1594), .B2(DP_sw0_2_), .C1(
        DP_mult_214_n1595), .C2(DP_sw0_1_), .A(DP_mult_214_n1966), .ZN(
        DP_mult_214_n1965) );
  XNOR2_X1 DP_mult_214_U1656 ( .A(DP_mult_214_n1608), .B(DP_mult_214_n1965), 
        .ZN(DP_mult_214_n772) );
  OAI222_X1 DP_mult_214_U1655 ( .A1(DP_mult_214_n1649), .A2(DP_mult_214_n1543), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1555), .C1(DP_mult_214_n1650), 
        .C2(DP_mult_214_n1593), .ZN(DP_mult_214_n1964) );
  XOR2_X1 DP_mult_214_U1654 ( .A(DP_mult_214_n1964), .B(DP_mult_214_n1608), 
        .Z(DP_mult_214_n773) );
  OAI22_X1 DP_mult_214_U1653 ( .A1(DP_mult_214_n1565), .A2(DP_mult_214_n1543), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1593), .ZN(DP_mult_214_n1963)
         );
  XOR2_X1 DP_mult_214_U1652 ( .A(DP_mult_214_n1963), .B(DP_mult_214_n1608), 
        .Z(DP_mult_214_n774) );
  XOR2_X1 DP_mult_214_U1651 ( .A(DP_coeff_ret0[15]), .B(DP_mult_214_n1605), 
        .Z(DP_mult_214_n1962) );
  XNOR2_X1 DP_mult_214_U1650 ( .A(DP_coeff_ret0[16]), .B(DP_mult_214_n1607), 
        .ZN(DP_mult_214_n1961) );
  XNOR2_X1 DP_mult_214_U1649 ( .A(DP_coeff_ret0[15]), .B(DP_coeff_ret0[16]), 
        .ZN(DP_mult_214_n1960) );
  NAND3_X1 DP_mult_214_U1648 ( .A1(DP_mult_214_n1962), .A2(DP_mult_214_n1961), 
        .A3(DP_mult_214_n1960), .ZN(DP_mult_214_n1912) );
  INV_X1 DP_mult_214_U1647 ( .A(DP_mult_214_n1962), .ZN(DP_mult_214_n1959) );
  OAI21_X1 DP_mult_214_U1646 ( .B1(DP_mult_214_n1589), .B2(DP_mult_214_n1590), 
        .A(DP_mult_214_n1615), .ZN(DP_mult_214_n1958) );
  OAI221_X1 DP_mult_214_U1645 ( .B1(DP_mult_214_n1618), .B2(DP_mult_214_n1592), 
        .C1(DP_mult_214_n1617), .C2(DP_mult_214_n1588), .A(DP_mult_214_n1958), 
        .ZN(DP_mult_214_n1957) );
  XNOR2_X1 DP_mult_214_U1644 ( .A(DP_coeff_ret0[17]), .B(DP_mult_214_n1957), 
        .ZN(DP_mult_214_n775) );
  OAI22_X1 DP_mult_214_U1643 ( .A1(DP_mult_214_n1633), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1634), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1956)
         );
  AOI221_X1 DP_mult_214_U1642 ( .B1(DP_mult_214_n1589), .B2(DP_mult_214_n1613), 
        .C1(DP_mult_214_n1590), .C2(DP_mult_214_n1615), .A(DP_mult_214_n1956), 
        .ZN(DP_mult_214_n1955) );
  XNOR2_X1 DP_mult_214_U1641 ( .A(DP_coeff_ret0[17]), .B(DP_mult_214_n1955), 
        .ZN(DP_mult_214_n776) );
  OAI22_X1 DP_mult_214_U1640 ( .A1(DP_mult_214_n1620), .A2(DP_mult_214_n1549), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1954)
         );
  AOI221_X1 DP_mult_214_U1639 ( .B1(DP_mult_214_n1590), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1546), .C2(DP_mult_214_n1375), .A(DP_mult_214_n1954), 
        .ZN(DP_mult_214_n1953) );
  XNOR2_X1 DP_mult_214_U1638 ( .A(DP_coeff_ret0[17]), .B(DP_mult_214_n1953), 
        .ZN(DP_mult_214_n777) );
  OAI22_X1 DP_mult_214_U1637 ( .A1(DP_mult_214_n1640), .A2(DP_mult_214_n1592), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1554), .ZN(DP_mult_214_n1952)
         );
  AOI221_X1 DP_mult_214_U1636 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1546), .C2(DP_mult_214_n1376), .A(DP_mult_214_n1952), 
        .ZN(DP_mult_214_n1951) );
  XNOR2_X1 DP_mult_214_U1635 ( .A(DP_coeff_ret0[17]), .B(DP_mult_214_n1951), 
        .ZN(DP_mult_214_n778) );
  OAI22_X1 DP_mult_214_U1634 ( .A1(DP_mult_214_n1728), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1729), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1950)
         );
  AOI221_X1 DP_mult_214_U1633 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_21_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_20_), .A(DP_mult_214_n1950), .ZN(
        DP_mult_214_n1949) );
  XNOR2_X1 DP_mult_214_U1632 ( .A(DP_coeff_ret0[17]), .B(DP_mult_214_n1949), 
        .ZN(DP_mult_214_n779) );
  OAI22_X1 DP_mult_214_U1631 ( .A1(DP_mult_214_n1724), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1725), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1948)
         );
  AOI221_X1 DP_mult_214_U1630 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_20_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_19_), .A(DP_mult_214_n1948), .ZN(
        DP_mult_214_n1947) );
  XNOR2_X1 DP_mult_214_U1629 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1947), 
        .ZN(DP_mult_214_n780) );
  OAI22_X1 DP_mult_214_U1628 ( .A1(DP_mult_214_n1720), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1721), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1946)
         );
  AOI221_X1 DP_mult_214_U1627 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_19_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_18_), .A(DP_mult_214_n1946), .ZN(
        DP_mult_214_n1945) );
  XNOR2_X1 DP_mult_214_U1626 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1945), 
        .ZN(DP_mult_214_n781) );
  OAI22_X1 DP_mult_214_U1625 ( .A1(DP_mult_214_n1716), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1717), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1944)
         );
  AOI221_X1 DP_mult_214_U1624 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_18_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_17_), .A(DP_mult_214_n1944), .ZN(
        DP_mult_214_n1943) );
  XNOR2_X1 DP_mult_214_U1623 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1943), 
        .ZN(DP_mult_214_n782) );
  OAI22_X1 DP_mult_214_U1622 ( .A1(DP_mult_214_n1712), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1713), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1942)
         );
  AOI221_X1 DP_mult_214_U1621 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_17_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_16_), .A(DP_mult_214_n1942), .ZN(
        DP_mult_214_n1941) );
  XNOR2_X1 DP_mult_214_U1620 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1941), 
        .ZN(DP_mult_214_n783) );
  OAI22_X1 DP_mult_214_U1619 ( .A1(DP_mult_214_n1708), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1709), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1940)
         );
  AOI221_X1 DP_mult_214_U1618 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_16_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_15_), .A(DP_mult_214_n1940), .ZN(
        DP_mult_214_n1939) );
  XNOR2_X1 DP_mult_214_U1617 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1939), 
        .ZN(DP_mult_214_n784) );
  OAI22_X1 DP_mult_214_U1616 ( .A1(DP_mult_214_n1704), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1705), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1938)
         );
  AOI221_X1 DP_mult_214_U1615 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_15_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_14_), .A(DP_mult_214_n1938), .ZN(
        DP_mult_214_n1937) );
  XNOR2_X1 DP_mult_214_U1614 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1937), 
        .ZN(DP_mult_214_n785) );
  OAI22_X1 DP_mult_214_U1613 ( .A1(DP_mult_214_n1700), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1701), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1936)
         );
  AOI221_X1 DP_mult_214_U1612 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_14_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_13_), .A(DP_mult_214_n1936), .ZN(
        DP_mult_214_n1935) );
  XNOR2_X1 DP_mult_214_U1611 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1935), 
        .ZN(DP_mult_214_n786) );
  OAI22_X1 DP_mult_214_U1610 ( .A1(DP_mult_214_n1696), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1697), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1934)
         );
  AOI221_X1 DP_mult_214_U1609 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_13_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_12_), .A(DP_mult_214_n1934), .ZN(
        DP_mult_214_n1933) );
  XNOR2_X1 DP_mult_214_U1608 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1933), 
        .ZN(DP_mult_214_n787) );
  OAI22_X1 DP_mult_214_U1607 ( .A1(DP_mult_214_n1692), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1693), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1932)
         );
  AOI221_X1 DP_mult_214_U1606 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_12_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_11_), .A(DP_mult_214_n1932), .ZN(
        DP_mult_214_n1931) );
  XNOR2_X1 DP_mult_214_U1605 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1931), 
        .ZN(DP_mult_214_n788) );
  OAI22_X1 DP_mult_214_U1604 ( .A1(DP_mult_214_n1688), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1689), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1930)
         );
  AOI221_X1 DP_mult_214_U1603 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_11_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_10_), .A(DP_mult_214_n1930), .ZN(
        DP_mult_214_n1929) );
  XNOR2_X1 DP_mult_214_U1602 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1929), 
        .ZN(DP_mult_214_n789) );
  OAI22_X1 DP_mult_214_U1601 ( .A1(DP_mult_214_n1684), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1685), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1928)
         );
  AOI221_X1 DP_mult_214_U1600 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_10_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_9_), .A(DP_mult_214_n1928), .ZN(
        DP_mult_214_n1927) );
  XNOR2_X1 DP_mult_214_U1599 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1927), 
        .ZN(DP_mult_214_n790) );
  OAI22_X1 DP_mult_214_U1598 ( .A1(DP_mult_214_n1680), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1681), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1926)
         );
  AOI221_X1 DP_mult_214_U1597 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_9_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_8_), .A(DP_mult_214_n1926), .ZN(
        DP_mult_214_n1925) );
  XNOR2_X1 DP_mult_214_U1596 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1925), 
        .ZN(DP_mult_214_n791) );
  OAI22_X1 DP_mult_214_U1595 ( .A1(DP_mult_214_n1676), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1677), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1924)
         );
  AOI221_X1 DP_mult_214_U1594 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_8_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_7_), .A(DP_mult_214_n1924), .ZN(
        DP_mult_214_n1923) );
  XNOR2_X1 DP_mult_214_U1593 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1923), 
        .ZN(DP_mult_214_n792) );
  OAI22_X1 DP_mult_214_U1592 ( .A1(DP_mult_214_n1672), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1673), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1922)
         );
  AOI221_X1 DP_mult_214_U1591 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_7_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_6_), .A(DP_mult_214_n1922), .ZN(
        DP_mult_214_n1921) );
  XNOR2_X1 DP_mult_214_U1590 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1921), 
        .ZN(DP_mult_214_n793) );
  OAI22_X1 DP_mult_214_U1589 ( .A1(DP_mult_214_n1668), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1669), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1920)
         );
  AOI221_X1 DP_mult_214_U1588 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_6_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_5_), .A(DP_mult_214_n1920), .ZN(
        DP_mult_214_n1919) );
  XNOR2_X1 DP_mult_214_U1587 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1919), 
        .ZN(DP_mult_214_n794) );
  OAI22_X1 DP_mult_214_U1586 ( .A1(DP_mult_214_n1664), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1665), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1918)
         );
  AOI221_X1 DP_mult_214_U1585 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_5_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_4_), .A(DP_mult_214_n1918), .ZN(
        DP_mult_214_n1917) );
  XNOR2_X1 DP_mult_214_U1584 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1917), 
        .ZN(DP_mult_214_n795) );
  OAI22_X1 DP_mult_214_U1583 ( .A1(DP_mult_214_n1660), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1661), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1916)
         );
  AOI221_X1 DP_mult_214_U1582 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_4_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_3_), .A(DP_mult_214_n1916), .ZN(
        DP_mult_214_n1915) );
  XNOR2_X1 DP_mult_214_U1581 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1915), 
        .ZN(DP_mult_214_n796) );
  OAI22_X1 DP_mult_214_U1580 ( .A1(DP_mult_214_n1657), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1649), .B2(DP_mult_214_n1592), .ZN(DP_mult_214_n1914)
         );
  AOI221_X1 DP_mult_214_U1579 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_3_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_2_), .A(DP_mult_214_n1914), .ZN(
        DP_mult_214_n1913) );
  XNOR2_X1 DP_mult_214_U1578 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1913), 
        .ZN(DP_mult_214_n797) );
  OAI22_X1 DP_mult_214_U1577 ( .A1(DP_mult_214_n1653), .A2(DP_mult_214_n1588), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1591), .ZN(DP_mult_214_n1911)
         );
  AOI221_X1 DP_mult_214_U1576 ( .B1(DP_mult_214_n1589), .B2(DP_sw0_2_), .C1(
        DP_mult_214_n1590), .C2(DP_sw0_1_), .A(DP_mult_214_n1911), .ZN(
        DP_mult_214_n1910) );
  XNOR2_X1 DP_mult_214_U1575 ( .A(DP_mult_214_n1606), .B(DP_mult_214_n1910), 
        .ZN(DP_mult_214_n798) );
  OAI222_X1 DP_mult_214_U1574 ( .A1(DP_mult_214_n1649), .A2(DP_mult_214_n1549), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1554), .C1(DP_mult_214_n1650), 
        .C2(DP_mult_214_n1588), .ZN(DP_mult_214_n1909) );
  XNOR2_X1 DP_mult_214_U1573 ( .A(DP_mult_214_n1909), .B(DP_mult_214_n1607), 
        .ZN(DP_mult_214_n799) );
  OAI22_X1 DP_mult_214_U1572 ( .A1(DP_mult_214_n1565), .A2(DP_mult_214_n1549), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1588), .ZN(DP_mult_214_n1908)
         );
  XNOR2_X1 DP_mult_214_U1571 ( .A(DP_mult_214_n1908), .B(DP_mult_214_n1607), 
        .ZN(DP_mult_214_n800) );
  XOR2_X1 DP_mult_214_U1570 ( .A(DP_coeff_ret0[12]), .B(DP_mult_214_n1603), 
        .Z(DP_mult_214_n1907) );
  XNOR2_X1 DP_mult_214_U1569 ( .A(DP_coeff_ret0[13]), .B(DP_mult_214_n1605), 
        .ZN(DP_mult_214_n1906) );
  XNOR2_X1 DP_mult_214_U1568 ( .A(DP_coeff_ret0[12]), .B(DP_coeff_ret0[13]), 
        .ZN(DP_mult_214_n1905) );
  NAND3_X1 DP_mult_214_U1567 ( .A1(DP_mult_214_n1907), .A2(DP_mult_214_n1906), 
        .A3(DP_mult_214_n1905), .ZN(DP_mult_214_n1857) );
  INV_X1 DP_mult_214_U1566 ( .A(DP_mult_214_n1907), .ZN(DP_mult_214_n1904) );
  OAI21_X1 DP_mult_214_U1565 ( .B1(DP_mult_214_n1584), .B2(DP_mult_214_n1585), 
        .A(DP_mult_214_n1615), .ZN(DP_mult_214_n1903) );
  OAI221_X1 DP_mult_214_U1564 ( .B1(DP_mult_214_n1620), .B2(DP_mult_214_n1587), 
        .C1(DP_mult_214_n1619), .C2(DP_mult_214_n1583), .A(DP_mult_214_n1903), 
        .ZN(DP_mult_214_n1902) );
  XNOR2_X1 DP_mult_214_U1563 ( .A(DP_coeff_ret0[14]), .B(DP_mult_214_n1902), 
        .ZN(DP_mult_214_n801) );
  OAI22_X1 DP_mult_214_U1562 ( .A1(DP_mult_214_n1633), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1634), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1901)
         );
  AOI221_X1 DP_mult_214_U1561 ( .B1(DP_mult_214_n1584), .B2(DP_mult_214_n1615), 
        .C1(DP_mult_214_n1585), .C2(DP_mult_214_n1615), .A(DP_mult_214_n1901), 
        .ZN(DP_mult_214_n1900) );
  XNOR2_X1 DP_mult_214_U1560 ( .A(DP_coeff_ret0[14]), .B(DP_mult_214_n1900), 
        .ZN(DP_mult_214_n802) );
  OAI22_X1 DP_mult_214_U1559 ( .A1(DP_mult_214_n1617), .A2(DP_mult_214_n1548), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1899)
         );
  AOI221_X1 DP_mult_214_U1558 ( .B1(DP_mult_214_n1585), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1551), .C2(DP_mult_214_n1375), .A(DP_mult_214_n1899), 
        .ZN(DP_mult_214_n1898) );
  XNOR2_X1 DP_mult_214_U1557 ( .A(DP_coeff_ret0[14]), .B(DP_mult_214_n1898), 
        .ZN(DP_mult_214_n803) );
  OAI22_X1 DP_mult_214_U1556 ( .A1(DP_mult_214_n1640), .A2(DP_mult_214_n1587), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1553), .ZN(DP_mult_214_n1897)
         );
  AOI221_X1 DP_mult_214_U1555 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1551), .C2(DP_mult_214_n1376), .A(DP_mult_214_n1897), 
        .ZN(DP_mult_214_n1896) );
  XNOR2_X1 DP_mult_214_U1554 ( .A(DP_coeff_ret0[14]), .B(DP_mult_214_n1896), 
        .ZN(DP_mult_214_n804) );
  OAI22_X1 DP_mult_214_U1553 ( .A1(DP_mult_214_n1728), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1729), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1895)
         );
  AOI221_X1 DP_mult_214_U1552 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_21_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_20_), .A(DP_mult_214_n1895), .ZN(
        DP_mult_214_n1894) );
  XNOR2_X1 DP_mult_214_U1551 ( .A(DP_coeff_ret0[14]), .B(DP_mult_214_n1894), 
        .ZN(DP_mult_214_n805) );
  OAI22_X1 DP_mult_214_U1550 ( .A1(DP_mult_214_n1724), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1725), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1893)
         );
  AOI221_X1 DP_mult_214_U1549 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_20_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_19_), .A(DP_mult_214_n1893), .ZN(
        DP_mult_214_n1892) );
  XNOR2_X1 DP_mult_214_U1548 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1892), 
        .ZN(DP_mult_214_n806) );
  OAI22_X1 DP_mult_214_U1547 ( .A1(DP_mult_214_n1720), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1721), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1891)
         );
  AOI221_X1 DP_mult_214_U1546 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_19_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_18_), .A(DP_mult_214_n1891), .ZN(
        DP_mult_214_n1890) );
  XNOR2_X1 DP_mult_214_U1545 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1890), 
        .ZN(DP_mult_214_n807) );
  OAI22_X1 DP_mult_214_U1544 ( .A1(DP_mult_214_n1716), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1717), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1889)
         );
  AOI221_X1 DP_mult_214_U1543 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_18_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_17_), .A(DP_mult_214_n1889), .ZN(
        DP_mult_214_n1888) );
  XNOR2_X1 DP_mult_214_U1542 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1888), 
        .ZN(DP_mult_214_n808) );
  OAI22_X1 DP_mult_214_U1541 ( .A1(DP_mult_214_n1712), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1713), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1887)
         );
  AOI221_X1 DP_mult_214_U1540 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_17_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_16_), .A(DP_mult_214_n1887), .ZN(
        DP_mult_214_n1886) );
  XNOR2_X1 DP_mult_214_U1539 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1886), 
        .ZN(DP_mult_214_n809) );
  OAI22_X1 DP_mult_214_U1538 ( .A1(DP_mult_214_n1708), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1709), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1885)
         );
  AOI221_X1 DP_mult_214_U1537 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_16_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_15_), .A(DP_mult_214_n1885), .ZN(
        DP_mult_214_n1884) );
  XNOR2_X1 DP_mult_214_U1536 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1884), 
        .ZN(DP_mult_214_n810) );
  OAI22_X1 DP_mult_214_U1535 ( .A1(DP_mult_214_n1704), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1705), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1883)
         );
  AOI221_X1 DP_mult_214_U1534 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_15_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_14_), .A(DP_mult_214_n1883), .ZN(
        DP_mult_214_n1882) );
  XNOR2_X1 DP_mult_214_U1533 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1882), 
        .ZN(DP_mult_214_n811) );
  OAI22_X1 DP_mult_214_U1532 ( .A1(DP_mult_214_n1700), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1701), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1881)
         );
  AOI221_X1 DP_mult_214_U1531 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_14_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_13_), .A(DP_mult_214_n1881), .ZN(
        DP_mult_214_n1880) );
  XNOR2_X1 DP_mult_214_U1530 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1880), 
        .ZN(DP_mult_214_n812) );
  OAI22_X1 DP_mult_214_U1529 ( .A1(DP_mult_214_n1696), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1697), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1879)
         );
  AOI221_X1 DP_mult_214_U1528 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_13_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_12_), .A(DP_mult_214_n1879), .ZN(
        DP_mult_214_n1878) );
  XNOR2_X1 DP_mult_214_U1527 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1878), 
        .ZN(DP_mult_214_n813) );
  OAI22_X1 DP_mult_214_U1526 ( .A1(DP_mult_214_n1692), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1693), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1877)
         );
  AOI221_X1 DP_mult_214_U1525 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_12_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_11_), .A(DP_mult_214_n1877), .ZN(
        DP_mult_214_n1876) );
  XNOR2_X1 DP_mult_214_U1524 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1876), 
        .ZN(DP_mult_214_n814) );
  OAI22_X1 DP_mult_214_U1523 ( .A1(DP_mult_214_n1688), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1689), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1875)
         );
  AOI221_X1 DP_mult_214_U1522 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_11_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_10_), .A(DP_mult_214_n1875), .ZN(
        DP_mult_214_n1874) );
  XNOR2_X1 DP_mult_214_U1521 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1874), 
        .ZN(DP_mult_214_n815) );
  OAI22_X1 DP_mult_214_U1520 ( .A1(DP_mult_214_n1684), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1685), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1873)
         );
  AOI221_X1 DP_mult_214_U1519 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_10_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_9_), .A(DP_mult_214_n1873), .ZN(
        DP_mult_214_n1872) );
  XNOR2_X1 DP_mult_214_U1518 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1872), 
        .ZN(DP_mult_214_n816) );
  OAI22_X1 DP_mult_214_U1517 ( .A1(DP_mult_214_n1680), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1681), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1871)
         );
  AOI221_X1 DP_mult_214_U1516 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_9_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_8_), .A(DP_mult_214_n1871), .ZN(
        DP_mult_214_n1870) );
  XNOR2_X1 DP_mult_214_U1515 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1870), 
        .ZN(DP_mult_214_n817) );
  OAI22_X1 DP_mult_214_U1514 ( .A1(DP_mult_214_n1676), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1677), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1869)
         );
  AOI221_X1 DP_mult_214_U1513 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_8_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_7_), .A(DP_mult_214_n1869), .ZN(
        DP_mult_214_n1868) );
  XNOR2_X1 DP_mult_214_U1512 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1868), 
        .ZN(DP_mult_214_n818) );
  OAI22_X1 DP_mult_214_U1511 ( .A1(DP_mult_214_n1672), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1673), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1867)
         );
  AOI221_X1 DP_mult_214_U1510 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_7_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_6_), .A(DP_mult_214_n1867), .ZN(
        DP_mult_214_n1866) );
  XNOR2_X1 DP_mult_214_U1509 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1866), 
        .ZN(DP_mult_214_n819) );
  OAI22_X1 DP_mult_214_U1508 ( .A1(DP_mult_214_n1668), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1669), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1865)
         );
  AOI221_X1 DP_mult_214_U1507 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_6_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_5_), .A(DP_mult_214_n1865), .ZN(
        DP_mult_214_n1864) );
  XNOR2_X1 DP_mult_214_U1506 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1864), 
        .ZN(DP_mult_214_n820) );
  OAI22_X1 DP_mult_214_U1505 ( .A1(DP_mult_214_n1664), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1665), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1863)
         );
  AOI221_X1 DP_mult_214_U1504 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_5_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_4_), .A(DP_mult_214_n1863), .ZN(
        DP_mult_214_n1862) );
  XNOR2_X1 DP_mult_214_U1503 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1862), 
        .ZN(DP_mult_214_n821) );
  OAI22_X1 DP_mult_214_U1502 ( .A1(DP_mult_214_n1660), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1661), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1861)
         );
  AOI221_X1 DP_mult_214_U1501 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_4_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_3_), .A(DP_mult_214_n1861), .ZN(
        DP_mult_214_n1860) );
  XNOR2_X1 DP_mult_214_U1500 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1860), 
        .ZN(DP_mult_214_n822) );
  OAI22_X1 DP_mult_214_U1499 ( .A1(DP_mult_214_n1657), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1649), .B2(DP_mult_214_n1587), .ZN(DP_mult_214_n1859)
         );
  AOI221_X1 DP_mult_214_U1498 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_3_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_2_), .A(DP_mult_214_n1859), .ZN(
        DP_mult_214_n1858) );
  XNOR2_X1 DP_mult_214_U1497 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1858), 
        .ZN(DP_mult_214_n823) );
  OAI22_X1 DP_mult_214_U1496 ( .A1(DP_mult_214_n1653), .A2(DP_mult_214_n1583), 
        .B1(DP_mult_214_n1565), .B2(DP_mult_214_n1586), .ZN(DP_mult_214_n1856)
         );
  AOI221_X1 DP_mult_214_U1495 ( .B1(DP_mult_214_n1584), .B2(DP_sw0_2_), .C1(
        DP_mult_214_n1585), .C2(DP_sw0_1_), .A(DP_mult_214_n1856), .ZN(
        DP_mult_214_n1855) );
  XNOR2_X1 DP_mult_214_U1494 ( .A(DP_mult_214_n1604), .B(DP_mult_214_n1855), 
        .ZN(DP_mult_214_n824) );
  OAI222_X1 DP_mult_214_U1493 ( .A1(DP_mult_214_n1649), .A2(DP_mult_214_n1548), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1553), .C1(DP_mult_214_n1650), 
        .C2(DP_mult_214_n1583), .ZN(DP_mult_214_n1854) );
  XNOR2_X1 DP_mult_214_U1492 ( .A(DP_mult_214_n1854), .B(DP_mult_214_n1605), 
        .ZN(DP_mult_214_n825) );
  OAI22_X1 DP_mult_214_U1491 ( .A1(DP_mult_214_n1565), .A2(DP_mult_214_n1548), 
        .B1(DP_mult_214_n1565), .B2(DP_mult_214_n1583), .ZN(DP_mult_214_n1853)
         );
  XNOR2_X1 DP_mult_214_U1490 ( .A(DP_mult_214_n1853), .B(DP_mult_214_n1605), 
        .ZN(DP_mult_214_n826) );
  XOR2_X1 DP_mult_214_U1489 ( .A(DP_coeff_ret0[9]), .B(DP_mult_214_n1601), .Z(
        DP_mult_214_n1852) );
  XNOR2_X1 DP_mult_214_U1488 ( .A(DP_coeff_ret0[10]), .B(DP_mult_214_n1603), 
        .ZN(DP_mult_214_n1851) );
  XNOR2_X1 DP_mult_214_U1487 ( .A(DP_coeff_ret0[10]), .B(DP_coeff_ret0[9]), 
        .ZN(DP_mult_214_n1850) );
  NAND3_X1 DP_mult_214_U1486 ( .A1(DP_mult_214_n1852), .A2(DP_mult_214_n1851), 
        .A3(DP_mult_214_n1850), .ZN(DP_mult_214_n1802) );
  INV_X1 DP_mult_214_U1485 ( .A(DP_mult_214_n1852), .ZN(DP_mult_214_n1849) );
  OAI21_X1 DP_mult_214_U1484 ( .B1(DP_mult_214_n1579), .B2(DP_mult_214_n1580), 
        .A(DP_mult_214_n1615), .ZN(DP_mult_214_n1848) );
  OAI221_X1 DP_mult_214_U1483 ( .B1(DP_mult_214_n1617), .B2(DP_mult_214_n1582), 
        .C1(DP_mult_214_n1620), .C2(DP_mult_214_n1578), .A(DP_mult_214_n1848), 
        .ZN(DP_mult_214_n1847) );
  XNOR2_X1 DP_mult_214_U1482 ( .A(DP_coeff_ret0[11]), .B(DP_mult_214_n1847), 
        .ZN(DP_mult_214_n827) );
  OAI22_X1 DP_mult_214_U1481 ( .A1(DP_mult_214_n1633), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1634), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1846)
         );
  AOI221_X1 DP_mult_214_U1480 ( .B1(DP_mult_214_n1579), .B2(DP_mult_214_n1615), 
        .C1(DP_mult_214_n1580), .C2(DP_mult_214_n1615), .A(DP_mult_214_n1846), 
        .ZN(DP_mult_214_n1845) );
  XNOR2_X1 DP_mult_214_U1479 ( .A(DP_coeff_ret0[11]), .B(DP_mult_214_n1845), 
        .ZN(DP_mult_214_n828) );
  OAI22_X1 DP_mult_214_U1478 ( .A1(DP_mult_214_n1617), .A2(DP_mult_214_n1540), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1844)
         );
  AOI221_X1 DP_mult_214_U1477 ( .B1(DP_mult_214_n1580), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1542), .C2(DP_mult_214_n1375), .A(DP_mult_214_n1844), 
        .ZN(DP_mult_214_n1843) );
  XNOR2_X1 DP_mult_214_U1476 ( .A(DP_coeff_ret0[11]), .B(DP_mult_214_n1843), 
        .ZN(DP_mult_214_n829) );
  OAI22_X1 DP_mult_214_U1475 ( .A1(DP_mult_214_n1640), .A2(DP_mult_214_n1582), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1534), .ZN(DP_mult_214_n1842)
         );
  AOI221_X1 DP_mult_214_U1474 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1542), .C2(DP_mult_214_n1376), .A(DP_mult_214_n1842), 
        .ZN(DP_mult_214_n1841) );
  XNOR2_X1 DP_mult_214_U1473 ( .A(DP_coeff_ret0[11]), .B(DP_mult_214_n1841), 
        .ZN(DP_mult_214_n830) );
  OAI22_X1 DP_mult_214_U1472 ( .A1(DP_mult_214_n1728), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1729), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1840)
         );
  AOI221_X1 DP_mult_214_U1471 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_21_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_20_), .A(DP_mult_214_n1840), .ZN(
        DP_mult_214_n1839) );
  XNOR2_X1 DP_mult_214_U1470 ( .A(DP_coeff_ret0[11]), .B(DP_mult_214_n1839), 
        .ZN(DP_mult_214_n831) );
  OAI22_X1 DP_mult_214_U1469 ( .A1(DP_mult_214_n1724), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1725), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1838)
         );
  AOI221_X1 DP_mult_214_U1468 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_20_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_19_), .A(DP_mult_214_n1838), .ZN(
        DP_mult_214_n1837) );
  XNOR2_X1 DP_mult_214_U1467 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1837), 
        .ZN(DP_mult_214_n832) );
  OAI22_X1 DP_mult_214_U1466 ( .A1(DP_mult_214_n1720), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1721), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1836)
         );
  AOI221_X1 DP_mult_214_U1465 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_19_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_18_), .A(DP_mult_214_n1836), .ZN(
        DP_mult_214_n1835) );
  XNOR2_X1 DP_mult_214_U1464 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1835), 
        .ZN(DP_mult_214_n833) );
  OAI22_X1 DP_mult_214_U1463 ( .A1(DP_mult_214_n1716), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1717), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1834)
         );
  AOI221_X1 DP_mult_214_U1462 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_18_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_17_), .A(DP_mult_214_n1834), .ZN(
        DP_mult_214_n1833) );
  XNOR2_X1 DP_mult_214_U1461 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1833), 
        .ZN(DP_mult_214_n834) );
  OAI22_X1 DP_mult_214_U1460 ( .A1(DP_mult_214_n1712), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1713), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1832)
         );
  AOI221_X1 DP_mult_214_U1459 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_17_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_16_), .A(DP_mult_214_n1832), .ZN(
        DP_mult_214_n1831) );
  XNOR2_X1 DP_mult_214_U1458 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1831), 
        .ZN(DP_mult_214_n835) );
  OAI22_X1 DP_mult_214_U1457 ( .A1(DP_mult_214_n1708), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1709), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1830)
         );
  AOI221_X1 DP_mult_214_U1456 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_16_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_15_), .A(DP_mult_214_n1830), .ZN(
        DP_mult_214_n1829) );
  XNOR2_X1 DP_mult_214_U1455 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1829), 
        .ZN(DP_mult_214_n836) );
  OAI22_X1 DP_mult_214_U1454 ( .A1(DP_mult_214_n1704), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1705), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1828)
         );
  AOI221_X1 DP_mult_214_U1453 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_15_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_14_), .A(DP_mult_214_n1828), .ZN(
        DP_mult_214_n1827) );
  XNOR2_X1 DP_mult_214_U1452 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1827), 
        .ZN(DP_mult_214_n837) );
  OAI22_X1 DP_mult_214_U1451 ( .A1(DP_mult_214_n1700), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1701), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1826)
         );
  AOI221_X1 DP_mult_214_U1450 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_14_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_13_), .A(DP_mult_214_n1826), .ZN(
        DP_mult_214_n1825) );
  XNOR2_X1 DP_mult_214_U1449 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1825), 
        .ZN(DP_mult_214_n838) );
  OAI22_X1 DP_mult_214_U1448 ( .A1(DP_mult_214_n1696), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1697), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1824)
         );
  AOI221_X1 DP_mult_214_U1447 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_13_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_12_), .A(DP_mult_214_n1824), .ZN(
        DP_mult_214_n1823) );
  XNOR2_X1 DP_mult_214_U1446 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1823), 
        .ZN(DP_mult_214_n839) );
  OAI22_X1 DP_mult_214_U1445 ( .A1(DP_mult_214_n1692), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1693), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1822)
         );
  AOI221_X1 DP_mult_214_U1444 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_12_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_11_), .A(DP_mult_214_n1822), .ZN(
        DP_mult_214_n1821) );
  XNOR2_X1 DP_mult_214_U1443 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1821), 
        .ZN(DP_mult_214_n840) );
  OAI22_X1 DP_mult_214_U1442 ( .A1(DP_mult_214_n1688), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1689), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1820)
         );
  AOI221_X1 DP_mult_214_U1441 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_11_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_10_), .A(DP_mult_214_n1820), .ZN(
        DP_mult_214_n1819) );
  XNOR2_X1 DP_mult_214_U1440 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1819), 
        .ZN(DP_mult_214_n841) );
  OAI22_X1 DP_mult_214_U1439 ( .A1(DP_mult_214_n1684), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1685), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1818)
         );
  AOI221_X1 DP_mult_214_U1438 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_10_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_9_), .A(DP_mult_214_n1818), .ZN(
        DP_mult_214_n1817) );
  XNOR2_X1 DP_mult_214_U1437 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1817), 
        .ZN(DP_mult_214_n842) );
  OAI22_X1 DP_mult_214_U1436 ( .A1(DP_mult_214_n1680), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1681), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1816)
         );
  AOI221_X1 DP_mult_214_U1435 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_9_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_8_), .A(DP_mult_214_n1816), .ZN(
        DP_mult_214_n1815) );
  XNOR2_X1 DP_mult_214_U1434 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1815), 
        .ZN(DP_mult_214_n843) );
  OAI22_X1 DP_mult_214_U1433 ( .A1(DP_mult_214_n1676), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1677), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1814)
         );
  AOI221_X1 DP_mult_214_U1432 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_8_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_7_), .A(DP_mult_214_n1814), .ZN(
        DP_mult_214_n1813) );
  XNOR2_X1 DP_mult_214_U1431 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1813), 
        .ZN(DP_mult_214_n844) );
  OAI22_X1 DP_mult_214_U1430 ( .A1(DP_mult_214_n1672), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1673), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1812)
         );
  AOI221_X1 DP_mult_214_U1429 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_7_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_6_), .A(DP_mult_214_n1812), .ZN(
        DP_mult_214_n1811) );
  XNOR2_X1 DP_mult_214_U1428 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1811), 
        .ZN(DP_mult_214_n845) );
  OAI22_X1 DP_mult_214_U1427 ( .A1(DP_mult_214_n1668), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1669), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1810)
         );
  AOI221_X1 DP_mult_214_U1426 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_6_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_5_), .A(DP_mult_214_n1810), .ZN(
        DP_mult_214_n1809) );
  XNOR2_X1 DP_mult_214_U1425 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1809), 
        .ZN(DP_mult_214_n846) );
  OAI22_X1 DP_mult_214_U1424 ( .A1(DP_mult_214_n1664), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1665), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1808)
         );
  AOI221_X1 DP_mult_214_U1423 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_5_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_4_), .A(DP_mult_214_n1808), .ZN(
        DP_mult_214_n1807) );
  XNOR2_X1 DP_mult_214_U1422 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1807), 
        .ZN(DP_mult_214_n847) );
  OAI22_X1 DP_mult_214_U1421 ( .A1(DP_mult_214_n1660), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1661), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1806)
         );
  AOI221_X1 DP_mult_214_U1420 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_4_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_3_), .A(DP_mult_214_n1806), .ZN(
        DP_mult_214_n1805) );
  XNOR2_X1 DP_mult_214_U1419 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1805), 
        .ZN(DP_mult_214_n848) );
  OAI22_X1 DP_mult_214_U1418 ( .A1(DP_mult_214_n1657), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1649), .B2(DP_mult_214_n1582), .ZN(DP_mult_214_n1804)
         );
  AOI221_X1 DP_mult_214_U1417 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_3_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_2_), .A(DP_mult_214_n1804), .ZN(
        DP_mult_214_n1803) );
  XNOR2_X1 DP_mult_214_U1416 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1803), 
        .ZN(DP_mult_214_n849) );
  OAI22_X1 DP_mult_214_U1415 ( .A1(DP_mult_214_n1653), .A2(DP_mult_214_n1578), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1581), .ZN(DP_mult_214_n1801)
         );
  AOI221_X1 DP_mult_214_U1414 ( .B1(DP_mult_214_n1579), .B2(DP_sw0_2_), .C1(
        DP_mult_214_n1580), .C2(DP_sw0_1_), .A(DP_mult_214_n1801), .ZN(
        DP_mult_214_n1800) );
  XNOR2_X1 DP_mult_214_U1413 ( .A(DP_mult_214_n1602), .B(DP_mult_214_n1800), 
        .ZN(DP_mult_214_n850) );
  OAI222_X1 DP_mult_214_U1412 ( .A1(DP_mult_214_n1649), .A2(DP_mult_214_n1540), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1534), .C1(DP_mult_214_n1650), 
        .C2(DP_mult_214_n1578), .ZN(DP_mult_214_n1799) );
  XNOR2_X1 DP_mult_214_U1411 ( .A(DP_mult_214_n1799), .B(DP_mult_214_n1603), 
        .ZN(DP_mult_214_n851) );
  OAI22_X1 DP_mult_214_U1410 ( .A1(DP_mult_214_n1565), .A2(DP_mult_214_n1540), 
        .B1(DP_mult_214_n1565), .B2(DP_mult_214_n1578), .ZN(DP_mult_214_n1798)
         );
  XNOR2_X1 DP_mult_214_U1409 ( .A(DP_mult_214_n1798), .B(DP_mult_214_n1603), 
        .ZN(DP_mult_214_n852) );
  XOR2_X1 DP_mult_214_U1408 ( .A(DP_coeff_ret0[6]), .B(DP_mult_214_n1599), .Z(
        DP_mult_214_n1797) );
  XNOR2_X1 DP_mult_214_U1407 ( .A(DP_coeff_ret0[7]), .B(DP_mult_214_n1601), 
        .ZN(DP_mult_214_n1796) );
  XNOR2_X1 DP_mult_214_U1406 ( .A(DP_coeff_ret0[6]), .B(DP_coeff_ret0[7]), 
        .ZN(DP_mult_214_n1795) );
  NAND3_X1 DP_mult_214_U1405 ( .A1(DP_mult_214_n1797), .A2(DP_mult_214_n1796), 
        .A3(DP_mult_214_n1795), .ZN(DP_mult_214_n1747) );
  INV_X1 DP_mult_214_U1404 ( .A(DP_mult_214_n1797), .ZN(DP_mult_214_n1794) );
  OAI21_X1 DP_mult_214_U1403 ( .B1(DP_mult_214_n1574), .B2(DP_mult_214_n1575), 
        .A(DP_mult_214_n1615), .ZN(DP_mult_214_n1793) );
  OAI221_X1 DP_mult_214_U1402 ( .B1(DP_mult_214_n1617), .B2(DP_mult_214_n1577), 
        .C1(DP_mult_214_n1620), .C2(DP_mult_214_n1573), .A(DP_mult_214_n1793), 
        .ZN(DP_mult_214_n1792) );
  XNOR2_X1 DP_mult_214_U1401 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1792), 
        .ZN(DP_mult_214_n853) );
  OAI22_X1 DP_mult_214_U1400 ( .A1(DP_mult_214_n1633), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1634), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1791)
         );
  AOI221_X1 DP_mult_214_U1399 ( .B1(DP_mult_214_n1574), .B2(DP_mult_214_n1614), 
        .C1(DP_mult_214_n1575), .C2(DP_mult_214_n1615), .A(DP_mult_214_n1791), 
        .ZN(DP_mult_214_n1790) );
  XNOR2_X1 DP_mult_214_U1398 ( .A(DP_coeff_ret0[8]), .B(DP_mult_214_n1790), 
        .ZN(DP_mult_214_n854) );
  OAI22_X1 DP_mult_214_U1397 ( .A1(DP_mult_214_n1617), .A2(DP_mult_214_n1535), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1789)
         );
  AOI221_X1 DP_mult_214_U1396 ( .B1(DP_mult_214_n1575), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1533), .C2(DP_mult_214_n1375), .A(DP_mult_214_n1789), 
        .ZN(DP_mult_214_n1788) );
  XNOR2_X1 DP_mult_214_U1395 ( .A(DP_coeff_ret0[8]), .B(DP_mult_214_n1788), 
        .ZN(DP_mult_214_n855) );
  OAI22_X1 DP_mult_214_U1394 ( .A1(DP_mult_214_n1640), .A2(DP_mult_214_n1577), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1537), .ZN(DP_mult_214_n1787)
         );
  AOI221_X1 DP_mult_214_U1393 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1533), .C2(DP_mult_214_n1376), .A(DP_mult_214_n1787), 
        .ZN(DP_mult_214_n1786) );
  XNOR2_X1 DP_mult_214_U1392 ( .A(DP_coeff_ret0[8]), .B(DP_mult_214_n1786), 
        .ZN(DP_mult_214_n856) );
  OAI22_X1 DP_mult_214_U1391 ( .A1(DP_mult_214_n1728), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1729), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1785)
         );
  AOI221_X1 DP_mult_214_U1390 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_21_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_20_), .A(DP_mult_214_n1785), .ZN(
        DP_mult_214_n1784) );
  XNOR2_X1 DP_mult_214_U1389 ( .A(DP_coeff_ret0[8]), .B(DP_mult_214_n1784), 
        .ZN(DP_mult_214_n857) );
  OAI22_X1 DP_mult_214_U1388 ( .A1(DP_mult_214_n1724), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1725), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1783)
         );
  AOI221_X1 DP_mult_214_U1387 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_20_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_19_), .A(DP_mult_214_n1783), .ZN(
        DP_mult_214_n1782) );
  XNOR2_X1 DP_mult_214_U1386 ( .A(DP_coeff_ret0[8]), .B(DP_mult_214_n1782), 
        .ZN(DP_mult_214_n858) );
  OAI22_X1 DP_mult_214_U1385 ( .A1(DP_mult_214_n1720), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1721), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1781)
         );
  AOI221_X1 DP_mult_214_U1384 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_19_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_18_), .A(DP_mult_214_n1781), .ZN(
        DP_mult_214_n1780) );
  XNOR2_X1 DP_mult_214_U1383 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1780), 
        .ZN(DP_mult_214_n859) );
  OAI22_X1 DP_mult_214_U1382 ( .A1(DP_mult_214_n1716), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1717), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1779)
         );
  AOI221_X1 DP_mult_214_U1381 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_18_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_17_), .A(DP_mult_214_n1779), .ZN(
        DP_mult_214_n1778) );
  XNOR2_X1 DP_mult_214_U1380 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1778), 
        .ZN(DP_mult_214_n860) );
  OAI22_X1 DP_mult_214_U1379 ( .A1(DP_mult_214_n1712), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1713), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1777)
         );
  AOI221_X1 DP_mult_214_U1378 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_17_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_16_), .A(DP_mult_214_n1777), .ZN(
        DP_mult_214_n1776) );
  XNOR2_X1 DP_mult_214_U1377 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1776), 
        .ZN(DP_mult_214_n861) );
  OAI22_X1 DP_mult_214_U1376 ( .A1(DP_mult_214_n1708), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1709), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1775)
         );
  AOI221_X1 DP_mult_214_U1375 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_16_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_15_), .A(DP_mult_214_n1775), .ZN(
        DP_mult_214_n1774) );
  XNOR2_X1 DP_mult_214_U1374 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1774), 
        .ZN(DP_mult_214_n862) );
  OAI22_X1 DP_mult_214_U1373 ( .A1(DP_mult_214_n1704), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1705), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1773)
         );
  AOI221_X1 DP_mult_214_U1372 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_15_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_14_), .A(DP_mult_214_n1773), .ZN(
        DP_mult_214_n1772) );
  XNOR2_X1 DP_mult_214_U1371 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1772), 
        .ZN(DP_mult_214_n863) );
  OAI22_X1 DP_mult_214_U1370 ( .A1(DP_mult_214_n1700), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1701), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1771)
         );
  AOI221_X1 DP_mult_214_U1369 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_14_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_13_), .A(DP_mult_214_n1771), .ZN(
        DP_mult_214_n1770) );
  XNOR2_X1 DP_mult_214_U1368 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1770), 
        .ZN(DP_mult_214_n864) );
  OAI22_X1 DP_mult_214_U1367 ( .A1(DP_mult_214_n1696), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1697), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1769)
         );
  AOI221_X1 DP_mult_214_U1366 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_13_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_12_), .A(DP_mult_214_n1769), .ZN(
        DP_mult_214_n1768) );
  XNOR2_X1 DP_mult_214_U1365 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1768), 
        .ZN(DP_mult_214_n865) );
  OAI22_X1 DP_mult_214_U1364 ( .A1(DP_mult_214_n1692), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1693), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1767)
         );
  AOI221_X1 DP_mult_214_U1363 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_12_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_11_), .A(DP_mult_214_n1767), .ZN(
        DP_mult_214_n1766) );
  XNOR2_X1 DP_mult_214_U1362 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1766), 
        .ZN(DP_mult_214_n866) );
  OAI22_X1 DP_mult_214_U1361 ( .A1(DP_mult_214_n1688), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1689), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1765)
         );
  AOI221_X1 DP_mult_214_U1360 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_11_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_10_), .A(DP_mult_214_n1765), .ZN(
        DP_mult_214_n1764) );
  XNOR2_X1 DP_mult_214_U1359 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1764), 
        .ZN(DP_mult_214_n867) );
  OAI22_X1 DP_mult_214_U1358 ( .A1(DP_mult_214_n1684), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1685), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1763)
         );
  AOI221_X1 DP_mult_214_U1357 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_10_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_9_), .A(DP_mult_214_n1763), .ZN(
        DP_mult_214_n1762) );
  XNOR2_X1 DP_mult_214_U1356 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1762), 
        .ZN(DP_mult_214_n868) );
  OAI22_X1 DP_mult_214_U1355 ( .A1(DP_mult_214_n1680), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1681), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1761)
         );
  AOI221_X1 DP_mult_214_U1354 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_9_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_8_), .A(DP_mult_214_n1761), .ZN(
        DP_mult_214_n1760) );
  XNOR2_X1 DP_mult_214_U1353 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1760), 
        .ZN(DP_mult_214_n869) );
  OAI22_X1 DP_mult_214_U1352 ( .A1(DP_mult_214_n1676), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1677), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1759)
         );
  AOI221_X1 DP_mult_214_U1351 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_8_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_7_), .A(DP_mult_214_n1759), .ZN(
        DP_mult_214_n1758) );
  XNOR2_X1 DP_mult_214_U1350 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1758), 
        .ZN(DP_mult_214_n870) );
  OAI22_X1 DP_mult_214_U1349 ( .A1(DP_mult_214_n1672), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1673), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1757)
         );
  AOI221_X1 DP_mult_214_U1348 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_7_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_6_), .A(DP_mult_214_n1757), .ZN(
        DP_mult_214_n1756) );
  XNOR2_X1 DP_mult_214_U1347 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1756), 
        .ZN(DP_mult_214_n871) );
  OAI22_X1 DP_mult_214_U1346 ( .A1(DP_mult_214_n1668), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1669), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1755)
         );
  AOI221_X1 DP_mult_214_U1345 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_6_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_5_), .A(DP_mult_214_n1755), .ZN(
        DP_mult_214_n1754) );
  XNOR2_X1 DP_mult_214_U1344 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1754), 
        .ZN(DP_mult_214_n872) );
  OAI22_X1 DP_mult_214_U1343 ( .A1(DP_mult_214_n1664), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1665), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1753)
         );
  AOI221_X1 DP_mult_214_U1342 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_5_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_4_), .A(DP_mult_214_n1753), .ZN(
        DP_mult_214_n1752) );
  XNOR2_X1 DP_mult_214_U1341 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1752), 
        .ZN(DP_mult_214_n873) );
  OAI22_X1 DP_mult_214_U1340 ( .A1(DP_mult_214_n1660), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1661), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1751)
         );
  AOI221_X1 DP_mult_214_U1339 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_4_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_3_), .A(DP_mult_214_n1751), .ZN(
        DP_mult_214_n1750) );
  XNOR2_X1 DP_mult_214_U1338 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1750), 
        .ZN(DP_mult_214_n874) );
  OAI22_X1 DP_mult_214_U1337 ( .A1(DP_mult_214_n1657), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1649), .B2(DP_mult_214_n1577), .ZN(DP_mult_214_n1749)
         );
  AOI221_X1 DP_mult_214_U1336 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_3_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_2_), .A(DP_mult_214_n1749), .ZN(
        DP_mult_214_n1748) );
  XNOR2_X1 DP_mult_214_U1335 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1748), 
        .ZN(DP_mult_214_n875) );
  OAI22_X1 DP_mult_214_U1334 ( .A1(DP_mult_214_n1653), .A2(DP_mult_214_n1573), 
        .B1(DP_mult_214_n1565), .B2(DP_mult_214_n1576), .ZN(DP_mult_214_n1746)
         );
  AOI221_X1 DP_mult_214_U1333 ( .B1(DP_mult_214_n1574), .B2(DP_sw0_2_), .C1(
        DP_mult_214_n1575), .C2(DP_sw0_1_), .A(DP_mult_214_n1746), .ZN(
        DP_mult_214_n1745) );
  XNOR2_X1 DP_mult_214_U1332 ( .A(DP_mult_214_n1600), .B(DP_mult_214_n1745), 
        .ZN(DP_mult_214_n876) );
  OAI222_X1 DP_mult_214_U1331 ( .A1(DP_mult_214_n1649), .A2(DP_mult_214_n1535), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1537), .C1(DP_mult_214_n1650), 
        .C2(DP_mult_214_n1573), .ZN(DP_mult_214_n1744) );
  XNOR2_X1 DP_mult_214_U1330 ( .A(DP_mult_214_n1744), .B(DP_mult_214_n1601), 
        .ZN(DP_mult_214_n877) );
  OAI22_X1 DP_mult_214_U1329 ( .A1(DP_mult_214_n1565), .A2(DP_mult_214_n1535), 
        .B1(DP_mult_214_n1565), .B2(DP_mult_214_n1573), .ZN(DP_mult_214_n1743)
         );
  XNOR2_X1 DP_mult_214_U1328 ( .A(DP_mult_214_n1743), .B(DP_mult_214_n1601), 
        .ZN(DP_mult_214_n878) );
  XOR2_X1 DP_mult_214_U1327 ( .A(DP_coeff_ret0[3]), .B(DP_mult_214_n1742), .Z(
        DP_mult_214_n1741) );
  XNOR2_X1 DP_mult_214_U1326 ( .A(DP_coeff_ret0[4]), .B(DP_mult_214_n1599), 
        .ZN(DP_mult_214_n1740) );
  XNOR2_X1 DP_mult_214_U1325 ( .A(DP_coeff_ret0[3]), .B(DP_coeff_ret0[4]), 
        .ZN(DP_mult_214_n1739) );
  NAND3_X1 DP_mult_214_U1324 ( .A1(DP_mult_214_n1741), .A2(DP_mult_214_n1740), 
        .A3(DP_mult_214_n1739), .ZN(DP_mult_214_n1654) );
  INV_X1 DP_mult_214_U1323 ( .A(DP_mult_214_n1741), .ZN(DP_mult_214_n1738) );
  OAI21_X1 DP_mult_214_U1322 ( .B1(DP_mult_214_n1569), .B2(DP_mult_214_n1570), 
        .A(DP_mult_214_n1615), .ZN(DP_mult_214_n1737) );
  OAI221_X1 DP_mult_214_U1321 ( .B1(DP_mult_214_n1617), .B2(DP_mult_214_n1572), 
        .C1(DP_mult_214_n1620), .C2(DP_mult_214_n1568), .A(DP_mult_214_n1737), 
        .ZN(DP_mult_214_n1736) );
  XNOR2_X1 DP_mult_214_U1320 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1736), 
        .ZN(DP_mult_214_n879) );
  OAI22_X1 DP_mult_214_U1319 ( .A1(DP_mult_214_n1633), .A2(DP_mult_214_n1568), 
        .B1(DP_mult_214_n1634), .B2(DP_mult_214_n1572), .ZN(DP_mult_214_n1735)
         );
  AOI221_X1 DP_mult_214_U1318 ( .B1(DP_mult_214_n1569), .B2(DP_mult_214_n1614), 
        .C1(DP_mult_214_n1570), .C2(DP_mult_214_n1615), .A(DP_mult_214_n1735), 
        .ZN(DP_mult_214_n1734) );
  XNOR2_X1 DP_mult_214_U1317 ( .A(DP_coeff_ret0[5]), .B(DP_mult_214_n1734), 
        .ZN(DP_mult_214_n880) );
  OAI22_X1 DP_mult_214_U1316 ( .A1(DP_mult_214_n1616), .A2(DP_mult_214_n1539), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1572), .ZN(DP_mult_214_n1733)
         );
  AOI221_X1 DP_mult_214_U1315 ( .B1(DP_mult_214_n1570), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1536), .C2(DP_mult_214_n1375), .A(DP_mult_214_n1733), 
        .ZN(DP_mult_214_n1732) );
  XNOR2_X1 DP_mult_214_U1314 ( .A(DP_coeff_ret0[5]), .B(DP_mult_214_n1732), 
        .ZN(DP_mult_214_n881) );
  OAI22_X1 DP_mult_214_U1313 ( .A1(DP_mult_214_n1640), .A2(DP_mult_214_n1572), 
        .B1(DP_mult_214_n1643), .B2(DP_mult_214_n1538), .ZN(DP_mult_214_n1731)
         );
  AOI221_X1 DP_mult_214_U1312 ( .B1(DP_mult_214_n1569), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1536), .C2(DP_mult_214_n1376), .A(DP_mult_214_n1731), 
        .ZN(DP_mult_214_n1730) );
  XNOR2_X1 DP_mult_214_U1311 ( .A(DP_coeff_ret0[5]), .B(DP_mult_214_n1730), 
        .ZN(DP_mult_214_n882) );
  OAI22_X1 DP_mult_214_U1310 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1728), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1729), .ZN(DP_mult_214_n1727)
         );
  AOI221_X1 DP_mult_214_U1309 ( .B1(DP_mult_214_n1569), .B2(DP_sw0_21_), .C1(
        DP_mult_214_n1570), .C2(DP_sw0_20_), .A(DP_mult_214_n1727), .ZN(
        DP_mult_214_n1726) );
  XNOR2_X1 DP_mult_214_U1308 ( .A(DP_coeff_ret0[5]), .B(DP_mult_214_n1726), 
        .ZN(DP_mult_214_n883) );
  OAI22_X1 DP_mult_214_U1307 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1724), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1725), .ZN(DP_mult_214_n1723)
         );
  AOI221_X1 DP_mult_214_U1306 ( .B1(DP_mult_214_n1569), .B2(DP_sw0_20_), .C1(
        DP_sw0_19_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1723), .ZN(
        DP_mult_214_n1722) );
  XNOR2_X1 DP_mult_214_U1305 ( .A(DP_coeff_ret0[5]), .B(DP_mult_214_n1722), 
        .ZN(DP_mult_214_n884) );
  OAI22_X1 DP_mult_214_U1304 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1720), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1721), .ZN(DP_mult_214_n1719)
         );
  AOI221_X1 DP_mult_214_U1303 ( .B1(DP_sw0_19_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_18_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1719), .ZN(
        DP_mult_214_n1718) );
  XNOR2_X1 DP_mult_214_U1302 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1718), 
        .ZN(DP_mult_214_n885) );
  OAI22_X1 DP_mult_214_U1301 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1716), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1717), .ZN(DP_mult_214_n1715)
         );
  AOI221_X1 DP_mult_214_U1300 ( .B1(DP_sw0_18_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_17_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1715), .ZN(
        DP_mult_214_n1714) );
  XNOR2_X1 DP_mult_214_U1299 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1714), 
        .ZN(DP_mult_214_n886) );
  OAI22_X1 DP_mult_214_U1298 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1712), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1713), .ZN(DP_mult_214_n1711)
         );
  AOI221_X1 DP_mult_214_U1297 ( .B1(DP_sw0_17_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_16_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1711), .ZN(
        DP_mult_214_n1710) );
  XNOR2_X1 DP_mult_214_U1296 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1710), 
        .ZN(DP_mult_214_n887) );
  OAI22_X1 DP_mult_214_U1295 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1708), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1709), .ZN(DP_mult_214_n1707)
         );
  AOI221_X1 DP_mult_214_U1294 ( .B1(DP_sw0_16_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_15_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1707), .ZN(
        DP_mult_214_n1706) );
  XNOR2_X1 DP_mult_214_U1293 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1706), 
        .ZN(DP_mult_214_n888) );
  OAI22_X1 DP_mult_214_U1292 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1704), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1705), .ZN(DP_mult_214_n1703)
         );
  AOI221_X1 DP_mult_214_U1291 ( .B1(DP_sw0_15_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_14_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1703), .ZN(
        DP_mult_214_n1702) );
  XNOR2_X1 DP_mult_214_U1290 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1702), 
        .ZN(DP_mult_214_n889) );
  OAI22_X1 DP_mult_214_U1289 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1700), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1701), .ZN(DP_mult_214_n1699)
         );
  AOI221_X1 DP_mult_214_U1288 ( .B1(DP_sw0_14_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_13_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1699), .ZN(
        DP_mult_214_n1698) );
  XNOR2_X1 DP_mult_214_U1287 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1698), 
        .ZN(DP_mult_214_n890) );
  OAI22_X1 DP_mult_214_U1286 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1696), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1697), .ZN(DP_mult_214_n1695)
         );
  AOI221_X1 DP_mult_214_U1285 ( .B1(DP_sw0_13_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_12_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1695), .ZN(
        DP_mult_214_n1694) );
  XNOR2_X1 DP_mult_214_U1284 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1694), 
        .ZN(DP_mult_214_n891) );
  OAI22_X1 DP_mult_214_U1283 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1692), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1693), .ZN(DP_mult_214_n1691)
         );
  AOI221_X1 DP_mult_214_U1282 ( .B1(DP_sw0_12_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_11_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1691), .ZN(
        DP_mult_214_n1690) );
  XNOR2_X1 DP_mult_214_U1281 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1690), 
        .ZN(DP_mult_214_n892) );
  OAI22_X1 DP_mult_214_U1280 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1688), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1689), .ZN(DP_mult_214_n1687)
         );
  AOI221_X1 DP_mult_214_U1279 ( .B1(DP_sw0_11_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_10_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1687), .ZN(
        DP_mult_214_n1686) );
  XNOR2_X1 DP_mult_214_U1278 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1686), 
        .ZN(DP_mult_214_n893) );
  OAI22_X1 DP_mult_214_U1277 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1684), 
        .B1(DP_mult_214_n1572), .B2(DP_mult_214_n1685), .ZN(DP_mult_214_n1683)
         );
  AOI221_X1 DP_mult_214_U1276 ( .B1(DP_sw0_10_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_9_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1683), .ZN(
        DP_mult_214_n1682) );
  XNOR2_X1 DP_mult_214_U1275 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1682), 
        .ZN(DP_mult_214_n894) );
  OAI22_X1 DP_mult_214_U1274 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1680), 
        .B1(DP_mult_214_n1572), .B2(DP_mult_214_n1681), .ZN(DP_mult_214_n1679)
         );
  AOI221_X1 DP_mult_214_U1273 ( .B1(DP_sw0_9_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_8_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1679), .ZN(
        DP_mult_214_n1678) );
  XNOR2_X1 DP_mult_214_U1272 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1678), 
        .ZN(DP_mult_214_n895) );
  OAI22_X1 DP_mult_214_U1271 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1676), 
        .B1(DP_mult_214_n1571), .B2(DP_mult_214_n1677), .ZN(DP_mult_214_n1675)
         );
  AOI221_X1 DP_mult_214_U1270 ( .B1(DP_sw0_8_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_7_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1675), .ZN(
        DP_mult_214_n1674) );
  XNOR2_X1 DP_mult_214_U1269 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1674), 
        .ZN(DP_mult_214_n896) );
  OAI22_X1 DP_mult_214_U1268 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1672), 
        .B1(DP_mult_214_n1572), .B2(DP_mult_214_n1673), .ZN(DP_mult_214_n1671)
         );
  AOI221_X1 DP_mult_214_U1267 ( .B1(DP_sw0_7_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_6_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1671), .ZN(
        DP_mult_214_n1670) );
  XNOR2_X1 DP_mult_214_U1266 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1670), 
        .ZN(DP_mult_214_n897) );
  OAI22_X1 DP_mult_214_U1265 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1668), 
        .B1(DP_mult_214_n1572), .B2(DP_mult_214_n1669), .ZN(DP_mult_214_n1667)
         );
  AOI221_X1 DP_mult_214_U1264 ( .B1(DP_sw0_6_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_5_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1667), .ZN(
        DP_mult_214_n1666) );
  XNOR2_X1 DP_mult_214_U1263 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1666), 
        .ZN(DP_mult_214_n898) );
  OAI22_X1 DP_mult_214_U1262 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1664), 
        .B1(DP_mult_214_n1572), .B2(DP_mult_214_n1665), .ZN(DP_mult_214_n1663)
         );
  AOI221_X1 DP_mult_214_U1261 ( .B1(DP_sw0_5_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_4_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1663), .ZN(
        DP_mult_214_n1662) );
  XNOR2_X1 DP_mult_214_U1260 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1662), 
        .ZN(DP_mult_214_n899) );
  OAI22_X1 DP_mult_214_U1259 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1660), 
        .B1(DP_mult_214_n1661), .B2(DP_mult_214_n1572), .ZN(DP_mult_214_n1659)
         );
  AOI221_X1 DP_mult_214_U1258 ( .B1(DP_sw0_4_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_3_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1659), .ZN(
        DP_mult_214_n1658) );
  XNOR2_X1 DP_mult_214_U1257 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1658), 
        .ZN(DP_mult_214_n900) );
  OAI22_X1 DP_mult_214_U1256 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1657), 
        .B1(DP_mult_214_n1649), .B2(DP_mult_214_n1572), .ZN(DP_mult_214_n1656)
         );
  AOI221_X1 DP_mult_214_U1255 ( .B1(DP_sw0_3_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_2_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1656), .ZN(
        DP_mult_214_n1655) );
  XNOR2_X1 DP_mult_214_U1254 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1655), 
        .ZN(DP_mult_214_n901) );
  OAI22_X1 DP_mult_214_U1253 ( .A1(DP_mult_214_n1568), .A2(DP_mult_214_n1653), 
        .B1(DP_mult_214_n1565), .B2(DP_mult_214_n1572), .ZN(DP_mult_214_n1652)
         );
  AOI221_X1 DP_mult_214_U1252 ( .B1(DP_sw0_2_), .B2(DP_mult_214_n1569), .C1(
        DP_sw0_1_), .C2(DP_mult_214_n1570), .A(DP_mult_214_n1652), .ZN(
        DP_mult_214_n1651) );
  XNOR2_X1 DP_mult_214_U1251 ( .A(DP_mult_214_n1598), .B(DP_mult_214_n1651), 
        .ZN(DP_mult_214_n902) );
  OAI222_X1 DP_mult_214_U1250 ( .A1(DP_mult_214_n1539), .A2(DP_mult_214_n1649), 
        .B1(DP_mult_214_n1566), .B2(DP_mult_214_n1538), .C1(DP_mult_214_n1568), 
        .C2(DP_mult_214_n1650), .ZN(DP_mult_214_n1648) );
  XNOR2_X1 DP_mult_214_U1249 ( .A(DP_mult_214_n1648), .B(DP_mult_214_n1599), 
        .ZN(DP_mult_214_n903) );
  OAI22_X1 DP_mult_214_U1248 ( .A1(DP_mult_214_n1565), .A2(DP_mult_214_n1539), 
        .B1(DP_mult_214_n1568), .B2(DP_mult_214_n1567), .ZN(DP_mult_214_n1646)
         );
  XNOR2_X1 DP_mult_214_U1247 ( .A(DP_mult_214_n1646), .B(DP_mult_214_n1599), 
        .ZN(DP_mult_214_n904) );
  OAI22_X1 DP_mult_214_U1246 ( .A1(DP_mult_214_n1633), .A2(DP_mult_214_n1564), 
        .B1(DP_mult_214_n1634), .B2(DP_mult_214_n1639), .ZN(DP_mult_214_n1645)
         );
  AOI221_X1 DP_mult_214_U1245 ( .B1(DP_mult_214_n1561), .B2(DP_mult_214_n1614), 
        .C1(DP_mult_214_n1563), .C2(DP_mult_214_n1615), .A(DP_mult_214_n1645), 
        .ZN(DP_mult_214_n1644) );
  XNOR2_X1 DP_mult_214_U1244 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n1644), 
        .ZN(DP_mult_214_n906) );
  OAI22_X1 DP_mult_214_U1243 ( .A1(DP_mult_214_n1643), .A2(DP_mult_214_n1639), 
        .B1(DP_mult_214_n1617), .B2(DP_mult_214_n1541), .ZN(DP_mult_214_n1642)
         );
  AOI221_X1 DP_mult_214_U1242 ( .B1(DP_mult_214_n1563), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1550), .C2(DP_mult_214_n1375), .A(DP_mult_214_n1642), 
        .ZN(DP_mult_214_n1641) );
  XNOR2_X1 DP_mult_214_U1241 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n1641), 
        .ZN(DP_mult_214_n907) );
  INV_X1 DP_mult_214_U1240 ( .A(DP_mult_214_n1376), .ZN(DP_mult_214_n1638) );
  OAI22_X1 DP_mult_214_U1239 ( .A1(DP_mult_214_n1564), .A2(DP_mult_214_n1638), 
        .B1(DP_mult_214_n1639), .B2(DP_mult_214_n1640), .ZN(DP_mult_214_n1637)
         );
  AOI221_X1 DP_mult_214_U1238 ( .B1(DP_mult_214_n1561), .B2(DP_sw0_22_), .C1(
        DP_mult_214_n1563), .C2(DP_sw0_21_), .A(DP_mult_214_n1637), .ZN(
        DP_mult_214_n1635) );
  XNOR2_X1 DP_mult_214_U1237 ( .A(DP_coeff_ret0[2]), .B(DP_mult_214_n1635), 
        .ZN(DP_mult_214_n908) );
  OAI22_X1 DP_mult_214_U1236 ( .A1(DP_mult_214_n1558), .A2(DP_mult_214_n1633), 
        .B1(DP_mult_214_n1557), .B2(DP_mult_214_n1634), .ZN(DP_mult_214_n1632)
         );
  AOI221_X1 DP_mult_214_U1235 ( .B1(DP_mult_214_n1613), .B2(DP_mult_214_n1559), 
        .C1(DP_mult_214_n1560), .C2(DP_mult_214_n1615), .A(DP_mult_214_n1632), 
        .ZN(DP_mult_214_n1631) );
  XOR2_X1 DP_mult_214_U1234 ( .A(DP_coeff_ret0[23]), .B(DP_mult_214_n1631), 
        .Z(DP_mult_214_n1625) );
  INV_X1 DP_mult_214_U1233 ( .A(DP_mult_214_n1625), .ZN(DP_mult_214_n1621) );
  OAI21_X1 DP_mult_214_U1232 ( .B1(DP_mult_214_n1559), .B2(DP_mult_214_n1560), 
        .A(DP_mult_214_n1615), .ZN(DP_mult_214_n1630) );
  OAI221_X1 DP_mult_214_U1231 ( .B1(DP_mult_214_n1617), .B2(DP_mult_214_n1557), 
        .C1(DP_mult_214_n1620), .C2(DP_mult_214_n1558), .A(DP_mult_214_n1630), 
        .ZN(DP_mult_214_n1628) );
  XOR2_X1 DP_mult_214_U1230 ( .A(DP_mult_214_n1628), .B(DP_mult_214_n1611), 
        .Z(DP_mult_214_n1622) );
  AOI222_X1 DP_mult_214_U1229 ( .A1(DP_mult_214_n1627), .A2(DP_mult_214_n303), 
        .B1(DP_mult_214_n1625), .B2(DP_mult_214_n303), .C1(DP_mult_214_n1627), 
        .C2(DP_mult_214_n1625), .ZN(DP_mult_214_n1624) );
  INV_X1 DP_mult_214_U1228 ( .A(DP_mult_214_n1622), .ZN(DP_mult_214_n1626) );
  OAI22_X1 DP_mult_214_U1227 ( .A1(DP_mult_214_n1624), .A2(DP_mult_214_n1625), 
        .B1(DP_mult_214_n1624), .B2(DP_mult_214_n1626), .ZN(DP_mult_214_n1623)
         );
  AOI21_X1 DP_mult_214_U1226 ( .B1(DP_mult_214_n1621), .B2(DP_mult_214_n1622), 
        .A(DP_mult_214_n1623), .ZN(DP_sw0_coeff_ret0[23]) );
  INV_X1 DP_mult_214_U1225 ( .A(DP_mult_214_n1614), .ZN(DP_mult_214_n1620) );
  INV_X1 DP_mult_214_U1224 ( .A(DP_mult_214_n1614), .ZN(DP_mult_214_n1619) );
  INV_X1 DP_mult_214_U1223 ( .A(DP_mult_214_n1613), .ZN(DP_mult_214_n1618) );
  INV_X1 DP_mult_214_U1222 ( .A(DP_mult_214_n1613), .ZN(DP_mult_214_n1617) );
  INV_X1 DP_mult_214_U1221 ( .A(DP_mult_214_n1612), .ZN(DP_mult_214_n1616) );
  CLKBUF_X1 DP_mult_214_U1220 ( .A(DP_sw0_23_), .Z(DP_mult_214_n1614) );
  CLKBUF_X1 DP_mult_214_U1219 ( .A(DP_sw0_23_), .Z(DP_mult_214_n1613) );
  CLKBUF_X1 DP_mult_214_U1218 ( .A(DP_sw0_23_), .Z(DP_mult_214_n1612) );
  INV_X1 DP_mult_214_U1217 ( .A(DP_coeff_ret0[23]), .ZN(DP_mult_214_n1611) );
  BUF_X1 DP_mult_214_U1216 ( .A(DP_mult_214_n1647), .Z(DP_mult_214_n1567) );
  BUF_X1 DP_mult_214_U1215 ( .A(DP_mult_214_n1647), .Z(DP_mult_214_n1566) );
  BUF_X1 DP_mult_214_U1214 ( .A(DP_mult_214_n1647), .Z(DP_mult_214_n1565) );
  BUF_X1 DP_mult_214_U1213 ( .A(DP_coeff_ret0[20]), .Z(DP_mult_214_n1609) );
  INV_X1 DP_mult_214_U1212 ( .A(DP_coeff_ret0[14]), .ZN(DP_mult_214_n1605) );
  INV_X1 DP_mult_214_U1211 ( .A(DP_coeff_ret0[11]), .ZN(DP_mult_214_n1603) );
  INV_X1 DP_mult_214_U1210 ( .A(DP_coeff_ret0[17]), .ZN(DP_mult_214_n1607) );
  BUF_X1 DP_mult_214_U1209 ( .A(DP_coeff_ret0[20]), .Z(DP_mult_214_n1608) );
  INV_X1 DP_mult_214_U1208 ( .A(DP_mult_214_n1611), .ZN(DP_mult_214_n1610) );
  INV_X1 DP_mult_214_U1207 ( .A(DP_mult_214_n1616), .ZN(DP_mult_214_n1615) );
  OR2_X1 DP_mult_214_U1206 ( .A1(DP_mult_214_n2014), .A2(DP_mult_214_n2015), 
        .ZN(DP_mult_214_n1555) );
  OR2_X1 DP_mult_214_U1205 ( .A1(DP_mult_214_n1959), .A2(DP_mult_214_n1960), 
        .ZN(DP_mult_214_n1554) );
  OR2_X1 DP_mult_214_U1204 ( .A1(DP_mult_214_n1904), .A2(DP_mult_214_n1905), 
        .ZN(DP_mult_214_n1553) );
  OR2_X1 DP_mult_214_U1203 ( .A1(DP_mult_214_n2070), .A2(DP_mult_214_n2069), 
        .ZN(DP_mult_214_n1552) );
  AND2_X1 DP_mult_214_U1202 ( .A1(DP_mult_214_n1904), .A2(DP_mult_214_n1906), 
        .ZN(DP_mult_214_n1551) );
  AND2_X1 DP_mult_214_U1201 ( .A1(DP_coeff_ret0[1]), .A2(DP_mult_214_n2157), 
        .ZN(DP_mult_214_n1550) );
  OR2_X1 DP_mult_214_U1200 ( .A1(DP_mult_214_n1961), .A2(DP_mult_214_n1962), 
        .ZN(DP_mult_214_n1549) );
  OR2_X1 DP_mult_214_U1199 ( .A1(DP_mult_214_n1906), .A2(DP_mult_214_n1907), 
        .ZN(DP_mult_214_n1548) );
  INV_X1 DP_mult_214_U1198 ( .A(DP_mult_214_n1607), .ZN(DP_mult_214_n1606) );
  INV_X1 DP_mult_214_U1197 ( .A(DP_mult_214_n1605), .ZN(DP_mult_214_n1604) );
  INV_X1 DP_mult_214_U1196 ( .A(DP_mult_214_n1603), .ZN(DP_mult_214_n1602) );
  AND2_X1 DP_mult_214_U1195 ( .A1(DP_mult_214_n2070), .A2(DP_mult_214_n2068), 
        .ZN(DP_mult_214_n1547) );
  AND2_X1 DP_mult_214_U1194 ( .A1(DP_mult_214_n1959), .A2(DP_mult_214_n1961), 
        .ZN(DP_mult_214_n1546) );
  AND2_X1 DP_mult_214_U1193 ( .A1(DP_mult_214_n2014), .A2(DP_mult_214_n2016), 
        .ZN(DP_mult_214_n1545) );
  OR2_X1 DP_mult_214_U1192 ( .A1(DP_mult_214_n2068), .A2(DP_mult_214_n2067), 
        .ZN(DP_mult_214_n1544) );
  OR2_X1 DP_mult_214_U1191 ( .A1(DP_mult_214_n2016), .A2(DP_mult_214_n2017), 
        .ZN(DP_mult_214_n1543) );
  BUF_X1 DP_mult_214_U1190 ( .A(DP_mult_214_n1636), .Z(DP_mult_214_n1563) );
  BUF_X1 DP_mult_214_U1189 ( .A(DP_mult_214_n1636), .Z(DP_mult_214_n1562) );
  INV_X1 DP_mult_214_U1188 ( .A(DP_mult_214_n1543), .ZN(DP_mult_214_n1594) );
  INV_X1 DP_mult_214_U1187 ( .A(DP_mult_214_n1549), .ZN(DP_mult_214_n1589) );
  INV_X1 DP_mult_214_U1186 ( .A(DP_mult_214_n1548), .ZN(DP_mult_214_n1584) );
  INV_X1 DP_mult_214_U1185 ( .A(DP_coeff_ret0[5]), .ZN(DP_mult_214_n1599) );
  AND2_X1 DP_mult_214_U1184 ( .A1(DP_mult_214_n1849), .A2(DP_mult_214_n1851), 
        .ZN(DP_mult_214_n1542) );
  OR2_X1 DP_mult_214_U1183 ( .A1(DP_mult_214_n2158), .A2(DP_mult_214_n2157), 
        .ZN(DP_mult_214_n1541) );
  OR2_X1 DP_mult_214_U1182 ( .A1(DP_mult_214_n1851), .A2(DP_mult_214_n1852), 
        .ZN(DP_mult_214_n1540) );
  BUF_X1 DP_mult_214_U1181 ( .A(DP_mult_214_n1912), .Z(DP_mult_214_n1592) );
  BUF_X1 DP_mult_214_U1180 ( .A(DP_mult_214_n1857), .Z(DP_mult_214_n1587) );
  BUF_X1 DP_mult_214_U1179 ( .A(DP_mult_214_n1912), .Z(DP_mult_214_n1591) );
  BUF_X1 DP_mult_214_U1178 ( .A(DP_mult_214_n1857), .Z(DP_mult_214_n1586) );
  BUF_X1 DP_mult_214_U1177 ( .A(DP_mult_214_n1629), .Z(DP_mult_214_n1556) );
  INV_X1 DP_mult_214_U1176 ( .A(DP_mult_214_n1550), .ZN(DP_mult_214_n1564) );
  INV_X1 DP_mult_214_U1175 ( .A(DP_mult_214_n1551), .ZN(DP_mult_214_n1583) );
  INV_X1 DP_mult_214_U1174 ( .A(DP_mult_214_n1555), .ZN(DP_mult_214_n1595) );
  INV_X1 DP_mult_214_U1173 ( .A(DP_mult_214_n1554), .ZN(DP_mult_214_n1590) );
  INV_X1 DP_mult_214_U1172 ( .A(DP_mult_214_n1553), .ZN(DP_mult_214_n1585) );
  INV_X1 DP_mult_214_U1171 ( .A(DP_mult_214_n1552), .ZN(DP_mult_214_n1560) );
  NAND3_X1 DP_mult_214_U1170 ( .A1(DP_mult_214_n2157), .A2(DP_mult_214_n2158), 
        .A3(DP_mult_214_n2158), .ZN(DP_mult_214_n1639) );
  BUF_X1 DP_mult_214_U1169 ( .A(DP_mult_214_n1967), .Z(DP_mult_214_n1597) );
  BUF_X1 DP_mult_214_U1168 ( .A(DP_mult_214_n1967), .Z(DP_mult_214_n1596) );
  BUF_X1 DP_mult_214_U1167 ( .A(DP_mult_214_n1629), .Z(DP_mult_214_n1557) );
  INV_X1 DP_mult_214_U1166 ( .A(DP_mult_214_n1545), .ZN(DP_mult_214_n1593) );
  INV_X1 DP_mult_214_U1165 ( .A(DP_mult_214_n1546), .ZN(DP_mult_214_n1588) );
  INV_X1 DP_mult_214_U1164 ( .A(DP_mult_214_n1544), .ZN(DP_mult_214_n1559) );
  INV_X1 DP_mult_214_U1163 ( .A(DP_mult_214_n1547), .ZN(DP_mult_214_n1558) );
  INV_X1 DP_mult_214_U1162 ( .A(DP_mult_214_n1540), .ZN(DP_mult_214_n1579) );
  INV_X1 DP_mult_214_U1161 ( .A(DP_coeff_ret0[8]), .ZN(DP_mult_214_n1601) );
  OR2_X1 DP_mult_214_U1160 ( .A1(DP_mult_214_n1740), .A2(DP_mult_214_n1741), 
        .ZN(DP_mult_214_n1539) );
  BUF_X1 DP_mult_214_U1159 ( .A(DP_mult_214_n1802), .Z(DP_mult_214_n1582) );
  BUF_X1 DP_mult_214_U1158 ( .A(DP_mult_214_n1802), .Z(DP_mult_214_n1581) );
  OR2_X1 DP_mult_214_U1157 ( .A1(DP_mult_214_n1738), .A2(DP_mult_214_n1739), 
        .ZN(DP_mult_214_n1538) );
  INV_X1 DP_mult_214_U1156 ( .A(DP_mult_214_n1542), .ZN(DP_mult_214_n1578) );
  INV_X1 DP_mult_214_U1155 ( .A(DP_mult_214_n1541), .ZN(DP_mult_214_n1561) );
  INV_X1 DP_mult_214_U1154 ( .A(DP_mult_214_n1599), .ZN(DP_mult_214_n1598) );
  BUF_X1 DP_mult_214_U1153 ( .A(DP_mult_214_n1654), .Z(DP_mult_214_n1571) );
  OR2_X1 DP_mult_214_U1152 ( .A1(DP_mult_214_n1794), .A2(DP_mult_214_n1795), 
        .ZN(DP_mult_214_n1537) );
  AND2_X1 DP_mult_214_U1151 ( .A1(DP_mult_214_n1738), .A2(DP_mult_214_n1740), 
        .ZN(DP_mult_214_n1536) );
  OR2_X1 DP_mult_214_U1150 ( .A1(DP_mult_214_n1796), .A2(DP_mult_214_n1797), 
        .ZN(DP_mult_214_n1535) );
  BUF_X1 DP_mult_214_U1149 ( .A(DP_mult_214_n1654), .Z(DP_mult_214_n1572) );
  INV_X1 DP_mult_214_U1148 ( .A(DP_mult_214_n1539), .ZN(DP_mult_214_n1569) );
  INV_X1 DP_mult_214_U1147 ( .A(DP_mult_214_n1538), .ZN(DP_mult_214_n1570) );
  INV_X1 DP_mult_214_U1146 ( .A(DP_mult_214_n1601), .ZN(DP_mult_214_n1600) );
  INV_X1 DP_mult_214_U1145 ( .A(DP_mult_214_n1535), .ZN(DP_mult_214_n1574) );
  OR2_X1 DP_mult_214_U1144 ( .A1(DP_mult_214_n1849), .A2(DP_mult_214_n1850), 
        .ZN(DP_mult_214_n1534) );
  AND2_X1 DP_mult_214_U1143 ( .A1(DP_mult_214_n1794), .A2(DP_mult_214_n1796), 
        .ZN(DP_mult_214_n1533) );
  BUF_X1 DP_mult_214_U1142 ( .A(DP_mult_214_n1747), .Z(DP_mult_214_n1577) );
  BUF_X1 DP_mult_214_U1141 ( .A(DP_mult_214_n1747), .Z(DP_mult_214_n1576) );
  INV_X1 DP_mult_214_U1140 ( .A(DP_mult_214_n1537), .ZN(DP_mult_214_n1575) );
  INV_X1 DP_mult_214_U1139 ( .A(DP_mult_214_n1536), .ZN(DP_mult_214_n1568) );
  INV_X1 DP_mult_214_U1138 ( .A(DP_mult_214_n1533), .ZN(DP_mult_214_n1573) );
  INV_X1 DP_mult_214_U1137 ( .A(DP_mult_214_n1534), .ZN(DP_mult_214_n1580) );
  HA_X1 DP_mult_214_U1134 ( .A(DP_sw0_0_), .B(DP_sw0_1_), .CO(DP_mult_214_n727), .S(DP_mult_214_n1397) );
  FA_X1 DP_mult_214_U1133 ( .A(DP_sw0_1_), .B(DP_sw0_2_), .CI(DP_mult_214_n727), .CO(DP_mult_214_n726), .S(DP_mult_214_n1396) );
  FA_X1 DP_mult_214_U1132 ( .A(DP_sw0_2_), .B(DP_sw0_3_), .CI(DP_mult_214_n726), .CO(DP_mult_214_n725), .S(DP_mult_214_n1395) );
  FA_X1 DP_mult_214_U1131 ( .A(DP_sw0_3_), .B(DP_sw0_4_), .CI(DP_mult_214_n725), .CO(DP_mult_214_n724), .S(DP_mult_214_n1394) );
  FA_X1 DP_mult_214_U1130 ( .A(DP_sw0_4_), .B(DP_sw0_5_), .CI(DP_mult_214_n724), .CO(DP_mult_214_n723), .S(DP_mult_214_n1393) );
  FA_X1 DP_mult_214_U1129 ( .A(DP_sw0_5_), .B(DP_sw0_6_), .CI(DP_mult_214_n723), .CO(DP_mult_214_n722), .S(DP_mult_214_n1392) );
  FA_X1 DP_mult_214_U1128 ( .A(DP_sw0_6_), .B(DP_sw0_7_), .CI(DP_mult_214_n722), .CO(DP_mult_214_n721), .S(DP_mult_214_n1391) );
  FA_X1 DP_mult_214_U1127 ( .A(DP_sw0_7_), .B(DP_sw0_8_), .CI(DP_mult_214_n721), .CO(DP_mult_214_n720), .S(DP_mult_214_n1390) );
  FA_X1 DP_mult_214_U1126 ( .A(DP_sw0_8_), .B(DP_sw0_9_), .CI(DP_mult_214_n720), .CO(DP_mult_214_n719), .S(DP_mult_214_n1389) );
  FA_X1 DP_mult_214_U1125 ( .A(DP_sw0_9_), .B(DP_sw0_10_), .CI(
        DP_mult_214_n719), .CO(DP_mult_214_n718), .S(DP_mult_214_n1388) );
  FA_X1 DP_mult_214_U1124 ( .A(DP_sw0_10_), .B(DP_sw0_11_), .CI(
        DP_mult_214_n718), .CO(DP_mult_214_n717), .S(DP_mult_214_n1387) );
  FA_X1 DP_mult_214_U1123 ( .A(DP_sw0_11_), .B(DP_sw0_12_), .CI(
        DP_mult_214_n717), .CO(DP_mult_214_n716), .S(DP_mult_214_n1386) );
  FA_X1 DP_mult_214_U1122 ( .A(DP_sw0_12_), .B(DP_sw0_13_), .CI(
        DP_mult_214_n716), .CO(DP_mult_214_n715), .S(DP_mult_214_n1385) );
  FA_X1 DP_mult_214_U1121 ( .A(DP_sw0_13_), .B(DP_sw0_14_), .CI(
        DP_mult_214_n715), .CO(DP_mult_214_n714), .S(DP_mult_214_n1384) );
  FA_X1 DP_mult_214_U1120 ( .A(DP_sw0_14_), .B(DP_sw0_15_), .CI(
        DP_mult_214_n714), .CO(DP_mult_214_n713), .S(DP_mult_214_n1383) );
  FA_X1 DP_mult_214_U1119 ( .A(DP_sw0_15_), .B(DP_sw0_16_), .CI(
        DP_mult_214_n713), .CO(DP_mult_214_n712), .S(DP_mult_214_n1382) );
  FA_X1 DP_mult_214_U1118 ( .A(DP_sw0_16_), .B(DP_sw0_17_), .CI(
        DP_mult_214_n712), .CO(DP_mult_214_n711), .S(DP_mult_214_n1381) );
  FA_X1 DP_mult_214_U1117 ( .A(DP_sw0_17_), .B(DP_sw0_18_), .CI(
        DP_mult_214_n711), .CO(DP_mult_214_n710), .S(DP_mult_214_n1380) );
  FA_X1 DP_mult_214_U1116 ( .A(DP_sw0_18_), .B(DP_sw0_19_), .CI(
        DP_mult_214_n710), .CO(DP_mult_214_n709), .S(DP_mult_214_n1379) );
  FA_X1 DP_mult_214_U1115 ( .A(DP_sw0_19_), .B(DP_sw0_20_), .CI(
        DP_mult_214_n709), .CO(DP_mult_214_n708), .S(DP_mult_214_n1378) );
  FA_X1 DP_mult_214_U1114 ( .A(DP_sw0_20_), .B(DP_sw0_21_), .CI(
        DP_mult_214_n708), .CO(DP_mult_214_n707), .S(DP_mult_214_n1377) );
  FA_X1 DP_mult_214_U1113 ( .A(DP_sw0_21_), .B(DP_sw0_22_), .CI(
        DP_mult_214_n707), .CO(DP_mult_214_n706), .S(DP_mult_214_n1376) );
  FA_X1 DP_mult_214_U1112 ( .A(DP_sw0_22_), .B(DP_mult_214_n1615), .CI(
        DP_mult_214_n706), .CO(DP_mult_214_n1374), .S(DP_mult_214_n1375) );
  HA_X1 DP_mult_214_U408 ( .A(DP_mult_214_n904), .B(DP_mult_214_n1598), .CO(
        DP_mult_214_n687), .S(DP_mult_214_n688) );
  HA_X1 DP_mult_214_U407 ( .A(DP_mult_214_n687), .B(DP_mult_214_n903), .CO(
        DP_mult_214_n685), .S(DP_mult_214_n686) );
  HA_X1 DP_mult_214_U406 ( .A(DP_mult_214_n685), .B(DP_mult_214_n902), .CO(
        DP_mult_214_n683), .S(DP_mult_214_n684) );
  HA_X1 DP_mult_214_U405 ( .A(DP_mult_214_n878), .B(DP_mult_214_n1600), .CO(
        DP_mult_214_n681), .S(DP_mult_214_n682) );
  FA_X1 DP_mult_214_U404 ( .A(DP_mult_214_n901), .B(DP_mult_214_n682), .CI(
        DP_mult_214_n683), .CO(DP_mult_214_n679), .S(DP_mult_214_n680) );
  HA_X1 DP_mult_214_U403 ( .A(DP_mult_214_n681), .B(DP_mult_214_n877), .CO(
        DP_mult_214_n677), .S(DP_mult_214_n678) );
  FA_X1 DP_mult_214_U402 ( .A(DP_mult_214_n900), .B(DP_mult_214_n678), .CI(
        DP_mult_214_n679), .CO(DP_mult_214_n675), .S(DP_mult_214_n676) );
  HA_X1 DP_mult_214_U401 ( .A(DP_mult_214_n677), .B(DP_mult_214_n876), .CO(
        DP_mult_214_n673), .S(DP_mult_214_n674) );
  FA_X1 DP_mult_214_U400 ( .A(DP_mult_214_n899), .B(DP_mult_214_n674), .CI(
        DP_mult_214_n675), .CO(DP_mult_214_n671), .S(DP_mult_214_n672) );
  HA_X1 DP_mult_214_U399 ( .A(DP_mult_214_n852), .B(DP_mult_214_n1602), .CO(
        DP_mult_214_n669), .S(DP_mult_214_n670) );
  FA_X1 DP_mult_214_U398 ( .A(DP_mult_214_n875), .B(DP_mult_214_n670), .CI(
        DP_mult_214_n673), .CO(DP_mult_214_n667), .S(DP_mult_214_n668) );
  FA_X1 DP_mult_214_U397 ( .A(DP_mult_214_n898), .B(DP_mult_214_n668), .CI(
        DP_mult_214_n671), .CO(DP_mult_214_n665), .S(DP_mult_214_n666) );
  HA_X1 DP_mult_214_U396 ( .A(DP_mult_214_n669), .B(DP_mult_214_n851), .CO(
        DP_mult_214_n663), .S(DP_mult_214_n664) );
  FA_X1 DP_mult_214_U395 ( .A(DP_mult_214_n874), .B(DP_mult_214_n664), .CI(
        DP_mult_214_n667), .CO(DP_mult_214_n661), .S(DP_mult_214_n662) );
  FA_X1 DP_mult_214_U394 ( .A(DP_mult_214_n897), .B(DP_mult_214_n662), .CI(
        DP_mult_214_n665), .CO(DP_mult_214_n659), .S(DP_mult_214_n660) );
  HA_X1 DP_mult_214_U393 ( .A(DP_mult_214_n663), .B(DP_mult_214_n850), .CO(
        DP_mult_214_n657), .S(DP_mult_214_n658) );
  FA_X1 DP_mult_214_U392 ( .A(DP_mult_214_n873), .B(DP_mult_214_n658), .CI(
        DP_mult_214_n661), .CO(DP_mult_214_n655), .S(DP_mult_214_n656) );
  FA_X1 DP_mult_214_U391 ( .A(DP_mult_214_n896), .B(DP_mult_214_n656), .CI(
        DP_mult_214_n659), .CO(DP_mult_214_n653), .S(DP_mult_214_n654) );
  HA_X1 DP_mult_214_U390 ( .A(DP_mult_214_n826), .B(DP_mult_214_n1604), .CO(
        DP_mult_214_n651), .S(DP_mult_214_n652) );
  FA_X1 DP_mult_214_U389 ( .A(DP_mult_214_n849), .B(DP_mult_214_n652), .CI(
        DP_mult_214_n657), .CO(DP_mult_214_n649), .S(DP_mult_214_n650) );
  FA_X1 DP_mult_214_U388 ( .A(DP_mult_214_n872), .B(DP_mult_214_n650), .CI(
        DP_mult_214_n655), .CO(DP_mult_214_n647), .S(DP_mult_214_n648) );
  FA_X1 DP_mult_214_U387 ( .A(DP_mult_214_n895), .B(DP_mult_214_n648), .CI(
        DP_mult_214_n653), .CO(DP_mult_214_n645), .S(DP_mult_214_n646) );
  HA_X1 DP_mult_214_U386 ( .A(DP_mult_214_n651), .B(DP_mult_214_n825), .CO(
        DP_mult_214_n643), .S(DP_mult_214_n644) );
  FA_X1 DP_mult_214_U385 ( .A(DP_mult_214_n848), .B(DP_mult_214_n644), .CI(
        DP_mult_214_n649), .CO(DP_mult_214_n641), .S(DP_mult_214_n642) );
  FA_X1 DP_mult_214_U384 ( .A(DP_mult_214_n871), .B(DP_mult_214_n642), .CI(
        DP_mult_214_n647), .CO(DP_mult_214_n639), .S(DP_mult_214_n640) );
  FA_X1 DP_mult_214_U383 ( .A(DP_mult_214_n894), .B(DP_mult_214_n640), .CI(
        DP_mult_214_n645), .CO(DP_mult_214_n637), .S(DP_mult_214_n638) );
  HA_X1 DP_mult_214_U382 ( .A(DP_mult_214_n643), .B(DP_mult_214_n824), .CO(
        DP_mult_214_n635), .S(DP_mult_214_n636) );
  FA_X1 DP_mult_214_U381 ( .A(DP_mult_214_n847), .B(DP_mult_214_n636), .CI(
        DP_mult_214_n641), .CO(DP_mult_214_n633), .S(DP_mult_214_n634) );
  FA_X1 DP_mult_214_U380 ( .A(DP_mult_214_n870), .B(DP_mult_214_n634), .CI(
        DP_mult_214_n639), .CO(DP_mult_214_n631), .S(DP_mult_214_n632) );
  FA_X1 DP_mult_214_U379 ( .A(DP_mult_214_n893), .B(DP_mult_214_n632), .CI(
        DP_mult_214_n637), .CO(DP_mult_214_n629), .S(DP_mult_214_n630) );
  HA_X1 DP_mult_214_U378 ( .A(DP_mult_214_n800), .B(DP_mult_214_n1606), .CO(
        DP_mult_214_n627), .S(DP_mult_214_n628) );
  FA_X1 DP_mult_214_U377 ( .A(DP_mult_214_n823), .B(DP_mult_214_n628), .CI(
        DP_mult_214_n635), .CO(DP_mult_214_n625), .S(DP_mult_214_n626) );
  FA_X1 DP_mult_214_U376 ( .A(DP_mult_214_n846), .B(DP_mult_214_n626), .CI(
        DP_mult_214_n633), .CO(DP_mult_214_n623), .S(DP_mult_214_n624) );
  FA_X1 DP_mult_214_U375 ( .A(DP_mult_214_n869), .B(DP_mult_214_n624), .CI(
        DP_mult_214_n631), .CO(DP_mult_214_n621), .S(DP_mult_214_n622) );
  FA_X1 DP_mult_214_U374 ( .A(DP_mult_214_n892), .B(DP_mult_214_n622), .CI(
        DP_mult_214_n629), .CO(DP_mult_214_n619), .S(DP_mult_214_n620) );
  HA_X1 DP_mult_214_U373 ( .A(DP_mult_214_n627), .B(DP_mult_214_n799), .CO(
        DP_mult_214_n617), .S(DP_mult_214_n618) );
  FA_X1 DP_mult_214_U372 ( .A(DP_mult_214_n822), .B(DP_mult_214_n618), .CI(
        DP_mult_214_n625), .CO(DP_mult_214_n615), .S(DP_mult_214_n616) );
  FA_X1 DP_mult_214_U371 ( .A(DP_mult_214_n845), .B(DP_mult_214_n616), .CI(
        DP_mult_214_n623), .CO(DP_mult_214_n613), .S(DP_mult_214_n614) );
  FA_X1 DP_mult_214_U370 ( .A(DP_mult_214_n868), .B(DP_mult_214_n614), .CI(
        DP_mult_214_n621), .CO(DP_mult_214_n611), .S(DP_mult_214_n612) );
  FA_X1 DP_mult_214_U369 ( .A(DP_mult_214_n891), .B(DP_mult_214_n612), .CI(
        DP_mult_214_n619), .CO(DP_mult_214_n609), .S(DP_mult_214_n610) );
  HA_X1 DP_mult_214_U368 ( .A(DP_mult_214_n617), .B(DP_mult_214_n798), .CO(
        DP_mult_214_n607), .S(DP_mult_214_n608) );
  FA_X1 DP_mult_214_U367 ( .A(DP_mult_214_n821), .B(DP_mult_214_n608), .CI(
        DP_mult_214_n615), .CO(DP_mult_214_n605), .S(DP_mult_214_n606) );
  FA_X1 DP_mult_214_U366 ( .A(DP_mult_214_n844), .B(DP_mult_214_n606), .CI(
        DP_mult_214_n613), .CO(DP_mult_214_n603), .S(DP_mult_214_n604) );
  FA_X1 DP_mult_214_U365 ( .A(DP_mult_214_n867), .B(DP_mult_214_n604), .CI(
        DP_mult_214_n611), .CO(DP_mult_214_n601), .S(DP_mult_214_n602) );
  FA_X1 DP_mult_214_U364 ( .A(DP_mult_214_n890), .B(DP_mult_214_n602), .CI(
        DP_mult_214_n609), .CO(DP_mult_214_n599), .S(DP_mult_214_n600) );
  HA_X1 DP_mult_214_U363 ( .A(DP_mult_214_n774), .B(DP_mult_214_n1608), .CO(
        DP_mult_214_n597), .S(DP_mult_214_n598) );
  FA_X1 DP_mult_214_U362 ( .A(DP_mult_214_n797), .B(DP_mult_214_n598), .CI(
        DP_mult_214_n607), .CO(DP_mult_214_n595), .S(DP_mult_214_n596) );
  FA_X1 DP_mult_214_U361 ( .A(DP_mult_214_n820), .B(DP_mult_214_n596), .CI(
        DP_mult_214_n605), .CO(DP_mult_214_n593), .S(DP_mult_214_n594) );
  FA_X1 DP_mult_214_U360 ( .A(DP_mult_214_n843), .B(DP_mult_214_n594), .CI(
        DP_mult_214_n603), .CO(DP_mult_214_n591), .S(DP_mult_214_n592) );
  FA_X1 DP_mult_214_U359 ( .A(DP_mult_214_n866), .B(DP_mult_214_n592), .CI(
        DP_mult_214_n601), .CO(DP_mult_214_n589), .S(DP_mult_214_n590) );
  FA_X1 DP_mult_214_U358 ( .A(DP_mult_214_n889), .B(DP_mult_214_n590), .CI(
        DP_mult_214_n599), .CO(DP_mult_214_n587), .S(DP_mult_214_n588) );
  HA_X1 DP_mult_214_U357 ( .A(DP_mult_214_n597), .B(DP_mult_214_n773), .CO(
        DP_mult_214_n585), .S(DP_mult_214_n586) );
  FA_X1 DP_mult_214_U356 ( .A(DP_mult_214_n796), .B(DP_mult_214_n586), .CI(
        DP_mult_214_n595), .CO(DP_mult_214_n583), .S(DP_mult_214_n584) );
  FA_X1 DP_mult_214_U355 ( .A(DP_mult_214_n819), .B(DP_mult_214_n584), .CI(
        DP_mult_214_n593), .CO(DP_mult_214_n581), .S(DP_mult_214_n582) );
  FA_X1 DP_mult_214_U354 ( .A(DP_mult_214_n842), .B(DP_mult_214_n582), .CI(
        DP_mult_214_n591), .CO(DP_mult_214_n579), .S(DP_mult_214_n580) );
  FA_X1 DP_mult_214_U353 ( .A(DP_mult_214_n865), .B(DP_mult_214_n580), .CI(
        DP_mult_214_n589), .CO(DP_mult_214_n577), .S(DP_mult_214_n578) );
  FA_X1 DP_mult_214_U352 ( .A(DP_mult_214_n888), .B(DP_mult_214_n578), .CI(
        DP_mult_214_n587), .CO(DP_mult_214_n575), .S(DP_mult_214_n576) );
  HA_X1 DP_mult_214_U351 ( .A(DP_mult_214_n585), .B(DP_mult_214_n772), .CO(
        DP_mult_214_n573), .S(DP_mult_214_n574) );
  FA_X1 DP_mult_214_U350 ( .A(DP_mult_214_n795), .B(DP_mult_214_n574), .CI(
        DP_mult_214_n583), .CO(DP_mult_214_n571), .S(DP_mult_214_n572) );
  FA_X1 DP_mult_214_U349 ( .A(DP_mult_214_n818), .B(DP_mult_214_n572), .CI(
        DP_mult_214_n581), .CO(DP_mult_214_n569), .S(DP_mult_214_n570) );
  FA_X1 DP_mult_214_U348 ( .A(DP_mult_214_n841), .B(DP_mult_214_n570), .CI(
        DP_mult_214_n579), .CO(DP_mult_214_n567), .S(DP_mult_214_n568) );
  FA_X1 DP_mult_214_U347 ( .A(DP_mult_214_n864), .B(DP_mult_214_n568), .CI(
        DP_mult_214_n577), .CO(DP_mult_214_n565), .S(DP_mult_214_n566) );
  FA_X1 DP_mult_214_U346 ( .A(DP_mult_214_n887), .B(DP_mult_214_n566), .CI(
        DP_mult_214_n575), .CO(DP_mult_214_n563), .S(DP_mult_214_n564) );
  HA_X1 DP_mult_214_U345 ( .A(DP_mult_214_n748), .B(DP_mult_214_n1610), .CO(
        DP_mult_214_n561), .S(DP_mult_214_n562) );
  FA_X1 DP_mult_214_U344 ( .A(DP_mult_214_n771), .B(DP_mult_214_n562), .CI(
        DP_mult_214_n573), .CO(DP_mult_214_n559), .S(DP_mult_214_n560) );
  FA_X1 DP_mult_214_U343 ( .A(DP_mult_214_n794), .B(DP_mult_214_n560), .CI(
        DP_mult_214_n571), .CO(DP_mult_214_n557), .S(DP_mult_214_n558) );
  FA_X1 DP_mult_214_U342 ( .A(DP_mult_214_n817), .B(DP_mult_214_n558), .CI(
        DP_mult_214_n569), .CO(DP_mult_214_n555), .S(DP_mult_214_n556) );
  FA_X1 DP_mult_214_U341 ( .A(DP_mult_214_n840), .B(DP_mult_214_n556), .CI(
        DP_mult_214_n567), .CO(DP_mult_214_n553), .S(DP_mult_214_n554) );
  FA_X1 DP_mult_214_U340 ( .A(DP_mult_214_n863), .B(DP_mult_214_n554), .CI(
        DP_mult_214_n565), .CO(DP_mult_214_n551), .S(DP_mult_214_n552) );
  FA_X1 DP_mult_214_U339 ( .A(DP_mult_214_n886), .B(DP_mult_214_n552), .CI(
        DP_mult_214_n563), .CO(DP_mult_214_n549), .S(DP_mult_214_n550) );
  HA_X1 DP_mult_214_U338 ( .A(DP_mult_214_n561), .B(DP_mult_214_n747), .CO(
        DP_mult_214_n547), .S(DP_mult_214_n548) );
  FA_X1 DP_mult_214_U337 ( .A(DP_mult_214_n770), .B(DP_mult_214_n548), .CI(
        DP_mult_214_n559), .CO(DP_mult_214_n545), .S(DP_mult_214_n546) );
  FA_X1 DP_mult_214_U336 ( .A(DP_mult_214_n793), .B(DP_mult_214_n546), .CI(
        DP_mult_214_n557), .CO(DP_mult_214_n543), .S(DP_mult_214_n544) );
  FA_X1 DP_mult_214_U335 ( .A(DP_mult_214_n816), .B(DP_mult_214_n544), .CI(
        DP_mult_214_n555), .CO(DP_mult_214_n541), .S(DP_mult_214_n542) );
  FA_X1 DP_mult_214_U334 ( .A(DP_mult_214_n839), .B(DP_mult_214_n542), .CI(
        DP_mult_214_n553), .CO(DP_mult_214_n539), .S(DP_mult_214_n540) );
  FA_X1 DP_mult_214_U333 ( .A(DP_mult_214_n862), .B(DP_mult_214_n540), .CI(
        DP_mult_214_n551), .CO(DP_mult_214_n537), .S(DP_mult_214_n538) );
  FA_X1 DP_mult_214_U332 ( .A(DP_mult_214_n885), .B(DP_mult_214_n538), .CI(
        DP_mult_214_n549), .CO(DP_mult_214_n535), .S(DP_mult_214_n536) );
  HA_X1 DP_mult_214_U331 ( .A(DP_mult_214_n547), .B(DP_mult_214_n746), .CO(
        DP_mult_214_n533), .S(DP_mult_214_n534) );
  FA_X1 DP_mult_214_U330 ( .A(DP_mult_214_n769), .B(DP_mult_214_n534), .CI(
        DP_mult_214_n545), .CO(DP_mult_214_n531), .S(DP_mult_214_n532) );
  FA_X1 DP_mult_214_U329 ( .A(DP_mult_214_n792), .B(DP_mult_214_n532), .CI(
        DP_mult_214_n543), .CO(DP_mult_214_n529), .S(DP_mult_214_n530) );
  FA_X1 DP_mult_214_U328 ( .A(DP_mult_214_n815), .B(DP_mult_214_n530), .CI(
        DP_mult_214_n541), .CO(DP_mult_214_n527), .S(DP_mult_214_n528) );
  FA_X1 DP_mult_214_U327 ( .A(DP_mult_214_n838), .B(DP_mult_214_n528), .CI(
        DP_mult_214_n539), .CO(DP_mult_214_n525), .S(DP_mult_214_n526) );
  FA_X1 DP_mult_214_U326 ( .A(DP_mult_214_n861), .B(DP_mult_214_n526), .CI(
        DP_mult_214_n537), .CO(DP_mult_214_n523), .S(DP_mult_214_n524) );
  FA_X1 DP_mult_214_U325 ( .A(DP_mult_214_n884), .B(DP_mult_214_n524), .CI(
        DP_mult_214_n535), .CO(DP_mult_214_n521), .S(DP_mult_214_n522) );
  HA_X1 DP_mult_214_U324 ( .A(DP_mult_214_n533), .B(DP_mult_214_n745), .CO(
        DP_mult_214_n519), .S(DP_mult_214_n520) );
  FA_X1 DP_mult_214_U323 ( .A(DP_mult_214_n768), .B(DP_mult_214_n520), .CI(
        DP_mult_214_n531), .CO(DP_mult_214_n517), .S(DP_mult_214_n518) );
  FA_X1 DP_mult_214_U322 ( .A(DP_mult_214_n791), .B(DP_mult_214_n518), .CI(
        DP_mult_214_n529), .CO(DP_mult_214_n515), .S(DP_mult_214_n516) );
  FA_X1 DP_mult_214_U321 ( .A(DP_mult_214_n814), .B(DP_mult_214_n516), .CI(
        DP_mult_214_n527), .CO(DP_mult_214_n513), .S(DP_mult_214_n514) );
  FA_X1 DP_mult_214_U320 ( .A(DP_mult_214_n837), .B(DP_mult_214_n514), .CI(
        DP_mult_214_n525), .CO(DP_mult_214_n511), .S(DP_mult_214_n512) );
  FA_X1 DP_mult_214_U319 ( .A(DP_mult_214_n860), .B(DP_mult_214_n512), .CI(
        DP_mult_214_n523), .CO(DP_mult_214_n509), .S(DP_mult_214_n510) );
  FA_X1 DP_mult_214_U318 ( .A(DP_mult_214_n883), .B(DP_mult_214_n510), .CI(
        DP_mult_214_n521), .CO(DP_mult_214_n507), .S(DP_mult_214_n508) );
  FA_X1 DP_mult_214_U315 ( .A(DP_mult_214_n506), .B(DP_mult_214_n744), .CI(
        DP_mult_214_n767), .CO(DP_mult_214_n504), .S(DP_mult_214_n505) );
  FA_X1 DP_mult_214_U314 ( .A(DP_mult_214_n505), .B(DP_mult_214_n517), .CI(
        DP_mult_214_n790), .CO(DP_mult_214_n502), .S(DP_mult_214_n503) );
  FA_X1 DP_mult_214_U313 ( .A(DP_mult_214_n503), .B(DP_mult_214_n515), .CI(
        DP_mult_214_n813), .CO(DP_mult_214_n500), .S(DP_mult_214_n501) );
  FA_X1 DP_mult_214_U312 ( .A(DP_mult_214_n501), .B(DP_mult_214_n513), .CI(
        DP_mult_214_n836), .CO(DP_mult_214_n498), .S(DP_mult_214_n499) );
  FA_X1 DP_mult_214_U311 ( .A(DP_mult_214_n499), .B(DP_mult_214_n511), .CI(
        DP_mult_214_n859), .CO(DP_mult_214_n496), .S(DP_mult_214_n497) );
  FA_X1 DP_mult_214_U310 ( .A(DP_mult_214_n497), .B(DP_mult_214_n509), .CI(
        DP_mult_214_n882), .CO(DP_mult_214_n494), .S(DP_mult_214_n495) );
  FA_X1 DP_mult_214_U308 ( .A(DP_mult_214_n743), .B(DP_mult_214_n493), .CI(
        DP_mult_214_n766), .CO(DP_mult_214_n491), .S(DP_mult_214_n492) );
  FA_X1 DP_mult_214_U307 ( .A(DP_mult_214_n492), .B(DP_mult_214_n504), .CI(
        DP_mult_214_n789), .CO(DP_mult_214_n489), .S(DP_mult_214_n490) );
  FA_X1 DP_mult_214_U306 ( .A(DP_mult_214_n490), .B(DP_mult_214_n502), .CI(
        DP_mult_214_n500), .CO(DP_mult_214_n487), .S(DP_mult_214_n488) );
  FA_X1 DP_mult_214_U305 ( .A(DP_mult_214_n488), .B(DP_mult_214_n812), .CI(
        DP_mult_214_n835), .CO(DP_mult_214_n485), .S(DP_mult_214_n486) );
  FA_X1 DP_mult_214_U304 ( .A(DP_mult_214_n486), .B(DP_mult_214_n498), .CI(
        DP_mult_214_n496), .CO(DP_mult_214_n483), .S(DP_mult_214_n484) );
  FA_X1 DP_mult_214_U303 ( .A(DP_mult_214_n484), .B(DP_mult_214_n858), .CI(
        DP_mult_214_n881), .CO(DP_mult_214_n481), .S(DP_mult_214_n482) );
  FA_X1 DP_mult_214_U301 ( .A(DP_mult_214_n742), .B(DP_mult_214_n493), .CI(
        DP_mult_214_n491), .CO(DP_mult_214_n477), .S(DP_mult_214_n478) );
  FA_X1 DP_mult_214_U300 ( .A(DP_mult_214_n478), .B(DP_mult_214_n765), .CI(
        DP_mult_214_n788), .CO(DP_mult_214_n475), .S(DP_mult_214_n476) );
  FA_X1 DP_mult_214_U299 ( .A(DP_mult_214_n476), .B(DP_mult_214_n489), .CI(
        DP_mult_214_n487), .CO(DP_mult_214_n473), .S(DP_mult_214_n474) );
  FA_X1 DP_mult_214_U298 ( .A(DP_mult_214_n474), .B(DP_mult_214_n811), .CI(
        DP_mult_214_n834), .CO(DP_mult_214_n471), .S(DP_mult_214_n472) );
  FA_X1 DP_mult_214_U297 ( .A(DP_mult_214_n472), .B(DP_mult_214_n485), .CI(
        DP_mult_214_n483), .CO(DP_mult_214_n469), .S(DP_mult_214_n470) );
  FA_X1 DP_mult_214_U296 ( .A(DP_mult_214_n880), .B(DP_mult_214_n857), .CI(
        DP_mult_214_n470), .CO(DP_mult_214_n467), .S(DP_mult_214_n468) );
  FA_X1 DP_mult_214_U295 ( .A(DP_mult_214_n479), .B(DP_mult_214_n879), .CI(
        DP_mult_214_n741), .CO(DP_mult_214_n465), .S(DP_mult_214_n466) );
  FA_X1 DP_mult_214_U294 ( .A(DP_mult_214_n764), .B(DP_mult_214_n466), .CI(
        DP_mult_214_n477), .CO(DP_mult_214_n463), .S(DP_mult_214_n464) );
  FA_X1 DP_mult_214_U293 ( .A(DP_mult_214_n475), .B(DP_mult_214_n464), .CI(
        DP_mult_214_n787), .CO(DP_mult_214_n461), .S(DP_mult_214_n462) );
  FA_X1 DP_mult_214_U292 ( .A(DP_mult_214_n810), .B(DP_mult_214_n462), .CI(
        DP_mult_214_n473), .CO(DP_mult_214_n459), .S(DP_mult_214_n460) );
  FA_X1 DP_mult_214_U291 ( .A(DP_mult_214_n471), .B(DP_mult_214_n460), .CI(
        DP_mult_214_n833), .CO(DP_mult_214_n457), .S(DP_mult_214_n458) );
  FA_X1 DP_mult_214_U290 ( .A(DP_mult_214_n856), .B(DP_mult_214_n458), .CI(
        DP_mult_214_n469), .CO(DP_mult_214_n455), .S(DP_mult_214_n456) );
  FA_X1 DP_mult_214_U288 ( .A(DP_mult_214_n454), .B(DP_mult_214_n465), .CI(
        DP_mult_214_n763), .CO(DP_mult_214_n452), .S(DP_mult_214_n453) );
  FA_X1 DP_mult_214_U287 ( .A(DP_mult_214_n453), .B(DP_mult_214_n463), .CI(
        DP_mult_214_n786), .CO(DP_mult_214_n450), .S(DP_mult_214_n451) );
  FA_X1 DP_mult_214_U286 ( .A(DP_mult_214_n451), .B(DP_mult_214_n461), .CI(
        DP_mult_214_n809), .CO(DP_mult_214_n448), .S(DP_mult_214_n449) );
  FA_X1 DP_mult_214_U285 ( .A(DP_mult_214_n449), .B(DP_mult_214_n459), .CI(
        DP_mult_214_n832), .CO(DP_mult_214_n446), .S(DP_mult_214_n447) );
  FA_X1 DP_mult_214_U284 ( .A(DP_mult_214_n447), .B(DP_mult_214_n457), .CI(
        DP_mult_214_n855), .CO(DP_mult_214_n444), .S(DP_mult_214_n445) );
  FA_X1 DP_mult_214_U282 ( .A(DP_mult_214_n740), .B(DP_mult_214_n454), .CI(
        DP_mult_214_n762), .CO(DP_mult_214_n440), .S(DP_mult_214_n441) );
  FA_X1 DP_mult_214_U281 ( .A(DP_mult_214_n441), .B(DP_mult_214_n452), .CI(
        DP_mult_214_n450), .CO(DP_mult_214_n438), .S(DP_mult_214_n439) );
  FA_X1 DP_mult_214_U280 ( .A(DP_mult_214_n439), .B(DP_mult_214_n785), .CI(
        DP_mult_214_n808), .CO(DP_mult_214_n436), .S(DP_mult_214_n437) );
  FA_X1 DP_mult_214_U279 ( .A(DP_mult_214_n437), .B(DP_mult_214_n448), .CI(
        DP_mult_214_n446), .CO(DP_mult_214_n434), .S(DP_mult_214_n435) );
  FA_X1 DP_mult_214_U278 ( .A(DP_mult_214_n854), .B(DP_mult_214_n831), .CI(
        DP_mult_214_n435), .CO(DP_mult_214_n432), .S(DP_mult_214_n433) );
  FA_X1 DP_mult_214_U277 ( .A(DP_mult_214_n442), .B(DP_mult_214_n853), .CI(
        DP_mult_214_n739), .CO(DP_mult_214_n430), .S(DP_mult_214_n431) );
  FA_X1 DP_mult_214_U276 ( .A(DP_mult_214_n440), .B(DP_mult_214_n431), .CI(
        DP_mult_214_n761), .CO(DP_mult_214_n428), .S(DP_mult_214_n429) );
  FA_X1 DP_mult_214_U275 ( .A(DP_mult_214_n784), .B(DP_mult_214_n429), .CI(
        DP_mult_214_n438), .CO(DP_mult_214_n426), .S(DP_mult_214_n427) );
  FA_X1 DP_mult_214_U274 ( .A(DP_mult_214_n436), .B(DP_mult_214_n427), .CI(
        DP_mult_214_n807), .CO(DP_mult_214_n424), .S(DP_mult_214_n425) );
  FA_X1 DP_mult_214_U273 ( .A(DP_mult_214_n830), .B(DP_mult_214_n425), .CI(
        DP_mult_214_n434), .CO(DP_mult_214_n422), .S(DP_mult_214_n423) );
  FA_X1 DP_mult_214_U271 ( .A(DP_mult_214_n421), .B(DP_mult_214_n430), .CI(
        DP_mult_214_n760), .CO(DP_mult_214_n419), .S(DP_mult_214_n420) );
  FA_X1 DP_mult_214_U270 ( .A(DP_mult_214_n420), .B(DP_mult_214_n428), .CI(
        DP_mult_214_n783), .CO(DP_mult_214_n417), .S(DP_mult_214_n418) );
  FA_X1 DP_mult_214_U269 ( .A(DP_mult_214_n418), .B(DP_mult_214_n426), .CI(
        DP_mult_214_n806), .CO(DP_mult_214_n415), .S(DP_mult_214_n416) );
  FA_X1 DP_mult_214_U268 ( .A(DP_mult_214_n416), .B(DP_mult_214_n424), .CI(
        DP_mult_214_n829), .CO(DP_mult_214_n413), .S(DP_mult_214_n414) );
  FA_X1 DP_mult_214_U266 ( .A(DP_mult_214_n738), .B(DP_mult_214_n421), .CI(
        DP_mult_214_n419), .CO(DP_mult_214_n409), .S(DP_mult_214_n410) );
  FA_X1 DP_mult_214_U265 ( .A(DP_mult_214_n410), .B(DP_mult_214_n759), .CI(
        DP_mult_214_n782), .CO(DP_mult_214_n407), .S(DP_mult_214_n408) );
  FA_X1 DP_mult_214_U264 ( .A(DP_mult_214_n408), .B(DP_mult_214_n417), .CI(
        DP_mult_214_n415), .CO(DP_mult_214_n405), .S(DP_mult_214_n406) );
  FA_X1 DP_mult_214_U263 ( .A(DP_mult_214_n828), .B(DP_mult_214_n805), .CI(
        DP_mult_214_n406), .CO(DP_mult_214_n403), .S(DP_mult_214_n404) );
  FA_X1 DP_mult_214_U262 ( .A(DP_mult_214_n411), .B(DP_mult_214_n827), .CI(
        DP_mult_214_n737), .CO(DP_mult_214_n387), .S(DP_mult_214_n402) );
  FA_X1 DP_mult_214_U261 ( .A(DP_mult_214_n758), .B(DP_mult_214_n402), .CI(
        DP_mult_214_n409), .CO(DP_mult_214_n400), .S(DP_mult_214_n401) );
  FA_X1 DP_mult_214_U260 ( .A(DP_mult_214_n407), .B(DP_mult_214_n401), .CI(
        DP_mult_214_n781), .CO(DP_mult_214_n398), .S(DP_mult_214_n399) );
  FA_X1 DP_mult_214_U259 ( .A(DP_mult_214_n804), .B(DP_mult_214_n399), .CI(
        DP_mult_214_n405), .CO(DP_mult_214_n396), .S(DP_mult_214_n397) );
  FA_X1 DP_mult_214_U257 ( .A(DP_mult_214_n395), .B(DP_mult_214_n736), .CI(
        DP_mult_214_n757), .CO(DP_mult_214_n393), .S(DP_mult_214_n394) );
  FA_X1 DP_mult_214_U256 ( .A(DP_mult_214_n394), .B(DP_mult_214_n400), .CI(
        DP_mult_214_n780), .CO(DP_mult_214_n391), .S(DP_mult_214_n392) );
  FA_X1 DP_mult_214_U255 ( .A(DP_mult_214_n392), .B(DP_mult_214_n398), .CI(
        DP_mult_214_n803), .CO(DP_mult_214_n389), .S(DP_mult_214_n390) );
  FA_X1 DP_mult_214_U253 ( .A(DP_mult_214_n735), .B(DP_mult_214_n395), .CI(
        DP_mult_214_n756), .CO(DP_mult_214_n385), .S(DP_mult_214_n386) );
  FA_X1 DP_mult_214_U252 ( .A(DP_mult_214_n386), .B(DP_mult_214_n393), .CI(
        DP_mult_214_n391), .CO(DP_mult_214_n383), .S(DP_mult_214_n384) );
  FA_X1 DP_mult_214_U251 ( .A(DP_mult_214_n802), .B(DP_mult_214_n779), .CI(
        DP_mult_214_n384), .CO(DP_mult_214_n381), .S(DP_mult_214_n382) );
  FA_X1 DP_mult_214_U250 ( .A(DP_mult_214_n387), .B(DP_mult_214_n801), .CI(
        DP_mult_214_n734), .CO(DP_mult_214_n379), .S(DP_mult_214_n380) );
  FA_X1 DP_mult_214_U249 ( .A(DP_mult_214_n385), .B(DP_mult_214_n380), .CI(
        DP_mult_214_n755), .CO(DP_mult_214_n377), .S(DP_mult_214_n378) );
  FA_X1 DP_mult_214_U248 ( .A(DP_mult_214_n778), .B(DP_mult_214_n378), .CI(
        DP_mult_214_n383), .CO(DP_mult_214_n375), .S(DP_mult_214_n376) );
  FA_X1 DP_mult_214_U246 ( .A(DP_mult_214_n374), .B(DP_mult_214_n379), .CI(
        DP_mult_214_n754), .CO(DP_mult_214_n372), .S(DP_mult_214_n373) );
  FA_X1 DP_mult_214_U245 ( .A(DP_mult_214_n373), .B(DP_mult_214_n377), .CI(
        DP_mult_214_n777), .CO(DP_mult_214_n370), .S(DP_mult_214_n371) );
  FA_X1 DP_mult_214_U243 ( .A(DP_mult_214_n733), .B(DP_mult_214_n374), .CI(
        DP_mult_214_n372), .CO(DP_mult_214_n366), .S(DP_mult_214_n367) );
  FA_X1 DP_mult_214_U242 ( .A(DP_mult_214_n776), .B(DP_mult_214_n753), .CI(
        DP_mult_214_n367), .CO(DP_mult_214_n364), .S(DP_mult_214_n365) );
  FA_X1 DP_mult_214_U241 ( .A(DP_mult_214_n368), .B(DP_mult_214_n775), .CI(
        DP_mult_214_n732), .CO(DP_mult_214_n356), .S(DP_mult_214_n363) );
  FA_X1 DP_mult_214_U240 ( .A(DP_mult_214_n752), .B(DP_mult_214_n363), .CI(
        DP_mult_214_n366), .CO(DP_mult_214_n361), .S(DP_mult_214_n362) );
  FA_X1 DP_mult_214_U238 ( .A(DP_mult_214_n360), .B(DP_mult_214_n731), .CI(
        DP_mult_214_n751), .CO(DP_mult_214_n358), .S(DP_mult_214_n359) );
  FA_X1 DP_mult_214_U236 ( .A(DP_mult_214_n730), .B(DP_mult_214_n360), .CI(
        DP_mult_214_n750), .CO(DP_mult_214_n354), .S(DP_mult_214_n355) );
  FA_X1 DP_mult_214_U235 ( .A(DP_mult_214_n356), .B(DP_mult_214_n749), .CI(
        DP_mult_214_n729), .CO(DP_mult_214_n352), .S(DP_mult_214_n353) );
  FA_X1 DP_mult_214_U204 ( .A(DP_mult_214_n908), .B(DP_mult_214_n536), .CI(
        DP_mult_214_n326), .CO(DP_mult_214_n325), .S(DP_sw0_coeff_ret0[0]) );
  FA_X1 DP_mult_214_U203 ( .A(DP_mult_214_n907), .B(DP_mult_214_n522), .CI(
        DP_mult_214_n325), .CO(DP_mult_214_n324), .S(DP_sw0_coeff_ret0[1]) );
  FA_X1 DP_mult_214_U202 ( .A(DP_mult_214_n508), .B(DP_mult_214_n906), .CI(
        DP_mult_214_n324), .CO(DP_mult_214_n323), .S(DP_sw0_coeff_ret0[2]) );
  FA_X1 DP_mult_214_U201 ( .A(DP_mult_214_n495), .B(DP_mult_214_n507), .CI(
        DP_mult_214_n323), .CO(DP_mult_214_n322), .S(DP_sw0_coeff_ret0[3]) );
  FA_X1 DP_mult_214_U200 ( .A(DP_mult_214_n482), .B(DP_mult_214_n494), .CI(
        DP_mult_214_n322), .CO(DP_mult_214_n321), .S(DP_sw0_coeff_ret0[4]) );
  FA_X1 DP_mult_214_U199 ( .A(DP_mult_214_n468), .B(DP_mult_214_n481), .CI(
        DP_mult_214_n321), .CO(DP_mult_214_n320), .S(DP_sw0_coeff_ret0[5]) );
  FA_X1 DP_mult_214_U198 ( .A(DP_mult_214_n456), .B(DP_mult_214_n467), .CI(
        DP_mult_214_n320), .CO(DP_mult_214_n319), .S(DP_sw0_coeff_ret0[6]) );
  FA_X1 DP_mult_214_U197 ( .A(DP_mult_214_n445), .B(DP_mult_214_n455), .CI(
        DP_mult_214_n319), .CO(DP_mult_214_n318), .S(DP_sw0_coeff_ret0[7]) );
  FA_X1 DP_mult_214_U196 ( .A(DP_mult_214_n433), .B(DP_mult_214_n444), .CI(
        DP_mult_214_n318), .CO(DP_mult_214_n317), .S(DP_sw0_coeff_ret0[8]) );
  FA_X1 DP_mult_214_U195 ( .A(DP_mult_214_n423), .B(DP_mult_214_n432), .CI(
        DP_mult_214_n317), .CO(DP_mult_214_n316), .S(DP_sw0_coeff_ret0[9]) );
  FA_X1 DP_mult_214_U194 ( .A(DP_mult_214_n414), .B(DP_mult_214_n422), .CI(
        DP_mult_214_n316), .CO(DP_mult_214_n315), .S(DP_sw0_coeff_ret0[10]) );
  FA_X1 DP_mult_214_U193 ( .A(DP_mult_214_n404), .B(DP_mult_214_n413), .CI(
        DP_mult_214_n315), .CO(DP_mult_214_n314), .S(DP_sw0_coeff_ret0[11]) );
  FA_X1 DP_mult_214_U192 ( .A(DP_mult_214_n397), .B(DP_mult_214_n403), .CI(
        DP_mult_214_n314), .CO(DP_mult_214_n313), .S(DP_sw0_coeff_ret0[12]) );
  FA_X1 DP_mult_214_U191 ( .A(DP_mult_214_n390), .B(DP_mult_214_n396), .CI(
        DP_mult_214_n313), .CO(DP_mult_214_n312), .S(DP_sw0_coeff_ret0[13]) );
  FA_X1 DP_mult_214_U190 ( .A(DP_mult_214_n382), .B(DP_mult_214_n389), .CI(
        DP_mult_214_n312), .CO(DP_mult_214_n311), .S(DP_sw0_coeff_ret0[14]) );
  FA_X1 DP_mult_214_U189 ( .A(DP_mult_214_n376), .B(DP_mult_214_n381), .CI(
        DP_mult_214_n311), .CO(DP_mult_214_n310), .S(DP_sw0_coeff_ret0[15]) );
  FA_X1 DP_mult_214_U188 ( .A(DP_mult_214_n371), .B(DP_mult_214_n375), .CI(
        DP_mult_214_n310), .CO(DP_mult_214_n309), .S(DP_sw0_coeff_ret0[16]) );
  FA_X1 DP_mult_214_U187 ( .A(DP_mult_214_n365), .B(DP_mult_214_n370), .CI(
        DP_mult_214_n309), .CO(DP_mult_214_n308), .S(DP_sw0_coeff_ret0[17]) );
  FA_X1 DP_mult_214_U186 ( .A(DP_mult_214_n362), .B(DP_mult_214_n364), .CI(
        DP_mult_214_n308), .CO(DP_mult_214_n307), .S(DP_sw0_coeff_ret0[18]) );
  FA_X1 DP_mult_214_U185 ( .A(DP_mult_214_n359), .B(DP_mult_214_n361), .CI(
        DP_mult_214_n307), .CO(DP_mult_214_n306), .S(DP_sw0_coeff_ret0[19]) );
  FA_X1 DP_mult_214_U184 ( .A(DP_mult_214_n355), .B(DP_mult_214_n358), .CI(
        DP_mult_214_n306), .CO(DP_mult_214_n305), .S(DP_sw0_coeff_ret0[20]) );
  FA_X1 DP_mult_214_U183 ( .A(DP_mult_214_n353), .B(DP_mult_214_n354), .CI(
        DP_mult_214_n305), .CO(DP_mult_214_n304), .S(DP_sw0_coeff_ret0[21]) );
  FA_X1 DP_mult_214_U182 ( .A(DP_mult_214_n351), .B(DP_mult_214_n352), .CI(
        DP_mult_214_n304), .CO(DP_mult_214_n303), .S(DP_sw0_coeff_ret0[22]) );
  INV_X1 DP_mult_207_U237 ( .A(DP_mult_207_n1), .ZN(DP_N25) );
  INV_X1 DP_mult_207_U236 ( .A(DP_coeff_ret0[1]), .ZN(DP_mult_207_n244) );
  NOR2_X1 DP_mult_207_U235 ( .A1(DP_mult_207_n239), .A2(DP_mult_207_n244), 
        .ZN(DP_mult_207_n177) );
  NOR2_X1 DP_mult_207_U234 ( .A1(DP_mult_207_n244), .A2(DP_mult_207_n245), 
        .ZN(DP_mult_207_n176) );
  NOR2_X1 DP_mult_207_U233 ( .A1(DP_mult_207_n239), .A2(DP_mult_207_n245), 
        .ZN(DP_mult_207_n175) );
  INV_X1 DP_mult_207_U232 ( .A(DP_a_int_1__2_), .ZN(DP_mult_207_n245) );
  NOR2_X1 DP_mult_207_U231 ( .A1(DP_mult_207_n244), .A2(DP_mult_207_n240), 
        .ZN(DP_mult_207_n174) );
  NOR2_X1 DP_mult_207_U230 ( .A1(DP_mult_207_n239), .A2(DP_mult_207_n240), 
        .ZN(DP_mult_207_n173) );
  NOR2_X1 DP_mult_207_U229 ( .A1(DP_mult_207_n245), .A2(DP_mult_207_n240), 
        .ZN(DP_mult_207_n172) );
  NOR2_X1 DP_mult_207_U228 ( .A1(DP_mult_207_n244), .A2(DP_mult_207_n246), 
        .ZN(DP_mult_207_n171) );
  NOR2_X1 DP_mult_207_U227 ( .A1(DP_mult_207_n239), .A2(DP_mult_207_n246), 
        .ZN(DP_mult_207_n170) );
  NOR2_X1 DP_mult_207_U226 ( .A1(DP_mult_207_n245), .A2(DP_mult_207_n246), 
        .ZN(DP_mult_207_n169) );
  NOR2_X1 DP_mult_207_U225 ( .A1(DP_mult_207_n240), .A2(DP_mult_207_n246), 
        .ZN(DP_mult_207_n168) );
  INV_X1 DP_mult_207_U224 ( .A(DP_a_int_1__4_), .ZN(DP_mult_207_n246) );
  NOR2_X1 DP_mult_207_U223 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n244), 
        .ZN(DP_mult_207_n167) );
  NOR2_X1 DP_mult_207_U222 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n239), 
        .ZN(DP_mult_207_n166) );
  NOR2_X1 DP_mult_207_U221 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n245), 
        .ZN(DP_mult_207_n165) );
  NOR2_X1 DP_mult_207_U220 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n240), 
        .ZN(DP_mult_207_n164) );
  NOR2_X1 DP_mult_207_U219 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n246), 
        .ZN(DP_mult_207_n163) );
  NOR2_X1 DP_mult_207_U218 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n244), 
        .ZN(DP_mult_207_n162) );
  NOR2_X1 DP_mult_207_U217 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n239), 
        .ZN(DP_mult_207_n161) );
  NOR2_X1 DP_mult_207_U216 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n245), 
        .ZN(DP_mult_207_n160) );
  NOR2_X1 DP_mult_207_U215 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n240), 
        .ZN(DP_mult_207_n159) );
  NAND2_X1 DP_mult_207_U214 ( .A1(DP_a_int_1__6_), .A2(DP_mult_207_n241), .ZN(
        DP_mult_207_n71) );
  NOR2_X1 DP_mult_207_U213 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n246), 
        .ZN(DP_mult_207_n158) );
  INV_X1 DP_mult_207_U212 ( .A(DP_a_int_1__6_), .ZN(DP_mult_207_n247) );
  NOR2_X1 DP_mult_207_U211 ( .A1(DP_mult_207_n244), .A2(DP_mult_207_n242), 
        .ZN(DP_mult_207_n156) );
  NOR2_X1 DP_mult_207_U210 ( .A1(DP_mult_207_n239), .A2(DP_mult_207_n242), 
        .ZN(DP_mult_207_n155) );
  NOR2_X1 DP_mult_207_U209 ( .A1(DP_mult_207_n245), .A2(DP_mult_207_n242), 
        .ZN(DP_mult_207_n154) );
  NOR2_X1 DP_mult_207_U208 ( .A1(DP_mult_207_n240), .A2(DP_mult_207_n242), 
        .ZN(DP_mult_207_n153) );
  NOR2_X1 DP_mult_207_U207 ( .A1(DP_mult_207_n246), .A2(DP_mult_207_n242), 
        .ZN(DP_mult_207_n152) );
  NOR2_X1 DP_mult_207_U206 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n242), 
        .ZN(DP_mult_207_n151) );
  NOR2_X1 DP_mult_207_U205 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n242), 
        .ZN(DP_mult_207_n150) );
  NOR2_X1 DP_mult_207_U204 ( .A1(DP_mult_207_n244), .A2(DP_mult_207_n248), 
        .ZN(DP_mult_207_n149) );
  NOR2_X1 DP_mult_207_U203 ( .A1(DP_mult_207_n239), .A2(DP_mult_207_n248), 
        .ZN(DP_mult_207_n148) );
  NOR2_X1 DP_mult_207_U202 ( .A1(DP_mult_207_n245), .A2(DP_mult_207_n248), 
        .ZN(DP_mult_207_n147) );
  NOR2_X1 DP_mult_207_U201 ( .A1(DP_mult_207_n240), .A2(DP_mult_207_n248), 
        .ZN(DP_mult_207_n146) );
  NOR2_X1 DP_mult_207_U200 ( .A1(DP_mult_207_n246), .A2(DP_mult_207_n248), 
        .ZN(DP_mult_207_n145) );
  NOR2_X1 DP_mult_207_U199 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n248), 
        .ZN(DP_mult_207_n144) );
  NOR2_X1 DP_mult_207_U198 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n248), 
        .ZN(DP_mult_207_n143) );
  NOR2_X1 DP_mult_207_U197 ( .A1(DP_mult_207_n242), .A2(DP_mult_207_n248), 
        .ZN(DP_mult_207_n142) );
  INV_X1 DP_mult_207_U196 ( .A(DP_a_int_1__8_), .ZN(DP_mult_207_n248) );
  NOR2_X1 DP_mult_207_U195 ( .A1(DP_mult_207_n244), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n141) );
  NOR2_X1 DP_mult_207_U194 ( .A1(DP_mult_207_n245), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n139) );
  NOR2_X1 DP_mult_207_U193 ( .A1(DP_mult_207_n239), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n140) );
  NOR2_X1 DP_mult_207_U192 ( .A1(DP_mult_207_n240), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n138) );
  NOR2_X1 DP_mult_207_U191 ( .A1(DP_mult_207_n246), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n137) );
  NOR2_X1 DP_mult_207_U190 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n136) );
  NOR2_X1 DP_mult_207_U189 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n135) );
  NOR2_X1 DP_mult_207_U188 ( .A1(DP_mult_207_n242), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n134) );
  NOR2_X1 DP_mult_207_U187 ( .A1(DP_mult_207_n248), .A2(DP_mult_207_n243), 
        .ZN(DP_mult_207_n133) );
  NOR2_X1 DP_mult_207_U186 ( .A1(DP_mult_207_n239), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n131) );
  NOR2_X1 DP_mult_207_U185 ( .A1(DP_mult_207_n244), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n132) );
  NOR2_X1 DP_mult_207_U184 ( .A1(DP_mult_207_n245), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n130) );
  NOR2_X1 DP_mult_207_U183 ( .A1(DP_mult_207_n240), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n129) );
  NOR2_X1 DP_mult_207_U182 ( .A1(DP_mult_207_n246), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n128) );
  NOR2_X1 DP_mult_207_U181 ( .A1(DP_mult_207_n241), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n127) );
  NOR2_X1 DP_mult_207_U180 ( .A1(DP_mult_207_n247), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n126) );
  NOR2_X1 DP_mult_207_U179 ( .A1(DP_mult_207_n242), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n125) );
  NOR2_X1 DP_mult_207_U178 ( .A1(DP_mult_207_n248), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n124) );
  NOR2_X1 DP_mult_207_U177 ( .A1(DP_mult_207_n243), .A2(DP_mult_207_n249), 
        .ZN(DP_mult_207_n123) );
  INV_X1 DP_mult_207_U176 ( .A(DP_a_int_1__10_), .ZN(DP_mult_207_n249) );
  NAND2_X1 DP_mult_207_U175 ( .A1(DP_a_int_1__11_), .A2(DP_coeff_ret0[1]), 
        .ZN(DP_mult_207_n122) );
  NAND2_X1 DP_mult_207_U174 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__1_), .ZN(
        DP_mult_207_n121) );
  NAND2_X1 DP_mult_207_U173 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__2_), .ZN(
        DP_mult_207_n120) );
  NAND2_X1 DP_mult_207_U172 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__3_), .ZN(
        DP_mult_207_n119) );
  NAND2_X1 DP_mult_207_U171 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__4_), .ZN(
        DP_mult_207_n118) );
  NAND2_X1 DP_mult_207_U170 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__6_), .ZN(
        DP_mult_207_n116) );
  NAND2_X1 DP_mult_207_U169 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__5_), .ZN(
        DP_mult_207_n117) );
  NAND2_X1 DP_mult_207_U168 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__7_), .ZN(
        DP_mult_207_n115) );
  NAND2_X1 DP_mult_207_U167 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__9_), .ZN(
        DP_mult_207_n113) );
  NAND2_X1 DP_mult_207_U166 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__8_), .ZN(
        DP_mult_207_n114) );
  NAND2_X1 DP_mult_207_U165 ( .A1(DP_a_int_1__11_), .A2(DP_a_int_1__10_), .ZN(
        DP_mult_207_n112) );
  INV_X1 DP_mult_207_U164 ( .A(DP_a_int_1__9_), .ZN(DP_mult_207_n243) );
  INV_X1 DP_mult_207_U163 ( .A(DP_a_int_1__7_), .ZN(DP_mult_207_n242) );
  INV_X1 DP_mult_207_U162 ( .A(DP_a_int_1__5_), .ZN(DP_mult_207_n241) );
  INV_X1 DP_mult_207_U161 ( .A(DP_a_int_1__3_), .ZN(DP_mult_207_n240) );
  INV_X1 DP_mult_207_U160 ( .A(DP_a_int_1__1_), .ZN(DP_mult_207_n239) );
  FA_X1 DP_mult_207_U23 ( .A(DP_mult_207_n123), .B(DP_a_int_1__10_), .CI(
        DP_mult_207_n114), .CO(DP_mult_207_n22), .S(DP_mult_207_n23) );
  FA_X1 DP_mult_207_U24 ( .A(DP_mult_207_n115), .B(DP_mult_207_n124), .CI(
        DP_mult_207_n28), .CO(DP_mult_207_n24), .S(DP_mult_207_n25) );
  FA_X1 DP_mult_207_U28 ( .A(DP_mult_207_n126), .B(DP_mult_207_n134), .CI(
        DP_mult_207_n117), .CO(DP_mult_207_n32), .S(DP_mult_207_n33) );
  FA_X1 DP_mult_207_U25 ( .A(DP_mult_207_n32), .B(DP_mult_207_n116), .CI(
        DP_mult_207_n29), .CO(DP_mult_207_n26), .S(DP_mult_207_n27) );
  FA_X1 DP_mult_207_U30 ( .A(DP_mult_207_n118), .B(DP_mult_207_n127), .CI(
        DP_mult_207_n44), .CO(DP_mult_207_n36), .S(DP_mult_207_n37) );
  FA_X1 DP_mult_207_U27 ( .A(DP_mult_207_n33), .B(DP_mult_207_n38), .CI(
        DP_mult_207_n36), .CO(DP_mult_207_n30), .S(DP_mult_207_n31) );
  FA_X1 DP_mult_207_U37 ( .A(DP_mult_207_n129), .B(DP_mult_207_n137), .CI(
        DP_mult_207_n120), .CO(DP_mult_207_n50), .S(DP_mult_207_n51) );
  FA_X1 DP_mult_207_U33 ( .A(DP_mult_207_n52), .B(DP_mult_207_n119), .CI(
        DP_mult_207_n50), .CO(DP_mult_207_n42), .S(DP_mult_207_n43) );
  FA_X1 DP_mult_207_U29 ( .A(DP_mult_207_n42), .B(DP_mult_207_n39), .CI(
        DP_mult_207_n37), .CO(DP_mult_207_n34), .S(DP_mult_207_n35) );
  FA_X1 DP_mult_207_U41 ( .A(DP_mult_207_n121), .B(DP_mult_207_n145), .CI(
        DP_a_int_1__6_), .CO(DP_mult_207_n58), .S(DP_mult_207_n59) );
  FA_X1 DP_mult_207_U36 ( .A(DP_mult_207_n58), .B(DP_mult_207_n60), .CI(
        DP_mult_207_n53), .CO(DP_mult_207_n48), .S(DP_mult_207_n49) );
  FA_X1 DP_mult_207_U32 ( .A(DP_mult_207_n48), .B(DP_mult_207_n45), .CI(
        DP_mult_207_n43), .CO(DP_mult_207_n40), .S(DP_mult_207_n41) );
  FA_X1 DP_mult_207_U45 ( .A(DP_mult_207_n122), .B(DP_mult_207_n146), .CI(
        DP_mult_207_n78), .CO(DP_mult_207_n66), .S(DP_mult_207_n67) );
  FA_X1 DP_mult_207_U40 ( .A(DP_mult_207_n66), .B(DP_mult_207_n68), .CI(
        DP_mult_207_n61), .CO(DP_mult_207_n56), .S(DP_mult_207_n57) );
  FA_X1 DP_mult_207_U35 ( .A(DP_mult_207_n56), .B(DP_mult_207_n51), .CI(
        DP_mult_207_n49), .CO(DP_mult_207_n46), .S(DP_mult_207_n47) );
  FA_X1 DP_mult_207_U39 ( .A(DP_mult_207_n64), .B(DP_mult_207_n59), .CI(
        DP_mult_207_n57), .CO(DP_mult_207_n54), .S(DP_mult_207_n55) );
  FA_X1 DP_mult_207_U43 ( .A(DP_mult_207_n74), .B(DP_mult_207_n67), .CI(
        DP_mult_207_n65), .CO(DP_mult_207_n62), .S(DP_mult_207_n63) );
  FA_X1 DP_mult_207_U12 ( .A(DP_mult_207_n63), .B(DP_mult_207_n72), .CI(
        DP_mult_207_n12), .CO(DP_mult_207_n11), .S(DP_N14) );
  FA_X1 DP_mult_207_U11 ( .A(DP_mult_207_n55), .B(DP_mult_207_n62), .CI(
        DP_mult_207_n11), .CO(DP_mult_207_n10), .S(DP_N15) );
  FA_X1 DP_mult_207_U10 ( .A(DP_mult_207_n47), .B(DP_mult_207_n54), .CI(
        DP_mult_207_n10), .CO(DP_mult_207_n9), .S(DP_N16) );
  FA_X1 DP_mult_207_U9 ( .A(DP_mult_207_n41), .B(DP_mult_207_n46), .CI(
        DP_mult_207_n9), .CO(DP_mult_207_n8), .S(DP_N17) );
  FA_X1 DP_mult_207_U8 ( .A(DP_mult_207_n35), .B(DP_mult_207_n40), .CI(
        DP_mult_207_n8), .CO(DP_mult_207_n7), .S(DP_N18) );
  FA_X1 DP_mult_207_U7 ( .A(DP_mult_207_n31), .B(DP_mult_207_n34), .CI(
        DP_mult_207_n7), .CO(DP_mult_207_n6), .S(DP_N19) );
  FA_X1 DP_mult_207_U6 ( .A(DP_mult_207_n27), .B(DP_mult_207_n30), .CI(
        DP_mult_207_n6), .CO(DP_mult_207_n5), .S(DP_N20) );
  FA_X1 DP_mult_207_U5 ( .A(DP_mult_207_n25), .B(DP_mult_207_n26), .CI(
        DP_mult_207_n5), .CO(DP_mult_207_n4), .S(DP_N21) );
  FA_X1 DP_mult_207_U4 ( .A(DP_mult_207_n24), .B(DP_mult_207_n23), .CI(
        DP_mult_207_n4), .CO(DP_mult_207_n3), .S(DP_N22) );
  FA_X1 DP_mult_207_U3 ( .A(DP_mult_207_n22), .B(DP_mult_207_n113), .CI(
        DP_mult_207_n3), .CO(DP_mult_207_n2), .S(DP_N23) );
  FA_X1 DP_mult_207_U2 ( .A(DP_mult_207_n112), .B(DP_a_int_1__11_), .CI(
        DP_mult_207_n2), .CO(DP_mult_207_n1), .S(DP_N24) );
  FA_X1 DP_mult_207_U26 ( .A(DP_mult_207_n133), .B(DP_a_int_1__9_), .CI(
        DP_mult_207_n125), .CO(DP_mult_207_n28), .S(DP_mult_207_n29) );
  FA_X1 DP_mult_207_U34 ( .A(DP_mult_207_n128), .B(DP_mult_207_n143), .CI(
        DP_mult_207_n136), .CO(DP_mult_207_n44), .S(DP_mult_207_n45) );
  FA_X1 DP_mult_207_U42 ( .A(DP_mult_207_n130), .B(DP_mult_207_n151), .CI(
        DP_mult_207_n138), .CO(DP_mult_207_n60), .S(DP_mult_207_n61) );
  HA_X1 DP_mult_207_U52 ( .A(DP_mult_207_n132), .B(DP_mult_207_n140), .CO(
        DP_mult_207_n78), .S(DP_mult_207_n79) );
  FA_X1 DP_mult_207_U46 ( .A(DP_mult_207_n131), .B(DP_mult_207_n152), .CI(
        DP_mult_207_n139), .CO(DP_mult_207_n68), .S(DP_mult_207_n69) );
  FA_X1 DP_mult_207_U44 ( .A(DP_mult_207_n76), .B(DP_mult_207_n71), .CI(
        DP_mult_207_n69), .CO(DP_mult_207_n64), .S(DP_mult_207_n65) );
  FA_X1 DP_mult_207_U50 ( .A(DP_mult_207_n79), .B(DP_mult_207_n86), .CI(
        DP_mult_207_n84), .CO(DP_mult_207_n74), .S(DP_mult_207_n75) );
  FA_X1 DP_mult_207_U49 ( .A(DP_mult_207_n82), .B(DP_mult_207_n77), .CI(
        DP_mult_207_n75), .CO(DP_mult_207_n72), .S(DP_mult_207_n73) );
  FA_X1 DP_mult_207_U13 ( .A(DP_mult_207_n73), .B(DP_mult_207_n80), .CI(
        DP_mult_207_n13), .CO(DP_mult_207_n12), .S(DP_N13) );
  FA_X1 DP_mult_207_U31 ( .A(DP_mult_207_n142), .B(DP_a_int_1__8_), .CI(
        DP_mult_207_n135), .CO(DP_mult_207_n38), .S(DP_mult_207_n39) );
  FA_X1 DP_mult_207_U55 ( .A(DP_mult_207_n141), .B(DP_mult_207_n163), .CI(
        DP_mult_207_n154), .CO(DP_mult_207_n84), .S(DP_mult_207_n85) );
  FA_X1 DP_mult_207_U53 ( .A(DP_mult_207_n85), .B(DP_mult_207_n90), .CI(
        DP_mult_207_n83), .CO(DP_mult_207_n80), .S(DP_mult_207_n81) );
  FA_X1 DP_mult_207_U14 ( .A(DP_mult_207_n81), .B(DP_mult_207_n88), .CI(
        DP_mult_207_n14), .CO(DP_mult_207_n13), .S(DP_N12) );
  FA_X1 DP_mult_207_U38 ( .A(DP_mult_207_n150), .B(DP_a_int_1__7_), .CI(
        DP_mult_207_n144), .CO(DP_mult_207_n52), .S(DP_mult_207_n53) );
  FA_X1 DP_mult_207_U51 ( .A(DP_mult_207_n153), .B(DP_mult_207_n147), .CI(
        DP_mult_207_n158), .CO(DP_mult_207_n76), .S(DP_mult_207_n77) );
  HA_X1 DP_mult_207_U56 ( .A(DP_mult_207_n148), .B(DP_a_int_1__5_), .CO(
        DP_mult_207_n86), .S(DP_mult_207_n87) );
  HA_X1 DP_mult_207_U59 ( .A(DP_mult_207_n149), .B(DP_mult_207_n155), .CO(
        DP_mult_207_n92), .S(DP_mult_207_n93) );
  FA_X1 DP_mult_207_U54 ( .A(DP_mult_207_n92), .B(DP_mult_207_n159), .CI(
        DP_mult_207_n87), .CO(DP_mult_207_n82), .S(DP_mult_207_n83) );
  FA_X1 DP_mult_207_U57 ( .A(DP_mult_207_n96), .B(DP_mult_207_n93), .CI(
        DP_mult_207_n91), .CO(DP_mult_207_n88), .S(DP_mult_207_n89) );
  FA_X1 DP_mult_207_U15 ( .A(DP_mult_207_n89), .B(DP_mult_207_n94), .CI(
        DP_mult_207_n15), .CO(DP_mult_207_n14), .S(DP_N11) );
  FA_X1 DP_mult_207_U61 ( .A(DP_mult_207_n156), .B(DP_mult_207_n168), .CI(
        DP_mult_207_n165), .CO(DP_mult_207_n96), .S(DP_mult_207_n97) );
  FA_X1 DP_mult_207_U60 ( .A(DP_mult_207_n99), .B(DP_mult_207_n102), .CI(
        DP_mult_207_n97), .CO(DP_mult_207_n94), .S(DP_mult_207_n95) );
  FA_X1 DP_mult_207_U16 ( .A(DP_mult_207_n95), .B(DP_mult_207_n100), .CI(
        DP_mult_207_n16), .CO(DP_mult_207_n15), .S(DP_N10) );
  HA_X1 DP_mult_207_U62 ( .A(DP_mult_207_n161), .B(DP_a_int_1__4_), .CO(
        DP_mult_207_n98), .S(DP_mult_207_n99) );
  FA_X1 DP_mult_207_U58 ( .A(DP_mult_207_n160), .B(DP_mult_207_n164), .CI(
        DP_mult_207_n98), .CO(DP_mult_207_n90), .S(DP_mult_207_n91) );
  HA_X1 DP_mult_207_U64 ( .A(DP_mult_207_n162), .B(DP_mult_207_n169), .CO(
        DP_mult_207_n102), .S(DP_mult_207_n103) );
  FA_X1 DP_mult_207_U63 ( .A(DP_mult_207_n106), .B(DP_mult_207_n166), .CI(
        DP_mult_207_n103), .CO(DP_mult_207_n100), .S(DP_mult_207_n101) );
  FA_X1 DP_mult_207_U17 ( .A(DP_mult_207_n101), .B(DP_mult_207_n104), .CI(
        DP_mult_207_n17), .CO(DP_mult_207_n16), .S(DP_N9) );
  FA_X1 DP_mult_207_U65 ( .A(DP_mult_207_n167), .B(DP_mult_207_n170), .CI(
        DP_mult_207_n108), .CO(DP_mult_207_n104), .S(DP_mult_207_n105) );
  FA_X1 DP_mult_207_U18 ( .A(DP_mult_207_n105), .B(DP_mult_207_n107), .CI(
        DP_mult_207_n18), .CO(DP_mult_207_n17), .S(DP_N8) );
  HA_X1 DP_mult_207_U67 ( .A(DP_mult_207_n171), .B(DP_mult_207_n173), .CO(
        DP_mult_207_n108), .S(DP_mult_207_n109) );
  FA_X1 DP_mult_207_U19 ( .A(DP_mult_207_n109), .B(DP_mult_207_n110), .CI(
        DP_mult_207_n19), .CO(DP_mult_207_n18), .S(DP_N7) );
  HA_X1 DP_mult_207_U66 ( .A(DP_mult_207_n172), .B(DP_a_int_1__3_), .CO(
        DP_mult_207_n106), .S(DP_mult_207_n107) );
  FA_X1 DP_mult_207_U20 ( .A(DP_mult_207_n111), .B(DP_mult_207_n174), .CI(
        DP_mult_207_n20), .CO(DP_mult_207_n19), .S(DP_N6) );
  HA_X1 DP_mult_207_U68 ( .A(DP_mult_207_n175), .B(DP_a_int_1__2_), .CO(
        DP_mult_207_n110), .S(DP_mult_207_n111) );
  HA_X1 DP_mult_207_U21 ( .A(DP_mult_207_n21), .B(DP_mult_207_n176), .CO(
        DP_mult_207_n20), .S(DP_N5) );
  HA_X1 DP_mult_207_U22 ( .A(DP_mult_207_n177), .B(DP_a_int_1__1_), .CO(
        DP_mult_207_n21), .S(DP_N4) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U41 ( .A(DP_coeff_ret0[1]), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_2_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U40 ( .A(DP_N12), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_10_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U39 ( .A(DP_N13), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_11_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U38 ( .A(DP_N14), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_12_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U37 ( .A(DP_N15), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_13_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U36 ( .A(DP_N16), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_14_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U35 ( .A(DP_N17), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_15_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U34 ( .A(DP_N18), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_16_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U33 ( .A(DP_N19), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_17_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U32 ( .A(DP_N20), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_18_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U31 ( .A(DP_N21), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_19_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U30 ( .A(DP_N22), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_20_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U29 ( .A(DP_N23), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_21_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U28 ( .A(DP_N24), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_22_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U27 ( .A(DP_N25), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_23_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U26 ( .A(DP_N4), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_2_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U25 ( .A(DP_N5), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_3_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U24 ( .A(DP_N6), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_4_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U23 ( .A(DP_N7), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_5_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U22 ( .A(DP_N8), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_6_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U21 ( .A(DP_N9), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_7_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U20 ( .A(DP_N10), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_8_) );
  INV_X1 DP_sub_0_root_add_0_root_add_207_U19 ( .A(DP_N11), .ZN(
        DP_sub_0_root_add_0_root_add_207_B_not_9_) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U18 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_2_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_2_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_3_) );
  XOR2_X1 DP_sub_0_root_add_0_root_add_207_U17 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_3_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_3_), .Z(DP_coeff_ret0[3]) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U16 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_3_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_3_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_4_) );
  XOR2_X1 DP_sub_0_root_add_0_root_add_207_U15 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_4_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_4_), .Z(DP_coeff_ret0[4]) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U14 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_4_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_4_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_5_) );
  XOR2_X1 DP_sub_0_root_add_0_root_add_207_U13 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_5_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_5_), .Z(DP_coeff_ret0[5]) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U12 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_5_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_5_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_6_) );
  XOR2_X1 DP_sub_0_root_add_0_root_add_207_U11 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_6_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_6_), .Z(DP_coeff_ret0[6]) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U10 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_6_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_6_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_7_) );
  XOR2_X1 DP_sub_0_root_add_0_root_add_207_U9 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_7_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_7_), .Z(DP_coeff_ret0[7]) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U8 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_7_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_7_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_8_) );
  XOR2_X1 DP_sub_0_root_add_0_root_add_207_U7 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_8_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_8_), .Z(DP_coeff_ret0[8]) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U6 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_8_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_8_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_9_) );
  XOR2_X1 DP_sub_0_root_add_0_root_add_207_U5 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_9_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_9_), .Z(DP_coeff_ret0[9]) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U4 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_9_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_9_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_10_) );
  XOR2_X1 DP_sub_0_root_add_0_root_add_207_U3 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_10_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_10_), .Z(DP_coeff_ret0[10]) );
  AND2_X1 DP_sub_0_root_add_0_root_add_207_U2 ( .A1(
        DP_sub_0_root_add_0_root_add_207_carry_10_), .A2(
        DP_sub_0_root_add_0_root_add_207_B_not_10_), .ZN(
        DP_sub_0_root_add_0_root_add_207_carry_11_) );
  XOR2_X2 DP_sub_0_root_add_0_root_add_207_U1 ( .A(
        DP_sub_0_root_add_0_root_add_207_B_not_2_), .B(
        DP_sub_0_root_add_0_root_add_207_carry_2_), .Z(DP_coeff_ret0[2]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_11 ( .A(DP_N37), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_11_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_11_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_12_), .S(DP_coeff_ret0[11]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_12 ( .A(DP_N38), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_12_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_12_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_13_), .S(DP_coeff_ret0[12]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_13 ( .A(DP_N39), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_13_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_13_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_14_), .S(DP_coeff_ret0[13]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_14 ( .A(DP_N40), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_14_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_14_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_15_), .S(DP_coeff_ret0[14]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_15 ( .A(DP_N41), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_15_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_15_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_16_), .S(DP_coeff_ret0[15]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_16 ( .A(DP_N42), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_16_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_16_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_17_), .S(DP_coeff_ret0[16]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_17 ( .A(DP_N43), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_17_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_17_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_18_), .S(DP_coeff_ret0[17]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_18 ( .A(DP_N44), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_18_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_18_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_19_), .S(DP_coeff_ret0[18]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_19 ( .A(DP_N45), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_19_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_19_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_20_), .S(DP_coeff_ret0[19]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_20 ( .A(DP_N46), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_20_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_20_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_21_), .S(DP_coeff_ret0[20]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_21 ( .A(DP_N47), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_21_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_21_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_22_), .S(DP_coeff_ret0[21]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_22 ( .A(DP_N49), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_22_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_22_), .CO(
        DP_sub_0_root_add_0_root_add_207_carry_23_), .S(DP_coeff_ret0[22]) );
  FA_X1 DP_sub_0_root_add_0_root_add_207_U2_23 ( .A(DP_N49), .B(
        DP_sub_0_root_add_0_root_add_207_B_not_23_), .CI(
        DP_sub_0_root_add_0_root_add_207_carry_23_), .S(DP_coeff_ret0[23]) );
  XNOR2_X1 DP_mult_208_U520 ( .A(DP_N47), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n612) );
  XNOR2_X1 DP_mult_208_U519 ( .A(DP_mult_208_n524), .B(DP_a_int_1__10_), .ZN(
        DP_mult_208_n626) );
  NAND2_X1 DP_mult_208_U518 ( .A1(DP_mult_208_n600), .A2(DP_mult_208_n626), 
        .ZN(DP_mult_208_n602) );
  XNOR2_X1 DP_mult_208_U517 ( .A(DP_N49), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n614) );
  OAI22_X1 DP_mult_208_U516 ( .A1(DP_mult_208_n612), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n614), .ZN(DP_mult_208_n142) );
  INV_X1 DP_mult_208_U515 ( .A(DP_mult_208_n142), .ZN(DP_mult_208_n143) );
  XNOR2_X1 DP_mult_208_U514 ( .A(DP_N47), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n597) );
  XNOR2_X1 DP_mult_208_U513 ( .A(DP_mult_208_n522), .B(DP_a_int_1__8_), .ZN(
        DP_mult_208_n625) );
  NAND2_X1 DP_mult_208_U512 ( .A1(DP_mult_208_n585), .A2(DP_mult_208_n625), 
        .ZN(DP_mult_208_n587) );
  XNOR2_X1 DP_mult_208_U511 ( .A(DP_N49), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n599) );
  OAI22_X1 DP_mult_208_U510 ( .A1(DP_mult_208_n597), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n599), .ZN(DP_mult_208_n148) );
  INV_X1 DP_mult_208_U509 ( .A(DP_mult_208_n148), .ZN(DP_mult_208_n149) );
  XNOR2_X1 DP_mult_208_U508 ( .A(DP_N47), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n582) );
  XNOR2_X1 DP_mult_208_U507 ( .A(DP_mult_208_n520), .B(DP_a_int_1__6_), .ZN(
        DP_mult_208_n624) );
  NAND2_X1 DP_mult_208_U506 ( .A1(DP_mult_208_n570), .A2(DP_mult_208_n624), 
        .ZN(DP_mult_208_n572) );
  XNOR2_X1 DP_mult_208_U505 ( .A(DP_N49), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n584) );
  OAI22_X1 DP_mult_208_U504 ( .A1(DP_mult_208_n582), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n584), .ZN(DP_mult_208_n158) );
  INV_X1 DP_mult_208_U503 ( .A(DP_mult_208_n158), .ZN(DP_mult_208_n159) );
  XNOR2_X1 DP_mult_208_U502 ( .A(DP_N47), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n567) );
  XNOR2_X1 DP_mult_208_U501 ( .A(DP_mult_208_n518), .B(DP_a_int_1__4_), .ZN(
        DP_mult_208_n623) );
  NAND2_X1 DP_mult_208_U500 ( .A1(DP_mult_208_n555), .A2(DP_mult_208_n623), 
        .ZN(DP_mult_208_n557) );
  XNOR2_X1 DP_mult_208_U499 ( .A(DP_N49), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n569) );
  OAI22_X1 DP_mult_208_U498 ( .A1(DP_mult_208_n567), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n569), .ZN(DP_mult_208_n172) );
  INV_X1 DP_mult_208_U497 ( .A(DP_mult_208_n172), .ZN(DP_mult_208_n173) );
  XNOR2_X1 DP_mult_208_U496 ( .A(DP_N47), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n552) );
  XNOR2_X1 DP_mult_208_U495 ( .A(DP_mult_208_n516), .B(DP_a_int_1__2_), .ZN(
        DP_mult_208_n622) );
  NAND2_X1 DP_mult_208_U494 ( .A1(DP_mult_208_n540), .A2(DP_mult_208_n622), 
        .ZN(DP_mult_208_n542) );
  XNOR2_X1 DP_mult_208_U493 ( .A(DP_N49), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n554) );
  OAI22_X1 DP_mult_208_U492 ( .A1(DP_mult_208_n552), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n554), .ZN(DP_mult_208_n190) );
  INV_X1 DP_mult_208_U491 ( .A(DP_mult_208_n190), .ZN(DP_mult_208_n191) );
  XNOR2_X1 DP_mult_208_U490 ( .A(DP_N40), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n590) );
  XNOR2_X1 DP_mult_208_U489 ( .A(DP_N41), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n591) );
  OAI22_X1 DP_mult_208_U488 ( .A1(DP_mult_208_n590), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n591), .ZN(DP_mult_208_n620) );
  XNOR2_X1 DP_mult_208_U487 ( .A(DP_N44), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n564) );
  XNOR2_X1 DP_mult_208_U486 ( .A(DP_N45), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n565) );
  OAI22_X1 DP_mult_208_U485 ( .A1(DP_mult_208_n564), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n565), .ZN(DP_mult_208_n621) );
  OR2_X1 DP_mult_208_U484 ( .A1(DP_mult_208_n620), .A2(DP_mult_208_n621), .ZN(
        DP_mult_208_n200) );
  XNOR2_X1 DP_mult_208_U483 ( .A(DP_mult_208_n620), .B(DP_mult_208_n621), .ZN(
        DP_mult_208_n201) );
  OR3_X1 DP_mult_208_U482 ( .A1(DP_mult_208_n600), .A2(DP_N37), .A3(
        DP_mult_208_n524), .ZN(DP_mult_208_n619) );
  OAI21_X1 DP_mult_208_U481 ( .B1(DP_mult_208_n524), .B2(DP_mult_208_n602), 
        .A(DP_mult_208_n619), .ZN(DP_mult_208_n252) );
  OR3_X1 DP_mult_208_U480 ( .A1(DP_mult_208_n585), .A2(DP_N37), .A3(
        DP_mult_208_n522), .ZN(DP_mult_208_n618) );
  OAI21_X1 DP_mult_208_U479 ( .B1(DP_mult_208_n522), .B2(DP_mult_208_n587), 
        .A(DP_mult_208_n618), .ZN(DP_mult_208_n253) );
  OR3_X1 DP_mult_208_U478 ( .A1(DP_mult_208_n570), .A2(DP_N37), .A3(
        DP_mult_208_n520), .ZN(DP_mult_208_n617) );
  OAI21_X1 DP_mult_208_U477 ( .B1(DP_mult_208_n520), .B2(DP_mult_208_n572), 
        .A(DP_mult_208_n617), .ZN(DP_mult_208_n254) );
  OR3_X1 DP_mult_208_U476 ( .A1(DP_mult_208_n555), .A2(DP_N37), .A3(
        DP_mult_208_n518), .ZN(DP_mult_208_n616) );
  OAI21_X1 DP_mult_208_U475 ( .B1(DP_mult_208_n518), .B2(DP_mult_208_n557), 
        .A(DP_mult_208_n616), .ZN(DP_mult_208_n255) );
  OR3_X1 DP_mult_208_U474 ( .A1(DP_mult_208_n540), .A2(DP_N37), .A3(
        DP_mult_208_n516), .ZN(DP_mult_208_n615) );
  OAI21_X1 DP_mult_208_U473 ( .B1(DP_mult_208_n516), .B2(DP_mult_208_n542), 
        .A(DP_mult_208_n615), .ZN(DP_mult_208_n256) );
  INV_X1 DP_mult_208_U472 ( .A(DP_coeff_ret0[1]), .ZN(DP_mult_208_n526) );
  NAND2_X1 DP_mult_208_U471 ( .A1(DP_mult_208_n513), .A2(DP_mult_208_n526), 
        .ZN(DP_mult_208_n527) );
  OAI21_X1 DP_mult_208_U470 ( .B1(DP_N37), .B2(DP_mult_208_n514), .A(
        DP_mult_208_n527), .ZN(DP_mult_208_n257) );
  AOI21_X1 DP_mult_208_U469 ( .B1(DP_mult_208_n602), .B2(DP_mult_208_n600), 
        .A(DP_mult_208_n614), .ZN(DP_mult_208_n613) );
  INV_X1 DP_mult_208_U468 ( .A(DP_mult_208_n613), .ZN(DP_mult_208_n258) );
  XNOR2_X1 DP_mult_208_U467 ( .A(DP_N46), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n611) );
  OAI22_X1 DP_mult_208_U466 ( .A1(DP_mult_208_n611), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n612), .ZN(DP_mult_208_n259) );
  XNOR2_X1 DP_mult_208_U465 ( .A(DP_N45), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n610) );
  OAI22_X1 DP_mult_208_U464 ( .A1(DP_mult_208_n610), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n611), .ZN(DP_mult_208_n260) );
  XNOR2_X1 DP_mult_208_U463 ( .A(DP_N44), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n609) );
  OAI22_X1 DP_mult_208_U462 ( .A1(DP_mult_208_n609), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n610), .ZN(DP_mult_208_n261) );
  XNOR2_X1 DP_mult_208_U461 ( .A(DP_N43), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n608) );
  OAI22_X1 DP_mult_208_U460 ( .A1(DP_mult_208_n608), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n609), .ZN(DP_mult_208_n262) );
  XNOR2_X1 DP_mult_208_U459 ( .A(DP_N42), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n607) );
  OAI22_X1 DP_mult_208_U458 ( .A1(DP_mult_208_n607), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n608), .ZN(DP_mult_208_n263) );
  XNOR2_X1 DP_mult_208_U457 ( .A(DP_N41), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n606) );
  OAI22_X1 DP_mult_208_U456 ( .A1(DP_mult_208_n606), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n607), .ZN(DP_mult_208_n264) );
  XNOR2_X1 DP_mult_208_U455 ( .A(DP_N40), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n605) );
  OAI22_X1 DP_mult_208_U454 ( .A1(DP_mult_208_n605), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n606), .ZN(DP_mult_208_n265) );
  XNOR2_X1 DP_mult_208_U453 ( .A(DP_N39), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n604) );
  OAI22_X1 DP_mult_208_U452 ( .A1(DP_mult_208_n604), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n605), .ZN(DP_mult_208_n266) );
  XNOR2_X1 DP_mult_208_U451 ( .A(DP_N38), .B(DP_mult_208_n523), .ZN(
        DP_mult_208_n603) );
  OAI22_X1 DP_mult_208_U450 ( .A1(DP_mult_208_n603), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n604), .ZN(DP_mult_208_n267) );
  XNOR2_X1 DP_mult_208_U449 ( .A(DP_mult_208_n523), .B(DP_N37), .ZN(
        DP_mult_208_n601) );
  OAI22_X1 DP_mult_208_U448 ( .A1(DP_mult_208_n601), .A2(DP_mult_208_n602), 
        .B1(DP_mult_208_n600), .B2(DP_mult_208_n603), .ZN(DP_mult_208_n268) );
  INV_X1 DP_mult_208_U447 ( .A(DP_N37), .ZN(DP_mult_208_n525) );
  NOR2_X1 DP_mult_208_U446 ( .A1(DP_mult_208_n525), .A2(DP_mult_208_n600), 
        .ZN(DP_mult_208_n269) );
  AOI21_X1 DP_mult_208_U445 ( .B1(DP_mult_208_n587), .B2(DP_mult_208_n585), 
        .A(DP_mult_208_n599), .ZN(DP_mult_208_n598) );
  INV_X1 DP_mult_208_U444 ( .A(DP_mult_208_n598), .ZN(DP_mult_208_n270) );
  XNOR2_X1 DP_mult_208_U443 ( .A(DP_N46), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n596) );
  OAI22_X1 DP_mult_208_U442 ( .A1(DP_mult_208_n596), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n597), .ZN(DP_mult_208_n271) );
  XNOR2_X1 DP_mult_208_U441 ( .A(DP_N45), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n595) );
  OAI22_X1 DP_mult_208_U440 ( .A1(DP_mult_208_n595), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n596), .ZN(DP_mult_208_n272) );
  XNOR2_X1 DP_mult_208_U439 ( .A(DP_N44), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n594) );
  OAI22_X1 DP_mult_208_U438 ( .A1(DP_mult_208_n594), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n595), .ZN(DP_mult_208_n273) );
  XNOR2_X1 DP_mult_208_U437 ( .A(DP_N43), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n593) );
  OAI22_X1 DP_mult_208_U436 ( .A1(DP_mult_208_n593), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n594), .ZN(DP_mult_208_n274) );
  XNOR2_X1 DP_mult_208_U435 ( .A(DP_N42), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n592) );
  OAI22_X1 DP_mult_208_U434 ( .A1(DP_mult_208_n592), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n593), .ZN(DP_mult_208_n275) );
  OAI22_X1 DP_mult_208_U433 ( .A1(DP_mult_208_n591), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n592), .ZN(DP_mult_208_n276) );
  XNOR2_X1 DP_mult_208_U432 ( .A(DP_N39), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n589) );
  OAI22_X1 DP_mult_208_U431 ( .A1(DP_mult_208_n589), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n590), .ZN(DP_mult_208_n278) );
  XNOR2_X1 DP_mult_208_U430 ( .A(DP_N38), .B(DP_mult_208_n521), .ZN(
        DP_mult_208_n588) );
  OAI22_X1 DP_mult_208_U429 ( .A1(DP_mult_208_n588), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n589), .ZN(DP_mult_208_n279) );
  XNOR2_X1 DP_mult_208_U428 ( .A(DP_mult_208_n521), .B(DP_N37), .ZN(
        DP_mult_208_n586) );
  OAI22_X1 DP_mult_208_U427 ( .A1(DP_mult_208_n586), .A2(DP_mult_208_n587), 
        .B1(DP_mult_208_n585), .B2(DP_mult_208_n588), .ZN(DP_mult_208_n280) );
  NOR2_X1 DP_mult_208_U426 ( .A1(DP_mult_208_n525), .A2(DP_mult_208_n585), 
        .ZN(DP_mult_208_n281) );
  AOI21_X1 DP_mult_208_U425 ( .B1(DP_mult_208_n572), .B2(DP_mult_208_n570), 
        .A(DP_mult_208_n584), .ZN(DP_mult_208_n583) );
  INV_X1 DP_mult_208_U424 ( .A(DP_mult_208_n583), .ZN(DP_mult_208_n282) );
  XNOR2_X1 DP_mult_208_U423 ( .A(DP_N46), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n581) );
  OAI22_X1 DP_mult_208_U422 ( .A1(DP_mult_208_n581), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n582), .ZN(DP_mult_208_n283) );
  XNOR2_X1 DP_mult_208_U421 ( .A(DP_N45), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n580) );
  OAI22_X1 DP_mult_208_U420 ( .A1(DP_mult_208_n580), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n581), .ZN(DP_mult_208_n284) );
  XNOR2_X1 DP_mult_208_U419 ( .A(DP_N44), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n579) );
  OAI22_X1 DP_mult_208_U418 ( .A1(DP_mult_208_n579), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n580), .ZN(DP_mult_208_n285) );
  XNOR2_X1 DP_mult_208_U417 ( .A(DP_N43), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n578) );
  OAI22_X1 DP_mult_208_U416 ( .A1(DP_mult_208_n578), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n579), .ZN(DP_mult_208_n286) );
  XNOR2_X1 DP_mult_208_U415 ( .A(DP_N42), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n577) );
  OAI22_X1 DP_mult_208_U414 ( .A1(DP_mult_208_n577), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n578), .ZN(DP_mult_208_n287) );
  XNOR2_X1 DP_mult_208_U413 ( .A(DP_N41), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n576) );
  OAI22_X1 DP_mult_208_U412 ( .A1(DP_mult_208_n576), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n577), .ZN(DP_mult_208_n288) );
  XNOR2_X1 DP_mult_208_U411 ( .A(DP_N40), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n575) );
  OAI22_X1 DP_mult_208_U410 ( .A1(DP_mult_208_n575), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n576), .ZN(DP_mult_208_n289) );
  XNOR2_X1 DP_mult_208_U409 ( .A(DP_N39), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n574) );
  OAI22_X1 DP_mult_208_U408 ( .A1(DP_mult_208_n574), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n575), .ZN(DP_mult_208_n290) );
  XNOR2_X1 DP_mult_208_U407 ( .A(DP_N38), .B(DP_mult_208_n519), .ZN(
        DP_mult_208_n573) );
  OAI22_X1 DP_mult_208_U406 ( .A1(DP_mult_208_n573), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n574), .ZN(DP_mult_208_n291) );
  XNOR2_X1 DP_mult_208_U405 ( .A(DP_mult_208_n519), .B(DP_N37), .ZN(
        DP_mult_208_n571) );
  OAI22_X1 DP_mult_208_U404 ( .A1(DP_mult_208_n571), .A2(DP_mult_208_n572), 
        .B1(DP_mult_208_n570), .B2(DP_mult_208_n573), .ZN(DP_mult_208_n292) );
  NOR2_X1 DP_mult_208_U403 ( .A1(DP_mult_208_n525), .A2(DP_mult_208_n570), 
        .ZN(DP_mult_208_n293) );
  AOI21_X1 DP_mult_208_U402 ( .B1(DP_mult_208_n557), .B2(DP_mult_208_n555), 
        .A(DP_mult_208_n569), .ZN(DP_mult_208_n568) );
  INV_X1 DP_mult_208_U401 ( .A(DP_mult_208_n568), .ZN(DP_mult_208_n294) );
  XNOR2_X1 DP_mult_208_U400 ( .A(DP_N46), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n566) );
  OAI22_X1 DP_mult_208_U399 ( .A1(DP_mult_208_n566), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n567), .ZN(DP_mult_208_n295) );
  OAI22_X1 DP_mult_208_U398 ( .A1(DP_mult_208_n565), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n566), .ZN(DP_mult_208_n296) );
  XNOR2_X1 DP_mult_208_U397 ( .A(DP_N43), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n563) );
  OAI22_X1 DP_mult_208_U396 ( .A1(DP_mult_208_n563), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n564), .ZN(DP_mult_208_n298) );
  XNOR2_X1 DP_mult_208_U395 ( .A(DP_N42), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n562) );
  OAI22_X1 DP_mult_208_U394 ( .A1(DP_mult_208_n562), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n563), .ZN(DP_mult_208_n299) );
  XNOR2_X1 DP_mult_208_U393 ( .A(DP_N41), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n561) );
  OAI22_X1 DP_mult_208_U392 ( .A1(DP_mult_208_n561), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n562), .ZN(DP_mult_208_n300) );
  XNOR2_X1 DP_mult_208_U391 ( .A(DP_N40), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n560) );
  OAI22_X1 DP_mult_208_U390 ( .A1(DP_mult_208_n560), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n561), .ZN(DP_mult_208_n301) );
  XNOR2_X1 DP_mult_208_U389 ( .A(DP_N39), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n559) );
  OAI22_X1 DP_mult_208_U388 ( .A1(DP_mult_208_n559), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n560), .ZN(DP_mult_208_n302) );
  XNOR2_X1 DP_mult_208_U387 ( .A(DP_N38), .B(DP_mult_208_n517), .ZN(
        DP_mult_208_n558) );
  OAI22_X1 DP_mult_208_U386 ( .A1(DP_mult_208_n558), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n559), .ZN(DP_mult_208_n303) );
  XNOR2_X1 DP_mult_208_U385 ( .A(DP_mult_208_n517), .B(DP_N37), .ZN(
        DP_mult_208_n556) );
  OAI22_X1 DP_mult_208_U384 ( .A1(DP_mult_208_n556), .A2(DP_mult_208_n557), 
        .B1(DP_mult_208_n555), .B2(DP_mult_208_n558), .ZN(DP_mult_208_n304) );
  NOR2_X1 DP_mult_208_U383 ( .A1(DP_mult_208_n525), .A2(DP_mult_208_n555), 
        .ZN(DP_mult_208_n305) );
  AOI21_X1 DP_mult_208_U382 ( .B1(DP_mult_208_n542), .B2(DP_mult_208_n540), 
        .A(DP_mult_208_n554), .ZN(DP_mult_208_n553) );
  INV_X1 DP_mult_208_U381 ( .A(DP_mult_208_n553), .ZN(DP_mult_208_n306) );
  XNOR2_X1 DP_mult_208_U380 ( .A(DP_N46), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n551) );
  OAI22_X1 DP_mult_208_U379 ( .A1(DP_mult_208_n551), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n552), .ZN(DP_mult_208_n307) );
  XNOR2_X1 DP_mult_208_U378 ( .A(DP_N45), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n550) );
  OAI22_X1 DP_mult_208_U377 ( .A1(DP_mult_208_n550), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n551), .ZN(DP_mult_208_n308) );
  XNOR2_X1 DP_mult_208_U376 ( .A(DP_N44), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n549) );
  OAI22_X1 DP_mult_208_U375 ( .A1(DP_mult_208_n549), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n550), .ZN(DP_mult_208_n309) );
  XNOR2_X1 DP_mult_208_U374 ( .A(DP_N43), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n548) );
  OAI22_X1 DP_mult_208_U373 ( .A1(DP_mult_208_n548), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n549), .ZN(DP_mult_208_n310) );
  XNOR2_X1 DP_mult_208_U372 ( .A(DP_N42), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n547) );
  OAI22_X1 DP_mult_208_U371 ( .A1(DP_mult_208_n547), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n548), .ZN(DP_mult_208_n311) );
  XNOR2_X1 DP_mult_208_U370 ( .A(DP_N41), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n546) );
  OAI22_X1 DP_mult_208_U369 ( .A1(DP_mult_208_n546), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n547), .ZN(DP_mult_208_n312) );
  XNOR2_X1 DP_mult_208_U368 ( .A(DP_N40), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n545) );
  OAI22_X1 DP_mult_208_U367 ( .A1(DP_mult_208_n545), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n546), .ZN(DP_mult_208_n313) );
  XNOR2_X1 DP_mult_208_U366 ( .A(DP_N39), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n544) );
  OAI22_X1 DP_mult_208_U365 ( .A1(DP_mult_208_n544), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n545), .ZN(DP_mult_208_n314) );
  XNOR2_X1 DP_mult_208_U364 ( .A(DP_N38), .B(DP_mult_208_n515), .ZN(
        DP_mult_208_n543) );
  OAI22_X1 DP_mult_208_U363 ( .A1(DP_mult_208_n543), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n544), .ZN(DP_mult_208_n315) );
  XNOR2_X1 DP_mult_208_U362 ( .A(DP_mult_208_n515), .B(DP_N37), .ZN(
        DP_mult_208_n541) );
  OAI22_X1 DP_mult_208_U361 ( .A1(DP_mult_208_n541), .A2(DP_mult_208_n542), 
        .B1(DP_mult_208_n540), .B2(DP_mult_208_n543), .ZN(DP_mult_208_n316) );
  NOR2_X1 DP_mult_208_U360 ( .A1(DP_mult_208_n525), .A2(DP_mult_208_n540), 
        .ZN(DP_mult_208_n317) );
  XNOR2_X1 DP_mult_208_U359 ( .A(DP_N49), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n538) );
  AOI21_X1 DP_mult_208_U358 ( .B1(DP_mult_208_n527), .B2(DP_mult_208_n526), 
        .A(DP_mult_208_n538), .ZN(DP_mult_208_n539) );
  INV_X1 DP_mult_208_U357 ( .A(DP_mult_208_n539), .ZN(DP_mult_208_n318) );
  XNOR2_X1 DP_mult_208_U356 ( .A(DP_N47), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n537) );
  OAI22_X1 DP_mult_208_U355 ( .A1(DP_mult_208_n537), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n538), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n319) );
  XNOR2_X1 DP_mult_208_U354 ( .A(DP_N46), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n536) );
  OAI22_X1 DP_mult_208_U353 ( .A1(DP_mult_208_n536), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n537), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n320) );
  XNOR2_X1 DP_mult_208_U352 ( .A(DP_N45), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n535) );
  OAI22_X1 DP_mult_208_U351 ( .A1(DP_mult_208_n535), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n536), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n321) );
  XNOR2_X1 DP_mult_208_U350 ( .A(DP_N44), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n534) );
  OAI22_X1 DP_mult_208_U349 ( .A1(DP_mult_208_n534), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n535), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n322) );
  XNOR2_X1 DP_mult_208_U348 ( .A(DP_N43), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n533) );
  OAI22_X1 DP_mult_208_U347 ( .A1(DP_mult_208_n533), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n534), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n323) );
  XNOR2_X1 DP_mult_208_U346 ( .A(DP_N42), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n532) );
  OAI22_X1 DP_mult_208_U345 ( .A1(DP_mult_208_n532), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n533), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n324) );
  XNOR2_X1 DP_mult_208_U344 ( .A(DP_N41), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n531) );
  OAI22_X1 DP_mult_208_U343 ( .A1(DP_mult_208_n531), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n532), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n325) );
  XNOR2_X1 DP_mult_208_U342 ( .A(DP_N40), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n530) );
  OAI22_X1 DP_mult_208_U341 ( .A1(DP_mult_208_n530), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n531), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n326) );
  XNOR2_X1 DP_mult_208_U340 ( .A(DP_N39), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n529) );
  OAI22_X1 DP_mult_208_U339 ( .A1(DP_mult_208_n529), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n530), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n327) );
  XNOR2_X1 DP_mult_208_U338 ( .A(DP_N38), .B(DP_mult_208_n513), .ZN(
        DP_mult_208_n528) );
  OAI22_X1 DP_mult_208_U337 ( .A1(DP_mult_208_n528), .A2(DP_mult_208_n527), 
        .B1(DP_mult_208_n529), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n328) );
  OAI22_X1 DP_mult_208_U336 ( .A1(DP_N37), .A2(DP_mult_208_n527), .B1(
        DP_mult_208_n528), .B2(DP_mult_208_n526), .ZN(DP_mult_208_n329) );
  NOR2_X1 DP_mult_208_U335 ( .A1(DP_mult_208_n525), .A2(DP_mult_208_n526), 
        .ZN(DP_coeff_ret1[0]) );
  INV_X1 DP_mult_208_U334 ( .A(DP_mult_208_n120), .ZN(DP_N73) );
  INV_X1 DP_mult_208_U333 ( .A(DP_a_int_1__1_), .ZN(DP_mult_208_n514) );
  XOR2_X2 DP_mult_208_U332 ( .A(DP_a_int_1__10_), .B(DP_mult_208_n522), .Z(
        DP_mult_208_n600) );
  XOR2_X2 DP_mult_208_U331 ( .A(DP_a_int_1__8_), .B(DP_mult_208_n520), .Z(
        DP_mult_208_n585) );
  XOR2_X2 DP_mult_208_U330 ( .A(DP_a_int_1__4_), .B(DP_mult_208_n516), .Z(
        DP_mult_208_n555) );
  XOR2_X2 DP_mult_208_U329 ( .A(DP_a_int_1__2_), .B(DP_mult_208_n514), .Z(
        DP_mult_208_n540) );
  INV_X1 DP_mult_208_U328 ( .A(DP_a_int_1__11_), .ZN(DP_mult_208_n524) );
  INV_X1 DP_mult_208_U327 ( .A(DP_a_int_1__5_), .ZN(DP_mult_208_n518) );
  INV_X1 DP_mult_208_U326 ( .A(DP_a_int_1__3_), .ZN(DP_mult_208_n516) );
  INV_X1 DP_mult_208_U325 ( .A(DP_a_int_1__9_), .ZN(DP_mult_208_n522) );
  INV_X1 DP_mult_208_U324 ( .A(DP_a_int_1__7_), .ZN(DP_mult_208_n520) );
  INV_X1 DP_mult_208_U323 ( .A(DP_mult_208_n524), .ZN(DP_mult_208_n523) );
  INV_X1 DP_mult_208_U322 ( .A(DP_mult_208_n514), .ZN(DP_mult_208_n513) );
  INV_X1 DP_mult_208_U321 ( .A(DP_mult_208_n518), .ZN(DP_mult_208_n517) );
  INV_X1 DP_mult_208_U320 ( .A(DP_mult_208_n522), .ZN(DP_mult_208_n521) );
  INV_X1 DP_mult_208_U319 ( .A(DP_mult_208_n520), .ZN(DP_mult_208_n519) );
  INV_X1 DP_mult_208_U318 ( .A(DP_mult_208_n516), .ZN(DP_mult_208_n515) );
  XOR2_X2 DP_mult_208_U317 ( .A(DP_a_int_1__6_), .B(DP_mult_208_n518), .Z(
        DP_mult_208_n570) );
  HA_X1 DP_mult_208_U107 ( .A(DP_mult_208_n316), .B(DP_mult_208_n327), .CO(
        DP_mult_208_n250), .S(DP_mult_208_n251) );
  FA_X1 DP_mult_208_U106 ( .A(DP_mult_208_n326), .B(DP_mult_208_n305), .CI(
        DP_mult_208_n315), .CO(DP_mult_208_n248), .S(DP_mult_208_n249) );
  HA_X1 DP_mult_208_U105 ( .A(DP_mult_208_n255), .B(DP_mult_208_n304), .CO(
        DP_mult_208_n246), .S(DP_mult_208_n247) );
  FA_X1 DP_mult_208_U104 ( .A(DP_mult_208_n314), .B(DP_mult_208_n325), .CI(
        DP_mult_208_n247), .CO(DP_mult_208_n244), .S(DP_mult_208_n245) );
  FA_X1 DP_mult_208_U103 ( .A(DP_mult_208_n324), .B(DP_mult_208_n293), .CI(
        DP_mult_208_n313), .CO(DP_mult_208_n242), .S(DP_mult_208_n243) );
  FA_X1 DP_mult_208_U102 ( .A(DP_mult_208_n246), .B(DP_mult_208_n303), .CI(
        DP_mult_208_n243), .CO(DP_mult_208_n240), .S(DP_mult_208_n241) );
  HA_X1 DP_mult_208_U101 ( .A(DP_mult_208_n254), .B(DP_mult_208_n292), .CO(
        DP_mult_208_n238), .S(DP_mult_208_n239) );
  FA_X1 DP_mult_208_U100 ( .A(DP_mult_208_n302), .B(DP_mult_208_n323), .CI(
        DP_mult_208_n312), .CO(DP_mult_208_n236), .S(DP_mult_208_n237) );
  FA_X1 DP_mult_208_U99 ( .A(DP_mult_208_n242), .B(DP_mult_208_n239), .CI(
        DP_mult_208_n237), .CO(DP_mult_208_n234), .S(DP_mult_208_n235) );
  FA_X1 DP_mult_208_U98 ( .A(DP_mult_208_n301), .B(DP_mult_208_n281), .CI(
        DP_mult_208_n322), .CO(DP_mult_208_n232), .S(DP_mult_208_n233) );
  FA_X1 DP_mult_208_U97 ( .A(DP_mult_208_n291), .B(DP_mult_208_n311), .CI(
        DP_mult_208_n238), .CO(DP_mult_208_n230), .S(DP_mult_208_n231) );
  FA_X1 DP_mult_208_U96 ( .A(DP_mult_208_n233), .B(DP_mult_208_n236), .CI(
        DP_mult_208_n231), .CO(DP_mult_208_n228), .S(DP_mult_208_n229) );
  HA_X1 DP_mult_208_U95 ( .A(DP_mult_208_n253), .B(DP_mult_208_n280), .CO(
        DP_mult_208_n226), .S(DP_mult_208_n227) );
  FA_X1 DP_mult_208_U94 ( .A(DP_mult_208_n290), .B(DP_mult_208_n300), .CI(
        DP_mult_208_n310), .CO(DP_mult_208_n224), .S(DP_mult_208_n225) );
  FA_X1 DP_mult_208_U93 ( .A(DP_mult_208_n227), .B(DP_mult_208_n321), .CI(
        DP_mult_208_n232), .CO(DP_mult_208_n222), .S(DP_mult_208_n223) );
  FA_X1 DP_mult_208_U92 ( .A(DP_mult_208_n225), .B(DP_mult_208_n230), .CI(
        DP_mult_208_n223), .CO(DP_mult_208_n220), .S(DP_mult_208_n221) );
  FA_X1 DP_mult_208_U91 ( .A(DP_mult_208_n289), .B(DP_mult_208_n269), .CI(
        DP_mult_208_n320), .CO(DP_mult_208_n218), .S(DP_mult_208_n219) );
  FA_X1 DP_mult_208_U90 ( .A(DP_mult_208_n279), .B(DP_mult_208_n309), .CI(
        DP_mult_208_n299), .CO(DP_mult_208_n216), .S(DP_mult_208_n217) );
  FA_X1 DP_mult_208_U89 ( .A(DP_mult_208_n224), .B(DP_mult_208_n226), .CI(
        DP_mult_208_n219), .CO(DP_mult_208_n214), .S(DP_mult_208_n215) );
  FA_X1 DP_mult_208_U88 ( .A(DP_mult_208_n222), .B(DP_mult_208_n217), .CI(
        DP_mult_208_n215), .CO(DP_mult_208_n212), .S(DP_mult_208_n213) );
  HA_X1 DP_mult_208_U87 ( .A(DP_mult_208_n252), .B(DP_mult_208_n268), .CO(
        DP_mult_208_n210), .S(DP_mult_208_n211) );
  FA_X1 DP_mult_208_U86 ( .A(DP_mult_208_n278), .B(DP_mult_208_n298), .CI(
        DP_mult_208_n319), .CO(DP_mult_208_n208), .S(DP_mult_208_n209) );
  FA_X1 DP_mult_208_U85 ( .A(DP_mult_208_n288), .B(DP_mult_208_n308), .CI(
        DP_mult_208_n211), .CO(DP_mult_208_n206), .S(DP_mult_208_n207) );
  FA_X1 DP_mult_208_U84 ( .A(DP_mult_208_n216), .B(DP_mult_208_n218), .CI(
        DP_mult_208_n209), .CO(DP_mult_208_n204), .S(DP_mult_208_n205) );
  FA_X1 DP_mult_208_U83 ( .A(DP_mult_208_n214), .B(DP_mult_208_n207), .CI(
        DP_mult_208_n205), .CO(DP_mult_208_n202), .S(DP_mult_208_n203) );
  FA_X1 DP_mult_208_U80 ( .A(DP_mult_208_n267), .B(DP_mult_208_n287), .CI(
        DP_mult_208_n318), .CO(DP_mult_208_n198), .S(DP_mult_208_n199) );
  FA_X1 DP_mult_208_U79 ( .A(DP_mult_208_n210), .B(DP_mult_208_n307), .CI(
        DP_mult_208_n201), .CO(DP_mult_208_n196), .S(DP_mult_208_n197) );
  FA_X1 DP_mult_208_U78 ( .A(DP_mult_208_n199), .B(DP_mult_208_n208), .CI(
        DP_mult_208_n206), .CO(DP_mult_208_n194), .S(DP_mult_208_n195) );
  FA_X1 DP_mult_208_U77 ( .A(DP_mult_208_n204), .B(DP_mult_208_n197), .CI(
        DP_mult_208_n195), .CO(DP_mult_208_n192), .S(DP_mult_208_n193) );
  FA_X1 DP_mult_208_U75 ( .A(DP_mult_208_n296), .B(DP_mult_208_n276), .CI(
        DP_mult_208_n191), .CO(DP_mult_208_n188), .S(DP_mult_208_n189) );
  FA_X1 DP_mult_208_U74 ( .A(DP_mult_208_n266), .B(DP_mult_208_n286), .CI(
        DP_mult_208_n200), .CO(DP_mult_208_n186), .S(DP_mult_208_n187) );
  FA_X1 DP_mult_208_U73 ( .A(DP_mult_208_n196), .B(DP_mult_208_n198), .CI(
        DP_mult_208_n189), .CO(DP_mult_208_n184), .S(DP_mult_208_n185) );
  FA_X1 DP_mult_208_U72 ( .A(DP_mult_208_n194), .B(DP_mult_208_n187), .CI(
        DP_mult_208_n185), .CO(DP_mult_208_n182), .S(DP_mult_208_n183) );
  FA_X1 DP_mult_208_U71 ( .A(DP_mult_208_n190), .B(DP_mult_208_n265), .CI(
        DP_mult_208_n306), .CO(DP_mult_208_n180), .S(DP_mult_208_n181) );
  FA_X1 DP_mult_208_U70 ( .A(DP_mult_208_n275), .B(DP_mult_208_n295), .CI(
        DP_mult_208_n285), .CO(DP_mult_208_n178), .S(DP_mult_208_n179) );
  FA_X1 DP_mult_208_U69 ( .A(DP_mult_208_n186), .B(DP_mult_208_n188), .CI(
        DP_mult_208_n179), .CO(DP_mult_208_n176), .S(DP_mult_208_n177) );
  FA_X1 DP_mult_208_U68 ( .A(DP_mult_208_n184), .B(DP_mult_208_n181), .CI(
        DP_mult_208_n177), .CO(DP_mult_208_n174), .S(DP_mult_208_n175) );
  FA_X1 DP_mult_208_U66 ( .A(DP_mult_208_n264), .B(DP_mult_208_n274), .CI(
        DP_mult_208_n173), .CO(DP_mult_208_n170), .S(DP_mult_208_n171) );
  FA_X1 DP_mult_208_U65 ( .A(DP_mult_208_n180), .B(DP_mult_208_n284), .CI(
        DP_mult_208_n178), .CO(DP_mult_208_n168), .S(DP_mult_208_n169) );
  FA_X1 DP_mult_208_U64 ( .A(DP_mult_208_n176), .B(DP_mult_208_n171), .CI(
        DP_mult_208_n169), .CO(DP_mult_208_n166), .S(DP_mult_208_n167) );
  FA_X1 DP_mult_208_U63 ( .A(DP_mult_208_n172), .B(DP_mult_208_n263), .CI(
        DP_mult_208_n294), .CO(DP_mult_208_n164), .S(DP_mult_208_n165) );
  FA_X1 DP_mult_208_U62 ( .A(DP_mult_208_n273), .B(DP_mult_208_n283), .CI(
        DP_mult_208_n170), .CO(DP_mult_208_n162), .S(DP_mult_208_n163) );
  FA_X1 DP_mult_208_U61 ( .A(DP_mult_208_n168), .B(DP_mult_208_n165), .CI(
        DP_mult_208_n163), .CO(DP_mult_208_n160), .S(DP_mult_208_n161) );
  FA_X1 DP_mult_208_U59 ( .A(DP_mult_208_n262), .B(DP_mult_208_n272), .CI(
        DP_mult_208_n159), .CO(DP_mult_208_n156), .S(DP_mult_208_n157) );
  FA_X1 DP_mult_208_U58 ( .A(DP_mult_208_n157), .B(DP_mult_208_n164), .CI(
        DP_mult_208_n162), .CO(DP_mult_208_n154), .S(DP_mult_208_n155) );
  FA_X1 DP_mult_208_U57 ( .A(DP_mult_208_n261), .B(DP_mult_208_n158), .CI(
        DP_mult_208_n282), .CO(DP_mult_208_n152), .S(DP_mult_208_n153) );
  FA_X1 DP_mult_208_U56 ( .A(DP_mult_208_n156), .B(DP_mult_208_n271), .CI(
        DP_mult_208_n153), .CO(DP_mult_208_n150), .S(DP_mult_208_n151) );
  FA_X1 DP_mult_208_U54 ( .A(DP_mult_208_n149), .B(DP_mult_208_n260), .CI(
        DP_mult_208_n152), .CO(DP_mult_208_n146), .S(DP_mult_208_n147) );
  FA_X1 DP_mult_208_U53 ( .A(DP_mult_208_n259), .B(DP_mult_208_n148), .CI(
        DP_mult_208_n270), .CO(DP_mult_208_n144), .S(DP_mult_208_n145) );
  HA_X1 DP_mult_208_U51 ( .A(DP_mult_208_n329), .B(DP_mult_208_n257), .CO(
        DP_mult_208_n141), .S(DP_N51) );
  FA_X1 DP_mult_208_U50 ( .A(DP_mult_208_n328), .B(DP_mult_208_n317), .CI(
        DP_mult_208_n141), .CO(DP_mult_208_n140), .S(DP_N52) );
  FA_X1 DP_mult_208_U49 ( .A(DP_mult_208_n251), .B(DP_mult_208_n256), .CI(
        DP_mult_208_n140), .CO(DP_mult_208_n139), .S(DP_N53) );
  FA_X1 DP_mult_208_U48 ( .A(DP_mult_208_n249), .B(DP_mult_208_n250), .CI(
        DP_mult_208_n139), .CO(DP_mult_208_n138), .S(DP_N54) );
  FA_X1 DP_mult_208_U47 ( .A(DP_mult_208_n245), .B(DP_mult_208_n248), .CI(
        DP_mult_208_n138), .CO(DP_mult_208_n137), .S(DP_N55) );
  FA_X1 DP_mult_208_U46 ( .A(DP_mult_208_n241), .B(DP_mult_208_n244), .CI(
        DP_mult_208_n137), .CO(DP_mult_208_n136), .S(DP_N56) );
  FA_X1 DP_mult_208_U45 ( .A(DP_mult_208_n235), .B(DP_mult_208_n240), .CI(
        DP_mult_208_n136), .CO(DP_mult_208_n135), .S(DP_N57) );
  FA_X1 DP_mult_208_U44 ( .A(DP_mult_208_n229), .B(DP_mult_208_n234), .CI(
        DP_mult_208_n135), .CO(DP_mult_208_n134), .S(DP_N58) );
  FA_X1 DP_mult_208_U43 ( .A(DP_mult_208_n221), .B(DP_mult_208_n228), .CI(
        DP_mult_208_n134), .CO(DP_mult_208_n133), .S(DP_N59) );
  FA_X1 DP_mult_208_U42 ( .A(DP_mult_208_n213), .B(DP_mult_208_n220), .CI(
        DP_mult_208_n133), .CO(DP_mult_208_n132), .S(DP_N60) );
  FA_X1 DP_mult_208_U41 ( .A(DP_mult_208_n203), .B(DP_mult_208_n212), .CI(
        DP_mult_208_n132), .CO(DP_mult_208_n131), .S(DP_N61) );
  FA_X1 DP_mult_208_U40 ( .A(DP_mult_208_n193), .B(DP_mult_208_n202), .CI(
        DP_mult_208_n131), .CO(DP_mult_208_n130), .S(DP_N62) );
  FA_X1 DP_mult_208_U39 ( .A(DP_mult_208_n183), .B(DP_mult_208_n192), .CI(
        DP_mult_208_n130), .CO(DP_mult_208_n129), .S(DP_N63) );
  FA_X1 DP_mult_208_U38 ( .A(DP_mult_208_n175), .B(DP_mult_208_n182), .CI(
        DP_mult_208_n129), .CO(DP_mult_208_n128), .S(DP_N64) );
  FA_X1 DP_mult_208_U37 ( .A(DP_mult_208_n167), .B(DP_mult_208_n174), .CI(
        DP_mult_208_n128), .CO(DP_mult_208_n127), .S(DP_N65) );
  FA_X1 DP_mult_208_U36 ( .A(DP_mult_208_n161), .B(DP_mult_208_n166), .CI(
        DP_mult_208_n127), .CO(DP_mult_208_n126), .S(DP_N66) );
  FA_X1 DP_mult_208_U30 ( .A(DP_mult_208_n160), .B(DP_mult_208_n155), .CI(
        DP_mult_208_n126), .CO(DP_mult_208_n125), .S(DP_N67) );
  FA_X1 DP_mult_208_U20 ( .A(DP_mult_208_n151), .B(DP_mult_208_n154), .CI(
        DP_mult_208_n125), .CO(DP_mult_208_n124), .S(DP_N68) );
  FA_X1 DP_mult_208_U10 ( .A(DP_mult_208_n147), .B(DP_mult_208_n150), .CI(
        DP_mult_208_n124), .CO(DP_mult_208_n123), .S(DP_N69) );
  FA_X1 DP_mult_208_U9 ( .A(DP_mult_208_n146), .B(DP_mult_208_n145), .CI(
        DP_mult_208_n123), .CO(DP_mult_208_n122), .S(DP_N70) );
  FA_X1 DP_mult_208_U8 ( .A(DP_mult_208_n144), .B(DP_mult_208_n143), .CI(
        DP_mult_208_n122), .CO(DP_mult_208_n121), .S(DP_N71) );
  FA_X1 DP_mult_208_U7 ( .A(DP_mult_208_n258), .B(DP_mult_208_n142), .CI(
        DP_mult_208_n121), .CO(DP_mult_208_n120), .S(DP_N72) );
  INV_X1 DP_sub_208_U69 ( .A(DP_N60), .ZN(DP_sub_208_B_not_10_) );
  INV_X1 DP_sub_208_U68 ( .A(DP_N61), .ZN(DP_sub_208_B_not_11_) );
  INV_X1 DP_sub_208_U67 ( .A(DP_N62), .ZN(DP_sub_208_B_not_12_) );
  INV_X1 DP_sub_208_U66 ( .A(DP_N63), .ZN(DP_sub_208_B_not_13_) );
  INV_X1 DP_sub_208_U65 ( .A(DP_N64), .ZN(DP_sub_208_B_not_14_) );
  INV_X1 DP_sub_208_U64 ( .A(DP_N65), .ZN(DP_sub_208_B_not_15_) );
  INV_X1 DP_sub_208_U63 ( .A(DP_N66), .ZN(DP_sub_208_B_not_16_) );
  INV_X1 DP_sub_208_U62 ( .A(DP_N67), .ZN(DP_sub_208_B_not_17_) );
  INV_X1 DP_sub_208_U61 ( .A(DP_N68), .ZN(DP_sub_208_B_not_18_) );
  INV_X1 DP_sub_208_U60 ( .A(DP_N69), .ZN(DP_sub_208_B_not_19_) );
  INV_X1 DP_sub_208_U59 ( .A(DP_N51), .ZN(DP_sub_208_B_not_1_) );
  INV_X1 DP_sub_208_U58 ( .A(DP_N70), .ZN(DP_sub_208_B_not_20_) );
  INV_X1 DP_sub_208_U57 ( .A(DP_N71), .ZN(DP_sub_208_B_not_21_) );
  INV_X1 DP_sub_208_U56 ( .A(DP_N72), .ZN(DP_sub_208_B_not_22_) );
  INV_X1 DP_sub_208_U55 ( .A(DP_N73), .ZN(DP_sub_208_B_not_23_) );
  INV_X1 DP_sub_208_U54 ( .A(DP_N52), .ZN(DP_sub_208_B_not_2_) );
  INV_X1 DP_sub_208_U53 ( .A(DP_N53), .ZN(DP_sub_208_B_not_3_) );
  INV_X1 DP_sub_208_U52 ( .A(DP_N54), .ZN(DP_sub_208_B_not_4_) );
  INV_X1 DP_sub_208_U51 ( .A(DP_N55), .ZN(DP_sub_208_B_not_5_) );
  INV_X1 DP_sub_208_U50 ( .A(DP_N56), .ZN(DP_sub_208_B_not_6_) );
  INV_X1 DP_sub_208_U49 ( .A(DP_N57), .ZN(DP_sub_208_B_not_7_) );
  INV_X1 DP_sub_208_U48 ( .A(DP_N58), .ZN(DP_sub_208_B_not_8_) );
  INV_X1 DP_sub_208_U47 ( .A(DP_N59), .ZN(DP_sub_208_B_not_9_) );
  INV_X1 DP_sub_208_U46 ( .A(DP_coeff_ret1[0]), .ZN(DP_sub_208_carry_1_) );
  XOR2_X1 DP_sub_208_U45 ( .A(DP_sub_208_B_not_1_), .B(DP_sub_208_carry_1_), 
        .Z(DP_coeff_ret1[1]) );
  AND2_X1 DP_sub_208_U44 ( .A1(DP_sub_208_carry_1_), .A2(DP_sub_208_B_not_1_), 
        .ZN(DP_sub_208_carry_2_) );
  AND2_X1 DP_sub_208_U43 ( .A1(DP_sub_208_carry_2_), .A2(DP_sub_208_B_not_2_), 
        .ZN(DP_sub_208_carry_3_) );
  XOR2_X1 DP_sub_208_U42 ( .A(DP_sub_208_B_not_3_), .B(DP_sub_208_carry_3_), 
        .Z(DP_coeff_ret1[3]) );
  AND2_X1 DP_sub_208_U41 ( .A1(DP_sub_208_carry_3_), .A2(DP_sub_208_B_not_3_), 
        .ZN(DP_sub_208_carry_4_) );
  XOR2_X1 DP_sub_208_U40 ( .A(DP_sub_208_B_not_4_), .B(DP_sub_208_carry_4_), 
        .Z(DP_coeff_ret1[4]) );
  AND2_X1 DP_sub_208_U39 ( .A1(DP_sub_208_carry_4_), .A2(DP_sub_208_B_not_4_), 
        .ZN(DP_sub_208_carry_5_) );
  XOR2_X1 DP_sub_208_U38 ( .A(DP_sub_208_B_not_5_), .B(DP_sub_208_carry_5_), 
        .Z(DP_coeff_ret1[5]) );
  AND2_X1 DP_sub_208_U37 ( .A1(DP_sub_208_carry_5_), .A2(DP_sub_208_B_not_5_), 
        .ZN(DP_sub_208_carry_6_) );
  XOR2_X1 DP_sub_208_U36 ( .A(DP_sub_208_B_not_6_), .B(DP_sub_208_carry_6_), 
        .Z(DP_coeff_ret1[6]) );
  AND2_X1 DP_sub_208_U35 ( .A1(DP_sub_208_carry_6_), .A2(DP_sub_208_B_not_6_), 
        .ZN(DP_sub_208_carry_7_) );
  XOR2_X1 DP_sub_208_U34 ( .A(DP_sub_208_B_not_7_), .B(DP_sub_208_carry_7_), 
        .Z(DP_coeff_ret1[7]) );
  AND2_X1 DP_sub_208_U33 ( .A1(DP_sub_208_carry_7_), .A2(DP_sub_208_B_not_7_), 
        .ZN(DP_sub_208_carry_8_) );
  XOR2_X1 DP_sub_208_U32 ( .A(DP_sub_208_B_not_8_), .B(DP_sub_208_carry_8_), 
        .Z(DP_coeff_ret1[8]) );
  AND2_X1 DP_sub_208_U31 ( .A1(DP_sub_208_carry_8_), .A2(DP_sub_208_B_not_8_), 
        .ZN(DP_sub_208_carry_9_) );
  XOR2_X1 DP_sub_208_U30 ( .A(DP_sub_208_B_not_9_), .B(DP_sub_208_carry_9_), 
        .Z(DP_coeff_ret1[9]) );
  AND2_X1 DP_sub_208_U29 ( .A1(DP_sub_208_carry_9_), .A2(DP_sub_208_B_not_9_), 
        .ZN(DP_sub_208_carry_10_) );
  XOR2_X1 DP_sub_208_U28 ( .A(DP_sub_208_B_not_10_), .B(DP_sub_208_carry_10_), 
        .Z(DP_coeff_ret1[10]) );
  AND2_X1 DP_sub_208_U27 ( .A1(DP_sub_208_carry_10_), .A2(DP_sub_208_B_not_10_), .ZN(DP_sub_208_carry_11_) );
  XOR2_X1 DP_sub_208_U26 ( .A(DP_sub_208_B_not_11_), .B(DP_sub_208_carry_11_), 
        .Z(DP_coeff_ret1[11]) );
  AND2_X1 DP_sub_208_U25 ( .A1(DP_sub_208_carry_11_), .A2(DP_sub_208_B_not_11_), .ZN(DP_sub_208_carry_12_) );
  XOR2_X1 DP_sub_208_U24 ( .A(DP_sub_208_B_not_12_), .B(DP_sub_208_carry_12_), 
        .Z(DP_coeff_ret1[12]) );
  AND2_X1 DP_sub_208_U23 ( .A1(DP_sub_208_carry_12_), .A2(DP_sub_208_B_not_12_), .ZN(DP_sub_208_carry_13_) );
  XOR2_X1 DP_sub_208_U22 ( .A(DP_sub_208_B_not_13_), .B(DP_sub_208_carry_13_), 
        .Z(DP_coeff_ret1[13]) );
  AND2_X1 DP_sub_208_U21 ( .A1(DP_sub_208_carry_13_), .A2(DP_sub_208_B_not_13_), .ZN(DP_sub_208_carry_14_) );
  XOR2_X1 DP_sub_208_U20 ( .A(DP_sub_208_B_not_14_), .B(DP_sub_208_carry_14_), 
        .Z(DP_coeff_ret1[14]) );
  AND2_X1 DP_sub_208_U19 ( .A1(DP_sub_208_carry_14_), .A2(DP_sub_208_B_not_14_), .ZN(DP_sub_208_carry_15_) );
  XOR2_X1 DP_sub_208_U18 ( .A(DP_sub_208_B_not_15_), .B(DP_sub_208_carry_15_), 
        .Z(DP_coeff_ret1[15]) );
  AND2_X1 DP_sub_208_U17 ( .A1(DP_sub_208_carry_15_), .A2(DP_sub_208_B_not_15_), .ZN(DP_sub_208_carry_16_) );
  XOR2_X1 DP_sub_208_U16 ( .A(DP_sub_208_B_not_16_), .B(DP_sub_208_carry_16_), 
        .Z(DP_coeff_ret1[16]) );
  AND2_X1 DP_sub_208_U15 ( .A1(DP_sub_208_carry_16_), .A2(DP_sub_208_B_not_16_), .ZN(DP_sub_208_carry_17_) );
  XOR2_X1 DP_sub_208_U14 ( .A(DP_sub_208_B_not_17_), .B(DP_sub_208_carry_17_), 
        .Z(DP_coeff_ret1[17]) );
  AND2_X1 DP_sub_208_U13 ( .A1(DP_sub_208_carry_17_), .A2(DP_sub_208_B_not_17_), .ZN(DP_sub_208_carry_18_) );
  XOR2_X1 DP_sub_208_U12 ( .A(DP_sub_208_B_not_18_), .B(DP_sub_208_carry_18_), 
        .Z(DP_coeff_ret1[18]) );
  AND2_X1 DP_sub_208_U11 ( .A1(DP_sub_208_carry_18_), .A2(DP_sub_208_B_not_18_), .ZN(DP_sub_208_carry_19_) );
  XOR2_X1 DP_sub_208_U10 ( .A(DP_sub_208_B_not_19_), .B(DP_sub_208_carry_19_), 
        .Z(DP_coeff_ret1[19]) );
  AND2_X1 DP_sub_208_U9 ( .A1(DP_sub_208_carry_19_), .A2(DP_sub_208_B_not_19_), 
        .ZN(DP_sub_208_carry_20_) );
  XOR2_X1 DP_sub_208_U8 ( .A(DP_sub_208_B_not_20_), .B(DP_sub_208_carry_20_), 
        .Z(DP_coeff_ret1[20]) );
  AND2_X1 DP_sub_208_U7 ( .A1(DP_sub_208_carry_20_), .A2(DP_sub_208_B_not_20_), 
        .ZN(DP_sub_208_carry_21_) );
  XOR2_X1 DP_sub_208_U6 ( .A(DP_sub_208_B_not_21_), .B(DP_sub_208_carry_21_), 
        .Z(DP_coeff_ret1[21]) );
  AND2_X1 DP_sub_208_U5 ( .A1(DP_sub_208_carry_21_), .A2(DP_sub_208_B_not_21_), 
        .ZN(DP_sub_208_carry_22_) );
  XOR2_X1 DP_sub_208_U4 ( .A(DP_sub_208_B_not_22_), .B(DP_sub_208_carry_22_), 
        .Z(DP_coeff_ret1[22]) );
  AND2_X1 DP_sub_208_U3 ( .A1(DP_sub_208_carry_22_), .A2(DP_sub_208_B_not_22_), 
        .ZN(DP_sub_208_carry_23_) );
  XOR2_X1 DP_sub_208_U2 ( .A(DP_sub_208_B_not_23_), .B(DP_sub_208_carry_23_), 
        .Z(DP_coeff_ret1[23]) );
  XOR2_X2 DP_sub_208_U1 ( .A(DP_sub_208_B_not_2_), .B(DP_sub_208_carry_2_), 
        .Z(DP_coeff_ret1[2]) );
  XNOR2_X1 DP_mult_209_U520 ( .A(DP_b_int_0__10_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n612) );
  XNOR2_X1 DP_mult_209_U519 ( .A(DP_mult_209_n524), .B(DP_a_int_1__10_), .ZN(
        DP_mult_209_n626) );
  NAND2_X1 DP_mult_209_U518 ( .A1(DP_mult_209_n600), .A2(DP_mult_209_n626), 
        .ZN(DP_mult_209_n602) );
  XNOR2_X1 DP_mult_209_U517 ( .A(DP_b_int_0__11_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n614) );
  OAI22_X1 DP_mult_209_U516 ( .A1(DP_mult_209_n612), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n614), .ZN(DP_mult_209_n142) );
  INV_X1 DP_mult_209_U515 ( .A(DP_mult_209_n142), .ZN(DP_mult_209_n143) );
  XNOR2_X1 DP_mult_209_U514 ( .A(DP_b_int_0__10_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n597) );
  XNOR2_X1 DP_mult_209_U513 ( .A(DP_mult_209_n522), .B(DP_a_int_1__8_), .ZN(
        DP_mult_209_n625) );
  NAND2_X1 DP_mult_209_U512 ( .A1(DP_mult_209_n585), .A2(DP_mult_209_n625), 
        .ZN(DP_mult_209_n587) );
  XNOR2_X1 DP_mult_209_U511 ( .A(DP_b_int_0__11_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n599) );
  OAI22_X1 DP_mult_209_U510 ( .A1(DP_mult_209_n597), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n599), .ZN(DP_mult_209_n148) );
  INV_X1 DP_mult_209_U509 ( .A(DP_mult_209_n148), .ZN(DP_mult_209_n149) );
  XNOR2_X1 DP_mult_209_U508 ( .A(DP_b_int_0__10_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n582) );
  XNOR2_X1 DP_mult_209_U507 ( .A(DP_mult_209_n520), .B(DP_a_int_1__6_), .ZN(
        DP_mult_209_n624) );
  NAND2_X1 DP_mult_209_U506 ( .A1(DP_mult_209_n570), .A2(DP_mult_209_n624), 
        .ZN(DP_mult_209_n572) );
  XNOR2_X1 DP_mult_209_U505 ( .A(DP_b_int_0__11_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n584) );
  OAI22_X1 DP_mult_209_U504 ( .A1(DP_mult_209_n582), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n584), .ZN(DP_mult_209_n158) );
  INV_X1 DP_mult_209_U503 ( .A(DP_mult_209_n158), .ZN(DP_mult_209_n159) );
  XNOR2_X1 DP_mult_209_U502 ( .A(DP_b_int_0__10_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n567) );
  XNOR2_X1 DP_mult_209_U501 ( .A(DP_mult_209_n518), .B(DP_a_int_1__4_), .ZN(
        DP_mult_209_n623) );
  NAND2_X1 DP_mult_209_U500 ( .A1(DP_mult_209_n555), .A2(DP_mult_209_n623), 
        .ZN(DP_mult_209_n557) );
  XNOR2_X1 DP_mult_209_U499 ( .A(DP_b_int_0__11_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n569) );
  OAI22_X1 DP_mult_209_U498 ( .A1(DP_mult_209_n567), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n569), .ZN(DP_mult_209_n172) );
  INV_X1 DP_mult_209_U497 ( .A(DP_mult_209_n172), .ZN(DP_mult_209_n173) );
  XNOR2_X1 DP_mult_209_U496 ( .A(DP_b_int_0__10_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n552) );
  XNOR2_X1 DP_mult_209_U495 ( .A(DP_mult_209_n516), .B(DP_a_int_1__2_), .ZN(
        DP_mult_209_n622) );
  NAND2_X1 DP_mult_209_U494 ( .A1(DP_mult_209_n540), .A2(DP_mult_209_n622), 
        .ZN(DP_mult_209_n542) );
  XNOR2_X1 DP_mult_209_U493 ( .A(DP_b_int_0__11_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n554) );
  OAI22_X1 DP_mult_209_U492 ( .A1(DP_mult_209_n552), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n554), .ZN(DP_mult_209_n190) );
  INV_X1 DP_mult_209_U491 ( .A(DP_mult_209_n190), .ZN(DP_mult_209_n191) );
  XNOR2_X1 DP_mult_209_U490 ( .A(DP_b_int_0__3_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n590) );
  XNOR2_X1 DP_mult_209_U489 ( .A(DP_b_int_0__4_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n591) );
  OAI22_X1 DP_mult_209_U488 ( .A1(DP_mult_209_n590), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n591), .ZN(DP_mult_209_n620) );
  XNOR2_X1 DP_mult_209_U487 ( .A(DP_b_int_0__7_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n564) );
  XNOR2_X1 DP_mult_209_U486 ( .A(DP_b_int_0__8_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n565) );
  OAI22_X1 DP_mult_209_U485 ( .A1(DP_mult_209_n564), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n565), .ZN(DP_mult_209_n621) );
  OR2_X1 DP_mult_209_U484 ( .A1(DP_mult_209_n620), .A2(DP_mult_209_n621), .ZN(
        DP_mult_209_n200) );
  XNOR2_X1 DP_mult_209_U483 ( .A(DP_mult_209_n620), .B(DP_mult_209_n621), .ZN(
        DP_mult_209_n201) );
  OR3_X1 DP_mult_209_U482 ( .A1(DP_mult_209_n600), .A2(DP_b_int_0__0_), .A3(
        DP_mult_209_n524), .ZN(DP_mult_209_n619) );
  OAI21_X1 DP_mult_209_U481 ( .B1(DP_mult_209_n524), .B2(DP_mult_209_n602), 
        .A(DP_mult_209_n619), .ZN(DP_mult_209_n252) );
  OR3_X1 DP_mult_209_U480 ( .A1(DP_mult_209_n585), .A2(DP_b_int_0__0_), .A3(
        DP_mult_209_n522), .ZN(DP_mult_209_n618) );
  OAI21_X1 DP_mult_209_U479 ( .B1(DP_mult_209_n522), .B2(DP_mult_209_n587), 
        .A(DP_mult_209_n618), .ZN(DP_mult_209_n253) );
  OR3_X1 DP_mult_209_U478 ( .A1(DP_mult_209_n570), .A2(DP_b_int_0__0_), .A3(
        DP_mult_209_n520), .ZN(DP_mult_209_n617) );
  OAI21_X1 DP_mult_209_U477 ( .B1(DP_mult_209_n520), .B2(DP_mult_209_n572), 
        .A(DP_mult_209_n617), .ZN(DP_mult_209_n254) );
  OR3_X1 DP_mult_209_U476 ( .A1(DP_mult_209_n555), .A2(DP_b_int_0__0_), .A3(
        DP_mult_209_n518), .ZN(DP_mult_209_n616) );
  OAI21_X1 DP_mult_209_U475 ( .B1(DP_mult_209_n518), .B2(DP_mult_209_n557), 
        .A(DP_mult_209_n616), .ZN(DP_mult_209_n255) );
  OR3_X1 DP_mult_209_U474 ( .A1(DP_mult_209_n540), .A2(DP_b_int_0__0_), .A3(
        DP_mult_209_n516), .ZN(DP_mult_209_n615) );
  OAI21_X1 DP_mult_209_U473 ( .B1(DP_mult_209_n516), .B2(DP_mult_209_n542), 
        .A(DP_mult_209_n615), .ZN(DP_mult_209_n256) );
  INV_X1 DP_mult_209_U472 ( .A(DP_coeff_ret0[1]), .ZN(DP_mult_209_n526) );
  NAND2_X1 DP_mult_209_U471 ( .A1(DP_mult_209_n513), .A2(DP_mult_209_n526), 
        .ZN(DP_mult_209_n527) );
  OAI21_X1 DP_mult_209_U470 ( .B1(DP_b_int_0__0_), .B2(DP_mult_209_n514), .A(
        DP_mult_209_n527), .ZN(DP_mult_209_n257) );
  AOI21_X1 DP_mult_209_U469 ( .B1(DP_mult_209_n602), .B2(DP_mult_209_n600), 
        .A(DP_mult_209_n614), .ZN(DP_mult_209_n613) );
  INV_X1 DP_mult_209_U468 ( .A(DP_mult_209_n613), .ZN(DP_mult_209_n258) );
  XNOR2_X1 DP_mult_209_U467 ( .A(DP_b_int_0__9_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n611) );
  OAI22_X1 DP_mult_209_U466 ( .A1(DP_mult_209_n611), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n612), .ZN(DP_mult_209_n259) );
  XNOR2_X1 DP_mult_209_U465 ( .A(DP_b_int_0__8_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n610) );
  OAI22_X1 DP_mult_209_U464 ( .A1(DP_mult_209_n610), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n611), .ZN(DP_mult_209_n260) );
  XNOR2_X1 DP_mult_209_U463 ( .A(DP_b_int_0__7_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n609) );
  OAI22_X1 DP_mult_209_U462 ( .A1(DP_mult_209_n609), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n610), .ZN(DP_mult_209_n261) );
  XNOR2_X1 DP_mult_209_U461 ( .A(DP_b_int_0__6_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n608) );
  OAI22_X1 DP_mult_209_U460 ( .A1(DP_mult_209_n608), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n609), .ZN(DP_mult_209_n262) );
  XNOR2_X1 DP_mult_209_U459 ( .A(DP_b_int_0__5_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n607) );
  OAI22_X1 DP_mult_209_U458 ( .A1(DP_mult_209_n607), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n608), .ZN(DP_mult_209_n263) );
  XNOR2_X1 DP_mult_209_U457 ( .A(DP_b_int_0__4_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n606) );
  OAI22_X1 DP_mult_209_U456 ( .A1(DP_mult_209_n606), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n607), .ZN(DP_mult_209_n264) );
  XNOR2_X1 DP_mult_209_U455 ( .A(DP_b_int_0__3_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n605) );
  OAI22_X1 DP_mult_209_U454 ( .A1(DP_mult_209_n605), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n606), .ZN(DP_mult_209_n265) );
  XNOR2_X1 DP_mult_209_U453 ( .A(DP_b_int_0__2_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n604) );
  OAI22_X1 DP_mult_209_U452 ( .A1(DP_mult_209_n604), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n605), .ZN(DP_mult_209_n266) );
  XNOR2_X1 DP_mult_209_U451 ( .A(DP_b_int_0__1_), .B(DP_mult_209_n523), .ZN(
        DP_mult_209_n603) );
  OAI22_X1 DP_mult_209_U450 ( .A1(DP_mult_209_n603), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n604), .ZN(DP_mult_209_n267) );
  XNOR2_X1 DP_mult_209_U449 ( .A(DP_mult_209_n523), .B(DP_b_int_0__0_), .ZN(
        DP_mult_209_n601) );
  OAI22_X1 DP_mult_209_U448 ( .A1(DP_mult_209_n601), .A2(DP_mult_209_n602), 
        .B1(DP_mult_209_n600), .B2(DP_mult_209_n603), .ZN(DP_mult_209_n268) );
  INV_X1 DP_mult_209_U447 ( .A(DP_b_int_0__0_), .ZN(DP_mult_209_n525) );
  NOR2_X1 DP_mult_209_U446 ( .A1(DP_mult_209_n525), .A2(DP_mult_209_n600), 
        .ZN(DP_mult_209_n269) );
  AOI21_X1 DP_mult_209_U445 ( .B1(DP_mult_209_n587), .B2(DP_mult_209_n585), 
        .A(DP_mult_209_n599), .ZN(DP_mult_209_n598) );
  INV_X1 DP_mult_209_U444 ( .A(DP_mult_209_n598), .ZN(DP_mult_209_n270) );
  XNOR2_X1 DP_mult_209_U443 ( .A(DP_b_int_0__9_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n596) );
  OAI22_X1 DP_mult_209_U442 ( .A1(DP_mult_209_n596), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n597), .ZN(DP_mult_209_n271) );
  XNOR2_X1 DP_mult_209_U441 ( .A(DP_b_int_0__8_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n595) );
  OAI22_X1 DP_mult_209_U440 ( .A1(DP_mult_209_n595), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n596), .ZN(DP_mult_209_n272) );
  XNOR2_X1 DP_mult_209_U439 ( .A(DP_b_int_0__7_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n594) );
  OAI22_X1 DP_mult_209_U438 ( .A1(DP_mult_209_n594), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n595), .ZN(DP_mult_209_n273) );
  XNOR2_X1 DP_mult_209_U437 ( .A(DP_b_int_0__6_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n593) );
  OAI22_X1 DP_mult_209_U436 ( .A1(DP_mult_209_n593), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n594), .ZN(DP_mult_209_n274) );
  XNOR2_X1 DP_mult_209_U435 ( .A(DP_b_int_0__5_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n592) );
  OAI22_X1 DP_mult_209_U434 ( .A1(DP_mult_209_n592), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n593), .ZN(DP_mult_209_n275) );
  OAI22_X1 DP_mult_209_U433 ( .A1(DP_mult_209_n591), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n592), .ZN(DP_mult_209_n276) );
  XNOR2_X1 DP_mult_209_U432 ( .A(DP_b_int_0__2_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n589) );
  OAI22_X1 DP_mult_209_U431 ( .A1(DP_mult_209_n589), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n590), .ZN(DP_mult_209_n278) );
  XNOR2_X1 DP_mult_209_U430 ( .A(DP_b_int_0__1_), .B(DP_mult_209_n521), .ZN(
        DP_mult_209_n588) );
  OAI22_X1 DP_mult_209_U429 ( .A1(DP_mult_209_n588), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n589), .ZN(DP_mult_209_n279) );
  XNOR2_X1 DP_mult_209_U428 ( .A(DP_mult_209_n521), .B(DP_b_int_0__0_), .ZN(
        DP_mult_209_n586) );
  OAI22_X1 DP_mult_209_U427 ( .A1(DP_mult_209_n586), .A2(DP_mult_209_n587), 
        .B1(DP_mult_209_n585), .B2(DP_mult_209_n588), .ZN(DP_mult_209_n280) );
  NOR2_X1 DP_mult_209_U426 ( .A1(DP_mult_209_n525), .A2(DP_mult_209_n585), 
        .ZN(DP_mult_209_n281) );
  AOI21_X1 DP_mult_209_U425 ( .B1(DP_mult_209_n572), .B2(DP_mult_209_n570), 
        .A(DP_mult_209_n584), .ZN(DP_mult_209_n583) );
  INV_X1 DP_mult_209_U424 ( .A(DP_mult_209_n583), .ZN(DP_mult_209_n282) );
  XNOR2_X1 DP_mult_209_U423 ( .A(DP_b_int_0__9_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n581) );
  OAI22_X1 DP_mult_209_U422 ( .A1(DP_mult_209_n581), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n582), .ZN(DP_mult_209_n283) );
  XNOR2_X1 DP_mult_209_U421 ( .A(DP_b_int_0__8_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n580) );
  OAI22_X1 DP_mult_209_U420 ( .A1(DP_mult_209_n580), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n581), .ZN(DP_mult_209_n284) );
  XNOR2_X1 DP_mult_209_U419 ( .A(DP_b_int_0__7_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n579) );
  OAI22_X1 DP_mult_209_U418 ( .A1(DP_mult_209_n579), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n580), .ZN(DP_mult_209_n285) );
  XNOR2_X1 DP_mult_209_U417 ( .A(DP_b_int_0__6_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n578) );
  OAI22_X1 DP_mult_209_U416 ( .A1(DP_mult_209_n578), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n579), .ZN(DP_mult_209_n286) );
  XNOR2_X1 DP_mult_209_U415 ( .A(DP_b_int_0__5_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n577) );
  OAI22_X1 DP_mult_209_U414 ( .A1(DP_mult_209_n577), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n578), .ZN(DP_mult_209_n287) );
  XNOR2_X1 DP_mult_209_U413 ( .A(DP_b_int_0__4_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n576) );
  OAI22_X1 DP_mult_209_U412 ( .A1(DP_mult_209_n576), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n577), .ZN(DP_mult_209_n288) );
  XNOR2_X1 DP_mult_209_U411 ( .A(DP_b_int_0__3_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n575) );
  OAI22_X1 DP_mult_209_U410 ( .A1(DP_mult_209_n575), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n576), .ZN(DP_mult_209_n289) );
  XNOR2_X1 DP_mult_209_U409 ( .A(DP_b_int_0__2_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n574) );
  OAI22_X1 DP_mult_209_U408 ( .A1(DP_mult_209_n574), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n575), .ZN(DP_mult_209_n290) );
  XNOR2_X1 DP_mult_209_U407 ( .A(DP_b_int_0__1_), .B(DP_mult_209_n519), .ZN(
        DP_mult_209_n573) );
  OAI22_X1 DP_mult_209_U406 ( .A1(DP_mult_209_n573), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n574), .ZN(DP_mult_209_n291) );
  XNOR2_X1 DP_mult_209_U405 ( .A(DP_mult_209_n519), .B(DP_b_int_0__0_), .ZN(
        DP_mult_209_n571) );
  OAI22_X1 DP_mult_209_U404 ( .A1(DP_mult_209_n571), .A2(DP_mult_209_n572), 
        .B1(DP_mult_209_n570), .B2(DP_mult_209_n573), .ZN(DP_mult_209_n292) );
  NOR2_X1 DP_mult_209_U403 ( .A1(DP_mult_209_n525), .A2(DP_mult_209_n570), 
        .ZN(DP_mult_209_n293) );
  AOI21_X1 DP_mult_209_U402 ( .B1(DP_mult_209_n557), .B2(DP_mult_209_n555), 
        .A(DP_mult_209_n569), .ZN(DP_mult_209_n568) );
  INV_X1 DP_mult_209_U401 ( .A(DP_mult_209_n568), .ZN(DP_mult_209_n294) );
  XNOR2_X1 DP_mult_209_U400 ( .A(DP_b_int_0__9_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n566) );
  OAI22_X1 DP_mult_209_U399 ( .A1(DP_mult_209_n566), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n567), .ZN(DP_mult_209_n295) );
  OAI22_X1 DP_mult_209_U398 ( .A1(DP_mult_209_n565), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n566), .ZN(DP_mult_209_n296) );
  XNOR2_X1 DP_mult_209_U397 ( .A(DP_b_int_0__6_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n563) );
  OAI22_X1 DP_mult_209_U396 ( .A1(DP_mult_209_n563), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n564), .ZN(DP_mult_209_n298) );
  XNOR2_X1 DP_mult_209_U395 ( .A(DP_b_int_0__5_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n562) );
  OAI22_X1 DP_mult_209_U394 ( .A1(DP_mult_209_n562), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n563), .ZN(DP_mult_209_n299) );
  XNOR2_X1 DP_mult_209_U393 ( .A(DP_b_int_0__4_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n561) );
  OAI22_X1 DP_mult_209_U392 ( .A1(DP_mult_209_n561), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n562), .ZN(DP_mult_209_n300) );
  XNOR2_X1 DP_mult_209_U391 ( .A(DP_b_int_0__3_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n560) );
  OAI22_X1 DP_mult_209_U390 ( .A1(DP_mult_209_n560), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n561), .ZN(DP_mult_209_n301) );
  XNOR2_X1 DP_mult_209_U389 ( .A(DP_b_int_0__2_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n559) );
  OAI22_X1 DP_mult_209_U388 ( .A1(DP_mult_209_n559), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n560), .ZN(DP_mult_209_n302) );
  XNOR2_X1 DP_mult_209_U387 ( .A(DP_b_int_0__1_), .B(DP_mult_209_n517), .ZN(
        DP_mult_209_n558) );
  OAI22_X1 DP_mult_209_U386 ( .A1(DP_mult_209_n558), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n559), .ZN(DP_mult_209_n303) );
  XNOR2_X1 DP_mult_209_U385 ( .A(DP_mult_209_n517), .B(DP_b_int_0__0_), .ZN(
        DP_mult_209_n556) );
  OAI22_X1 DP_mult_209_U384 ( .A1(DP_mult_209_n556), .A2(DP_mult_209_n557), 
        .B1(DP_mult_209_n555), .B2(DP_mult_209_n558), .ZN(DP_mult_209_n304) );
  NOR2_X1 DP_mult_209_U383 ( .A1(DP_mult_209_n525), .A2(DP_mult_209_n555), 
        .ZN(DP_mult_209_n305) );
  AOI21_X1 DP_mult_209_U382 ( .B1(DP_mult_209_n542), .B2(DP_mult_209_n540), 
        .A(DP_mult_209_n554), .ZN(DP_mult_209_n553) );
  INV_X1 DP_mult_209_U381 ( .A(DP_mult_209_n553), .ZN(DP_mult_209_n306) );
  XNOR2_X1 DP_mult_209_U380 ( .A(DP_b_int_0__9_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n551) );
  OAI22_X1 DP_mult_209_U379 ( .A1(DP_mult_209_n551), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n552), .ZN(DP_mult_209_n307) );
  XNOR2_X1 DP_mult_209_U378 ( .A(DP_b_int_0__8_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n550) );
  OAI22_X1 DP_mult_209_U377 ( .A1(DP_mult_209_n550), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n551), .ZN(DP_mult_209_n308) );
  XNOR2_X1 DP_mult_209_U376 ( .A(DP_b_int_0__7_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n549) );
  OAI22_X1 DP_mult_209_U375 ( .A1(DP_mult_209_n549), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n550), .ZN(DP_mult_209_n309) );
  XNOR2_X1 DP_mult_209_U374 ( .A(DP_b_int_0__6_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n548) );
  OAI22_X1 DP_mult_209_U373 ( .A1(DP_mult_209_n548), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n549), .ZN(DP_mult_209_n310) );
  XNOR2_X1 DP_mult_209_U372 ( .A(DP_b_int_0__5_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n547) );
  OAI22_X1 DP_mult_209_U371 ( .A1(DP_mult_209_n547), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n548), .ZN(DP_mult_209_n311) );
  XNOR2_X1 DP_mult_209_U370 ( .A(DP_b_int_0__4_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n546) );
  OAI22_X1 DP_mult_209_U369 ( .A1(DP_mult_209_n546), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n547), .ZN(DP_mult_209_n312) );
  XNOR2_X1 DP_mult_209_U368 ( .A(DP_b_int_0__3_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n545) );
  OAI22_X1 DP_mult_209_U367 ( .A1(DP_mult_209_n545), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n546), .ZN(DP_mult_209_n313) );
  XNOR2_X1 DP_mult_209_U366 ( .A(DP_b_int_0__2_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n544) );
  OAI22_X1 DP_mult_209_U365 ( .A1(DP_mult_209_n544), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n545), .ZN(DP_mult_209_n314) );
  XNOR2_X1 DP_mult_209_U364 ( .A(DP_b_int_0__1_), .B(DP_mult_209_n515), .ZN(
        DP_mult_209_n543) );
  OAI22_X1 DP_mult_209_U363 ( .A1(DP_mult_209_n543), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n544), .ZN(DP_mult_209_n315) );
  XNOR2_X1 DP_mult_209_U362 ( .A(DP_mult_209_n515), .B(DP_b_int_0__0_), .ZN(
        DP_mult_209_n541) );
  OAI22_X1 DP_mult_209_U361 ( .A1(DP_mult_209_n541), .A2(DP_mult_209_n542), 
        .B1(DP_mult_209_n540), .B2(DP_mult_209_n543), .ZN(DP_mult_209_n316) );
  NOR2_X1 DP_mult_209_U360 ( .A1(DP_mult_209_n525), .A2(DP_mult_209_n540), 
        .ZN(DP_mult_209_n317) );
  XNOR2_X1 DP_mult_209_U359 ( .A(DP_b_int_0__11_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n538) );
  AOI21_X1 DP_mult_209_U358 ( .B1(DP_mult_209_n527), .B2(DP_mult_209_n526), 
        .A(DP_mult_209_n538), .ZN(DP_mult_209_n539) );
  INV_X1 DP_mult_209_U357 ( .A(DP_mult_209_n539), .ZN(DP_mult_209_n318) );
  XNOR2_X1 DP_mult_209_U356 ( .A(DP_b_int_0__10_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n537) );
  OAI22_X1 DP_mult_209_U355 ( .A1(DP_mult_209_n537), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n538), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n319) );
  XNOR2_X1 DP_mult_209_U354 ( .A(DP_b_int_0__9_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n536) );
  OAI22_X1 DP_mult_209_U353 ( .A1(DP_mult_209_n536), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n537), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n320) );
  XNOR2_X1 DP_mult_209_U352 ( .A(DP_b_int_0__8_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n535) );
  OAI22_X1 DP_mult_209_U351 ( .A1(DP_mult_209_n535), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n536), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n321) );
  XNOR2_X1 DP_mult_209_U350 ( .A(DP_b_int_0__7_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n534) );
  OAI22_X1 DP_mult_209_U349 ( .A1(DP_mult_209_n534), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n535), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n322) );
  XNOR2_X1 DP_mult_209_U348 ( .A(DP_b_int_0__6_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n533) );
  OAI22_X1 DP_mult_209_U347 ( .A1(DP_mult_209_n533), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n534), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n323) );
  XNOR2_X1 DP_mult_209_U346 ( .A(DP_b_int_0__5_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n532) );
  OAI22_X1 DP_mult_209_U345 ( .A1(DP_mult_209_n532), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n533), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n324) );
  XNOR2_X1 DP_mult_209_U344 ( .A(DP_b_int_0__4_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n531) );
  OAI22_X1 DP_mult_209_U343 ( .A1(DP_mult_209_n531), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n532), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n325) );
  XNOR2_X1 DP_mult_209_U342 ( .A(DP_b_int_0__3_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n530) );
  OAI22_X1 DP_mult_209_U341 ( .A1(DP_mult_209_n530), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n531), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n326) );
  XNOR2_X1 DP_mult_209_U340 ( .A(DP_b_int_0__2_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n529) );
  OAI22_X1 DP_mult_209_U339 ( .A1(DP_mult_209_n529), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n530), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n327) );
  XNOR2_X1 DP_mult_209_U338 ( .A(DP_b_int_0__1_), .B(DP_mult_209_n513), .ZN(
        DP_mult_209_n528) );
  OAI22_X1 DP_mult_209_U337 ( .A1(DP_mult_209_n528), .A2(DP_mult_209_n527), 
        .B1(DP_mult_209_n529), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n328) );
  OAI22_X1 DP_mult_209_U336 ( .A1(DP_b_int_0__0_), .A2(DP_mult_209_n527), .B1(
        DP_mult_209_n528), .B2(DP_mult_209_n526), .ZN(DP_mult_209_n329) );
  NOR2_X1 DP_mult_209_U335 ( .A1(DP_mult_209_n525), .A2(DP_mult_209_n526), 
        .ZN(DP_coeff_pipe01[0]) );
  INV_X1 DP_mult_209_U334 ( .A(DP_mult_209_n120), .ZN(DP_N97) );
  INV_X1 DP_mult_209_U333 ( .A(DP_a_int_1__1_), .ZN(DP_mult_209_n514) );
  XOR2_X2 DP_mult_209_U332 ( .A(DP_a_int_1__10_), .B(DP_mult_209_n522), .Z(
        DP_mult_209_n600) );
  XOR2_X2 DP_mult_209_U331 ( .A(DP_a_int_1__8_), .B(DP_mult_209_n520), .Z(
        DP_mult_209_n585) );
  XOR2_X2 DP_mult_209_U330 ( .A(DP_a_int_1__6_), .B(DP_mult_209_n518), .Z(
        DP_mult_209_n570) );
  XOR2_X2 DP_mult_209_U329 ( .A(DP_a_int_1__4_), .B(DP_mult_209_n516), .Z(
        DP_mult_209_n555) );
  XOR2_X2 DP_mult_209_U328 ( .A(DP_a_int_1__2_), .B(DP_mult_209_n514), .Z(
        DP_mult_209_n540) );
  INV_X1 DP_mult_209_U327 ( .A(DP_a_int_1__5_), .ZN(DP_mult_209_n518) );
  INV_X1 DP_mult_209_U326 ( .A(DP_a_int_1__3_), .ZN(DP_mult_209_n516) );
  INV_X1 DP_mult_209_U325 ( .A(DP_a_int_1__9_), .ZN(DP_mult_209_n522) );
  INV_X1 DP_mult_209_U324 ( .A(DP_a_int_1__7_), .ZN(DP_mult_209_n520) );
  INV_X1 DP_mult_209_U323 ( .A(DP_a_int_1__11_), .ZN(DP_mult_209_n524) );
  INV_X1 DP_mult_209_U322 ( .A(DP_mult_209_n514), .ZN(DP_mult_209_n513) );
  INV_X1 DP_mult_209_U321 ( .A(DP_mult_209_n522), .ZN(DP_mult_209_n521) );
  INV_X1 DP_mult_209_U320 ( .A(DP_mult_209_n520), .ZN(DP_mult_209_n519) );
  INV_X1 DP_mult_209_U319 ( .A(DP_mult_209_n518), .ZN(DP_mult_209_n517) );
  INV_X1 DP_mult_209_U318 ( .A(DP_mult_209_n516), .ZN(DP_mult_209_n515) );
  INV_X1 DP_mult_209_U317 ( .A(DP_mult_209_n524), .ZN(DP_mult_209_n523) );
  HA_X1 DP_mult_209_U107 ( .A(DP_mult_209_n316), .B(DP_mult_209_n327), .CO(
        DP_mult_209_n250), .S(DP_mult_209_n251) );
  FA_X1 DP_mult_209_U106 ( .A(DP_mult_209_n326), .B(DP_mult_209_n305), .CI(
        DP_mult_209_n315), .CO(DP_mult_209_n248), .S(DP_mult_209_n249) );
  HA_X1 DP_mult_209_U105 ( .A(DP_mult_209_n255), .B(DP_mult_209_n304), .CO(
        DP_mult_209_n246), .S(DP_mult_209_n247) );
  FA_X1 DP_mult_209_U104 ( .A(DP_mult_209_n314), .B(DP_mult_209_n325), .CI(
        DP_mult_209_n247), .CO(DP_mult_209_n244), .S(DP_mult_209_n245) );
  FA_X1 DP_mult_209_U103 ( .A(DP_mult_209_n324), .B(DP_mult_209_n293), .CI(
        DP_mult_209_n313), .CO(DP_mult_209_n242), .S(DP_mult_209_n243) );
  FA_X1 DP_mult_209_U102 ( .A(DP_mult_209_n246), .B(DP_mult_209_n303), .CI(
        DP_mult_209_n243), .CO(DP_mult_209_n240), .S(DP_mult_209_n241) );
  HA_X1 DP_mult_209_U101 ( .A(DP_mult_209_n254), .B(DP_mult_209_n292), .CO(
        DP_mult_209_n238), .S(DP_mult_209_n239) );
  FA_X1 DP_mult_209_U100 ( .A(DP_mult_209_n302), .B(DP_mult_209_n323), .CI(
        DP_mult_209_n312), .CO(DP_mult_209_n236), .S(DP_mult_209_n237) );
  FA_X1 DP_mult_209_U99 ( .A(DP_mult_209_n242), .B(DP_mult_209_n239), .CI(
        DP_mult_209_n237), .CO(DP_mult_209_n234), .S(DP_mult_209_n235) );
  FA_X1 DP_mult_209_U98 ( .A(DP_mult_209_n301), .B(DP_mult_209_n281), .CI(
        DP_mult_209_n322), .CO(DP_mult_209_n232), .S(DP_mult_209_n233) );
  FA_X1 DP_mult_209_U97 ( .A(DP_mult_209_n291), .B(DP_mult_209_n311), .CI(
        DP_mult_209_n238), .CO(DP_mult_209_n230), .S(DP_mult_209_n231) );
  FA_X1 DP_mult_209_U96 ( .A(DP_mult_209_n233), .B(DP_mult_209_n236), .CI(
        DP_mult_209_n231), .CO(DP_mult_209_n228), .S(DP_mult_209_n229) );
  HA_X1 DP_mult_209_U95 ( .A(DP_mult_209_n253), .B(DP_mult_209_n280), .CO(
        DP_mult_209_n226), .S(DP_mult_209_n227) );
  FA_X1 DP_mult_209_U94 ( .A(DP_mult_209_n290), .B(DP_mult_209_n300), .CI(
        DP_mult_209_n310), .CO(DP_mult_209_n224), .S(DP_mult_209_n225) );
  FA_X1 DP_mult_209_U93 ( .A(DP_mult_209_n227), .B(DP_mult_209_n321), .CI(
        DP_mult_209_n232), .CO(DP_mult_209_n222), .S(DP_mult_209_n223) );
  FA_X1 DP_mult_209_U92 ( .A(DP_mult_209_n225), .B(DP_mult_209_n230), .CI(
        DP_mult_209_n223), .CO(DP_mult_209_n220), .S(DP_mult_209_n221) );
  FA_X1 DP_mult_209_U91 ( .A(DP_mult_209_n289), .B(DP_mult_209_n269), .CI(
        DP_mult_209_n320), .CO(DP_mult_209_n218), .S(DP_mult_209_n219) );
  FA_X1 DP_mult_209_U90 ( .A(DP_mult_209_n279), .B(DP_mult_209_n309), .CI(
        DP_mult_209_n299), .CO(DP_mult_209_n216), .S(DP_mult_209_n217) );
  FA_X1 DP_mult_209_U89 ( .A(DP_mult_209_n224), .B(DP_mult_209_n226), .CI(
        DP_mult_209_n219), .CO(DP_mult_209_n214), .S(DP_mult_209_n215) );
  FA_X1 DP_mult_209_U88 ( .A(DP_mult_209_n222), .B(DP_mult_209_n217), .CI(
        DP_mult_209_n215), .CO(DP_mult_209_n212), .S(DP_mult_209_n213) );
  HA_X1 DP_mult_209_U87 ( .A(DP_mult_209_n252), .B(DP_mult_209_n268), .CO(
        DP_mult_209_n210), .S(DP_mult_209_n211) );
  FA_X1 DP_mult_209_U86 ( .A(DP_mult_209_n278), .B(DP_mult_209_n298), .CI(
        DP_mult_209_n319), .CO(DP_mult_209_n208), .S(DP_mult_209_n209) );
  FA_X1 DP_mult_209_U85 ( .A(DP_mult_209_n288), .B(DP_mult_209_n308), .CI(
        DP_mult_209_n211), .CO(DP_mult_209_n206), .S(DP_mult_209_n207) );
  FA_X1 DP_mult_209_U84 ( .A(DP_mult_209_n216), .B(DP_mult_209_n218), .CI(
        DP_mult_209_n209), .CO(DP_mult_209_n204), .S(DP_mult_209_n205) );
  FA_X1 DP_mult_209_U83 ( .A(DP_mult_209_n214), .B(DP_mult_209_n207), .CI(
        DP_mult_209_n205), .CO(DP_mult_209_n202), .S(DP_mult_209_n203) );
  FA_X1 DP_mult_209_U80 ( .A(DP_mult_209_n267), .B(DP_mult_209_n287), .CI(
        DP_mult_209_n318), .CO(DP_mult_209_n198), .S(DP_mult_209_n199) );
  FA_X1 DP_mult_209_U79 ( .A(DP_mult_209_n210), .B(DP_mult_209_n307), .CI(
        DP_mult_209_n201), .CO(DP_mult_209_n196), .S(DP_mult_209_n197) );
  FA_X1 DP_mult_209_U78 ( .A(DP_mult_209_n199), .B(DP_mult_209_n208), .CI(
        DP_mult_209_n206), .CO(DP_mult_209_n194), .S(DP_mult_209_n195) );
  FA_X1 DP_mult_209_U77 ( .A(DP_mult_209_n204), .B(DP_mult_209_n197), .CI(
        DP_mult_209_n195), .CO(DP_mult_209_n192), .S(DP_mult_209_n193) );
  FA_X1 DP_mult_209_U75 ( .A(DP_mult_209_n296), .B(DP_mult_209_n276), .CI(
        DP_mult_209_n191), .CO(DP_mult_209_n188), .S(DP_mult_209_n189) );
  FA_X1 DP_mult_209_U74 ( .A(DP_mult_209_n266), .B(DP_mult_209_n286), .CI(
        DP_mult_209_n200), .CO(DP_mult_209_n186), .S(DP_mult_209_n187) );
  FA_X1 DP_mult_209_U73 ( .A(DP_mult_209_n196), .B(DP_mult_209_n198), .CI(
        DP_mult_209_n189), .CO(DP_mult_209_n184), .S(DP_mult_209_n185) );
  FA_X1 DP_mult_209_U72 ( .A(DP_mult_209_n194), .B(DP_mult_209_n187), .CI(
        DP_mult_209_n185), .CO(DP_mult_209_n182), .S(DP_mult_209_n183) );
  FA_X1 DP_mult_209_U71 ( .A(DP_mult_209_n190), .B(DP_mult_209_n265), .CI(
        DP_mult_209_n306), .CO(DP_mult_209_n180), .S(DP_mult_209_n181) );
  FA_X1 DP_mult_209_U70 ( .A(DP_mult_209_n275), .B(DP_mult_209_n295), .CI(
        DP_mult_209_n285), .CO(DP_mult_209_n178), .S(DP_mult_209_n179) );
  FA_X1 DP_mult_209_U69 ( .A(DP_mult_209_n186), .B(DP_mult_209_n188), .CI(
        DP_mult_209_n179), .CO(DP_mult_209_n176), .S(DP_mult_209_n177) );
  FA_X1 DP_mult_209_U68 ( .A(DP_mult_209_n184), .B(DP_mult_209_n181), .CI(
        DP_mult_209_n177), .CO(DP_mult_209_n174), .S(DP_mult_209_n175) );
  FA_X1 DP_mult_209_U66 ( .A(DP_mult_209_n264), .B(DP_mult_209_n274), .CI(
        DP_mult_209_n173), .CO(DP_mult_209_n170), .S(DP_mult_209_n171) );
  FA_X1 DP_mult_209_U65 ( .A(DP_mult_209_n180), .B(DP_mult_209_n284), .CI(
        DP_mult_209_n178), .CO(DP_mult_209_n168), .S(DP_mult_209_n169) );
  FA_X1 DP_mult_209_U64 ( .A(DP_mult_209_n176), .B(DP_mult_209_n171), .CI(
        DP_mult_209_n169), .CO(DP_mult_209_n166), .S(DP_mult_209_n167) );
  FA_X1 DP_mult_209_U63 ( .A(DP_mult_209_n172), .B(DP_mult_209_n263), .CI(
        DP_mult_209_n294), .CO(DP_mult_209_n164), .S(DP_mult_209_n165) );
  FA_X1 DP_mult_209_U62 ( .A(DP_mult_209_n273), .B(DP_mult_209_n283), .CI(
        DP_mult_209_n170), .CO(DP_mult_209_n162), .S(DP_mult_209_n163) );
  FA_X1 DP_mult_209_U61 ( .A(DP_mult_209_n168), .B(DP_mult_209_n165), .CI(
        DP_mult_209_n163), .CO(DP_mult_209_n160), .S(DP_mult_209_n161) );
  FA_X1 DP_mult_209_U59 ( .A(DP_mult_209_n262), .B(DP_mult_209_n272), .CI(
        DP_mult_209_n159), .CO(DP_mult_209_n156), .S(DP_mult_209_n157) );
  FA_X1 DP_mult_209_U58 ( .A(DP_mult_209_n157), .B(DP_mult_209_n164), .CI(
        DP_mult_209_n162), .CO(DP_mult_209_n154), .S(DP_mult_209_n155) );
  FA_X1 DP_mult_209_U57 ( .A(DP_mult_209_n261), .B(DP_mult_209_n158), .CI(
        DP_mult_209_n282), .CO(DP_mult_209_n152), .S(DP_mult_209_n153) );
  FA_X1 DP_mult_209_U56 ( .A(DP_mult_209_n156), .B(DP_mult_209_n271), .CI(
        DP_mult_209_n153), .CO(DP_mult_209_n150), .S(DP_mult_209_n151) );
  FA_X1 DP_mult_209_U54 ( .A(DP_mult_209_n149), .B(DP_mult_209_n260), .CI(
        DP_mult_209_n152), .CO(DP_mult_209_n146), .S(DP_mult_209_n147) );
  FA_X1 DP_mult_209_U53 ( .A(DP_mult_209_n259), .B(DP_mult_209_n148), .CI(
        DP_mult_209_n270), .CO(DP_mult_209_n144), .S(DP_mult_209_n145) );
  HA_X1 DP_mult_209_U51 ( .A(DP_mult_209_n329), .B(DP_mult_209_n257), .CO(
        DP_mult_209_n141), .S(DP_N75) );
  FA_X1 DP_mult_209_U50 ( .A(DP_mult_209_n328), .B(DP_mult_209_n317), .CI(
        DP_mult_209_n141), .CO(DP_mult_209_n140), .S(DP_N76) );
  FA_X1 DP_mult_209_U49 ( .A(DP_mult_209_n251), .B(DP_mult_209_n256), .CI(
        DP_mult_209_n140), .CO(DP_mult_209_n139), .S(DP_N77) );
  FA_X1 DP_mult_209_U48 ( .A(DP_mult_209_n249), .B(DP_mult_209_n250), .CI(
        DP_mult_209_n139), .CO(DP_mult_209_n138), .S(DP_N78) );
  FA_X1 DP_mult_209_U47 ( .A(DP_mult_209_n245), .B(DP_mult_209_n248), .CI(
        DP_mult_209_n138), .CO(DP_mult_209_n137), .S(DP_N79) );
  FA_X1 DP_mult_209_U46 ( .A(DP_mult_209_n241), .B(DP_mult_209_n244), .CI(
        DP_mult_209_n137), .CO(DP_mult_209_n136), .S(DP_N80) );
  FA_X1 DP_mult_209_U45 ( .A(DP_mult_209_n235), .B(DP_mult_209_n240), .CI(
        DP_mult_209_n136), .CO(DP_mult_209_n135), .S(DP_N81) );
  FA_X1 DP_mult_209_U44 ( .A(DP_mult_209_n229), .B(DP_mult_209_n234), .CI(
        DP_mult_209_n135), .CO(DP_mult_209_n134), .S(DP_N82) );
  FA_X1 DP_mult_209_U43 ( .A(DP_mult_209_n221), .B(DP_mult_209_n228), .CI(
        DP_mult_209_n134), .CO(DP_mult_209_n133), .S(DP_N83) );
  FA_X1 DP_mult_209_U42 ( .A(DP_mult_209_n213), .B(DP_mult_209_n220), .CI(
        DP_mult_209_n133), .CO(DP_mult_209_n132), .S(DP_N84) );
  FA_X1 DP_mult_209_U41 ( .A(DP_mult_209_n203), .B(DP_mult_209_n212), .CI(
        DP_mult_209_n132), .CO(DP_mult_209_n131), .S(DP_N85) );
  FA_X1 DP_mult_209_U40 ( .A(DP_mult_209_n193), .B(DP_mult_209_n202), .CI(
        DP_mult_209_n131), .CO(DP_mult_209_n130), .S(DP_N86) );
  FA_X1 DP_mult_209_U39 ( .A(DP_mult_209_n183), .B(DP_mult_209_n192), .CI(
        DP_mult_209_n130), .CO(DP_mult_209_n129), .S(DP_N87) );
  FA_X1 DP_mult_209_U38 ( .A(DP_mult_209_n175), .B(DP_mult_209_n182), .CI(
        DP_mult_209_n129), .CO(DP_mult_209_n128), .S(DP_N88) );
  FA_X1 DP_mult_209_U37 ( .A(DP_mult_209_n167), .B(DP_mult_209_n174), .CI(
        DP_mult_209_n128), .CO(DP_mult_209_n127), .S(DP_N89) );
  FA_X1 DP_mult_209_U36 ( .A(DP_mult_209_n161), .B(DP_mult_209_n166), .CI(
        DP_mult_209_n127), .CO(DP_mult_209_n126), .S(DP_N90) );
  FA_X1 DP_mult_209_U30 ( .A(DP_mult_209_n160), .B(DP_mult_209_n155), .CI(
        DP_mult_209_n126), .CO(DP_mult_209_n125), .S(DP_N91) );
  FA_X1 DP_mult_209_U20 ( .A(DP_mult_209_n151), .B(DP_mult_209_n154), .CI(
        DP_mult_209_n125), .CO(DP_mult_209_n124), .S(DP_N92) );
  FA_X1 DP_mult_209_U10 ( .A(DP_mult_209_n147), .B(DP_mult_209_n150), .CI(
        DP_mult_209_n124), .CO(DP_mult_209_n123), .S(DP_N93) );
  FA_X1 DP_mult_209_U9 ( .A(DP_mult_209_n146), .B(DP_mult_209_n145), .CI(
        DP_mult_209_n123), .CO(DP_mult_209_n122), .S(DP_N94) );
  FA_X1 DP_mult_209_U8 ( .A(DP_mult_209_n144), .B(DP_mult_209_n143), .CI(
        DP_mult_209_n122), .CO(DP_mult_209_n121), .S(DP_N95) );
  FA_X1 DP_mult_209_U7 ( .A(DP_mult_209_n258), .B(DP_mult_209_n142), .CI(
        DP_mult_209_n121), .CO(DP_mult_209_n120), .S(DP_N96) );
  INV_X1 DP_sub_209_U44 ( .A(DP_N84), .ZN(DP_sub_209_B_not_10_) );
  INV_X1 DP_sub_209_U43 ( .A(DP_N85), .ZN(DP_sub_209_B_not_11_) );
  INV_X1 DP_sub_209_U42 ( .A(DP_N86), .ZN(DP_sub_209_B_not_12_) );
  INV_X1 DP_sub_209_U41 ( .A(DP_N87), .ZN(DP_sub_209_B_not_13_) );
  INV_X1 DP_sub_209_U40 ( .A(DP_N88), .ZN(DP_sub_209_B_not_14_) );
  INV_X1 DP_sub_209_U39 ( .A(DP_N89), .ZN(DP_sub_209_B_not_15_) );
  INV_X1 DP_sub_209_U38 ( .A(DP_N90), .ZN(DP_sub_209_B_not_16_) );
  INV_X1 DP_sub_209_U37 ( .A(DP_N91), .ZN(DP_sub_209_B_not_17_) );
  INV_X1 DP_sub_209_U36 ( .A(DP_N92), .ZN(DP_sub_209_B_not_18_) );
  INV_X1 DP_sub_209_U35 ( .A(DP_N93), .ZN(DP_sub_209_B_not_19_) );
  INV_X1 DP_sub_209_U34 ( .A(DP_N75), .ZN(DP_sub_209_B_not_1_) );
  INV_X1 DP_sub_209_U33 ( .A(DP_N94), .ZN(DP_sub_209_B_not_20_) );
  INV_X1 DP_sub_209_U32 ( .A(DP_N95), .ZN(DP_sub_209_B_not_21_) );
  INV_X1 DP_sub_209_U31 ( .A(DP_N96), .ZN(DP_sub_209_B_not_22_) );
  INV_X1 DP_sub_209_U30 ( .A(DP_N97), .ZN(DP_sub_209_B_not_23_) );
  INV_X1 DP_sub_209_U29 ( .A(DP_N76), .ZN(DP_sub_209_B_not_2_) );
  INV_X1 DP_sub_209_U28 ( .A(DP_N77), .ZN(DP_sub_209_B_not_3_) );
  INV_X1 DP_sub_209_U27 ( .A(DP_N78), .ZN(DP_sub_209_B_not_4_) );
  INV_X1 DP_sub_209_U26 ( .A(DP_N79), .ZN(DP_sub_209_B_not_5_) );
  INV_X1 DP_sub_209_U25 ( .A(DP_N80), .ZN(DP_sub_209_B_not_6_) );
  INV_X1 DP_sub_209_U24 ( .A(DP_N81), .ZN(DP_sub_209_B_not_7_) );
  INV_X1 DP_sub_209_U23 ( .A(DP_N82), .ZN(DP_sub_209_B_not_8_) );
  INV_X1 DP_sub_209_U22 ( .A(DP_N83), .ZN(DP_sub_209_B_not_9_) );
  INV_X1 DP_sub_209_U21 ( .A(DP_coeff_pipe01[0]), .ZN(DP_sub_209_carry_1_) );
  XOR2_X1 DP_sub_209_U20 ( .A(DP_sub_209_B_not_1_), .B(DP_sub_209_carry_1_), 
        .Z(DP_coeff_pipe01[1]) );
  AND2_X1 DP_sub_209_U19 ( .A1(DP_sub_209_carry_1_), .A2(DP_sub_209_B_not_1_), 
        .ZN(DP_sub_209_carry_2_) );
  AND2_X1 DP_sub_209_U18 ( .A1(DP_sub_209_carry_2_), .A2(DP_sub_209_B_not_2_), 
        .ZN(DP_sub_209_carry_3_) );
  XOR2_X1 DP_sub_209_U17 ( .A(DP_sub_209_B_not_3_), .B(DP_sub_209_carry_3_), 
        .Z(DP_coeff_pipe01[3]) );
  AND2_X1 DP_sub_209_U16 ( .A1(DP_sub_209_carry_3_), .A2(DP_sub_209_B_not_3_), 
        .ZN(DP_sub_209_carry_4_) );
  XOR2_X1 DP_sub_209_U15 ( .A(DP_sub_209_B_not_4_), .B(DP_sub_209_carry_4_), 
        .Z(DP_coeff_pipe01[4]) );
  AND2_X1 DP_sub_209_U14 ( .A1(DP_sub_209_carry_4_), .A2(DP_sub_209_B_not_4_), 
        .ZN(DP_sub_209_carry_5_) );
  XOR2_X1 DP_sub_209_U13 ( .A(DP_sub_209_B_not_5_), .B(DP_sub_209_carry_5_), 
        .Z(DP_coeff_pipe01[5]) );
  AND2_X1 DP_sub_209_U12 ( .A1(DP_sub_209_carry_5_), .A2(DP_sub_209_B_not_5_), 
        .ZN(DP_sub_209_carry_6_) );
  XOR2_X1 DP_sub_209_U11 ( .A(DP_sub_209_B_not_6_), .B(DP_sub_209_carry_6_), 
        .Z(DP_coeff_pipe01[6]) );
  AND2_X1 DP_sub_209_U10 ( .A1(DP_sub_209_carry_6_), .A2(DP_sub_209_B_not_6_), 
        .ZN(DP_sub_209_carry_7_) );
  XOR2_X1 DP_sub_209_U9 ( .A(DP_sub_209_B_not_7_), .B(DP_sub_209_carry_7_), 
        .Z(DP_coeff_pipe01[7]) );
  AND2_X1 DP_sub_209_U8 ( .A1(DP_sub_209_carry_7_), .A2(DP_sub_209_B_not_7_), 
        .ZN(DP_sub_209_carry_8_) );
  XOR2_X1 DP_sub_209_U7 ( .A(DP_sub_209_B_not_8_), .B(DP_sub_209_carry_8_), 
        .Z(DP_coeff_pipe01[8]) );
  AND2_X1 DP_sub_209_U6 ( .A1(DP_sub_209_carry_8_), .A2(DP_sub_209_B_not_8_), 
        .ZN(DP_sub_209_carry_9_) );
  XOR2_X1 DP_sub_209_U5 ( .A(DP_sub_209_B_not_9_), .B(DP_sub_209_carry_9_), 
        .Z(DP_coeff_pipe01[9]) );
  AND2_X1 DP_sub_209_U4 ( .A1(DP_sub_209_carry_9_), .A2(DP_sub_209_B_not_9_), 
        .ZN(DP_sub_209_carry_10_) );
  XOR2_X1 DP_sub_209_U3 ( .A(DP_sub_209_B_not_10_), .B(DP_sub_209_carry_10_), 
        .Z(DP_coeff_pipe01[10]) );
  AND2_X1 DP_sub_209_U2 ( .A1(DP_sub_209_carry_10_), .A2(DP_sub_209_B_not_10_), 
        .ZN(DP_sub_209_carry_11_) );
  XOR2_X2 DP_sub_209_U1 ( .A(DP_sub_209_B_not_2_), .B(DP_sub_209_carry_2_), 
        .Z(DP_coeff_pipe01[2]) );
  FA_X1 DP_sub_209_U2_11 ( .A(DP_b_int_1__0_), .B(DP_sub_209_B_not_11_), .CI(
        DP_sub_209_carry_11_), .CO(DP_sub_209_carry_12_), .S(
        DP_coeff_pipe01[11]) );
  FA_X1 DP_sub_209_U2_12 ( .A(DP_b_int_1__1_), .B(DP_sub_209_B_not_12_), .CI(
        DP_sub_209_carry_12_), .CO(DP_sub_209_carry_13_), .S(
        DP_coeff_pipe01[12]) );
  FA_X1 DP_sub_209_U2_13 ( .A(DP_b_int_1__2_), .B(DP_sub_209_B_not_13_), .CI(
        DP_sub_209_carry_13_), .CO(DP_sub_209_carry_14_), .S(
        DP_coeff_pipe01[13]) );
  FA_X1 DP_sub_209_U2_14 ( .A(DP_b_int_1__3_), .B(DP_sub_209_B_not_14_), .CI(
        DP_sub_209_carry_14_), .CO(DP_sub_209_carry_15_), .S(
        DP_coeff_pipe01[14]) );
  FA_X1 DP_sub_209_U2_15 ( .A(DP_b_int_1__4_), .B(DP_sub_209_B_not_15_), .CI(
        DP_sub_209_carry_15_), .CO(DP_sub_209_carry_16_), .S(
        DP_coeff_pipe01[15]) );
  FA_X1 DP_sub_209_U2_16 ( .A(DP_b_int_1__5_), .B(DP_sub_209_B_not_16_), .CI(
        DP_sub_209_carry_16_), .CO(DP_sub_209_carry_17_), .S(
        DP_coeff_pipe01[16]) );
  FA_X1 DP_sub_209_U2_17 ( .A(DP_b_int_1__6_), .B(DP_sub_209_B_not_17_), .CI(
        DP_sub_209_carry_17_), .CO(DP_sub_209_carry_18_), .S(
        DP_coeff_pipe01[17]) );
  FA_X1 DP_sub_209_U2_18 ( .A(DP_b_int_1__7_), .B(DP_sub_209_B_not_18_), .CI(
        DP_sub_209_carry_18_), .CO(DP_sub_209_carry_19_), .S(
        DP_coeff_pipe01[18]) );
  FA_X1 DP_sub_209_U2_19 ( .A(DP_b_int_1__8_), .B(DP_sub_209_B_not_19_), .CI(
        DP_sub_209_carry_19_), .CO(DP_sub_209_carry_20_), .S(
        DP_coeff_pipe01[19]) );
  FA_X1 DP_sub_209_U2_20 ( .A(DP_b_int_1__9_), .B(DP_sub_209_B_not_20_), .CI(
        DP_sub_209_carry_20_), .CO(DP_sub_209_carry_21_), .S(
        DP_coeff_pipe01[20]) );
  FA_X1 DP_sub_209_U2_21 ( .A(DP_b_int_1__10_), .B(DP_sub_209_B_not_21_), .CI(
        DP_sub_209_carry_21_), .CO(DP_sub_209_carry_22_), .S(
        DP_coeff_pipe01[21]) );
  FA_X1 DP_sub_209_U2_22 ( .A(DP_b_int_1__11_), .B(DP_sub_209_B_not_22_), .CI(
        DP_sub_209_carry_22_), .CO(DP_sub_209_carry_23_), .S(
        DP_coeff_pipe01[22]) );
  FA_X1 DP_sub_209_U2_23 ( .A(DP_b_int_1__11_), .B(DP_sub_209_B_not_23_), .CI(
        DP_sub_209_carry_23_), .S(DP_coeff_pipe01[23]) );
  XNOR2_X1 DP_mult_210_U520 ( .A(DP_b_int_1__10_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n612) );
  XNOR2_X1 DP_mult_210_U519 ( .A(DP_mult_210_n524), .B(DP_a_int_1__10_), .ZN(
        DP_mult_210_n626) );
  NAND2_X1 DP_mult_210_U518 ( .A1(DP_mult_210_n600), .A2(DP_mult_210_n626), 
        .ZN(DP_mult_210_n602) );
  XNOR2_X1 DP_mult_210_U517 ( .A(DP_b_int_1__11_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n614) );
  OAI22_X1 DP_mult_210_U516 ( .A1(DP_mult_210_n612), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n614), .ZN(DP_mult_210_n142) );
  INV_X1 DP_mult_210_U515 ( .A(DP_mult_210_n142), .ZN(DP_mult_210_n143) );
  XNOR2_X1 DP_mult_210_U514 ( .A(DP_b_int_1__10_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n597) );
  XNOR2_X1 DP_mult_210_U513 ( .A(DP_mult_210_n522), .B(DP_a_int_1__8_), .ZN(
        DP_mult_210_n625) );
  NAND2_X1 DP_mult_210_U512 ( .A1(DP_mult_210_n585), .A2(DP_mult_210_n625), 
        .ZN(DP_mult_210_n587) );
  XNOR2_X1 DP_mult_210_U511 ( .A(DP_b_int_1__11_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n599) );
  OAI22_X1 DP_mult_210_U510 ( .A1(DP_mult_210_n597), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n599), .ZN(DP_mult_210_n148) );
  INV_X1 DP_mult_210_U509 ( .A(DP_mult_210_n148), .ZN(DP_mult_210_n149) );
  XNOR2_X1 DP_mult_210_U508 ( .A(DP_b_int_1__10_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n582) );
  XNOR2_X1 DP_mult_210_U507 ( .A(DP_mult_210_n520), .B(DP_a_int_1__6_), .ZN(
        DP_mult_210_n624) );
  NAND2_X1 DP_mult_210_U506 ( .A1(DP_mult_210_n570), .A2(DP_mult_210_n624), 
        .ZN(DP_mult_210_n572) );
  XNOR2_X1 DP_mult_210_U505 ( .A(DP_b_int_1__11_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n584) );
  OAI22_X1 DP_mult_210_U504 ( .A1(DP_mult_210_n582), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n584), .ZN(DP_mult_210_n158) );
  INV_X1 DP_mult_210_U503 ( .A(DP_mult_210_n158), .ZN(DP_mult_210_n159) );
  XNOR2_X1 DP_mult_210_U502 ( .A(DP_b_int_1__10_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n567) );
  XNOR2_X1 DP_mult_210_U501 ( .A(DP_mult_210_n518), .B(DP_a_int_1__4_), .ZN(
        DP_mult_210_n623) );
  NAND2_X1 DP_mult_210_U500 ( .A1(DP_mult_210_n555), .A2(DP_mult_210_n623), 
        .ZN(DP_mult_210_n557) );
  XNOR2_X1 DP_mult_210_U499 ( .A(DP_b_int_1__11_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n569) );
  OAI22_X1 DP_mult_210_U498 ( .A1(DP_mult_210_n567), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n569), .ZN(DP_mult_210_n172) );
  INV_X1 DP_mult_210_U497 ( .A(DP_mult_210_n172), .ZN(DP_mult_210_n173) );
  XNOR2_X1 DP_mult_210_U496 ( .A(DP_b_int_1__10_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n552) );
  XNOR2_X1 DP_mult_210_U495 ( .A(DP_mult_210_n516), .B(DP_a_int_1__2_), .ZN(
        DP_mult_210_n622) );
  NAND2_X1 DP_mult_210_U494 ( .A1(DP_mult_210_n540), .A2(DP_mult_210_n622), 
        .ZN(DP_mult_210_n542) );
  XNOR2_X1 DP_mult_210_U493 ( .A(DP_b_int_1__11_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n554) );
  OAI22_X1 DP_mult_210_U492 ( .A1(DP_mult_210_n552), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n554), .ZN(DP_mult_210_n190) );
  INV_X1 DP_mult_210_U491 ( .A(DP_mult_210_n190), .ZN(DP_mult_210_n191) );
  XNOR2_X1 DP_mult_210_U490 ( .A(DP_b_int_1__3_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n590) );
  XNOR2_X1 DP_mult_210_U489 ( .A(DP_b_int_1__4_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n591) );
  OAI22_X1 DP_mult_210_U488 ( .A1(DP_mult_210_n590), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n591), .ZN(DP_mult_210_n620) );
  XNOR2_X1 DP_mult_210_U487 ( .A(DP_b_int_1__7_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n564) );
  XNOR2_X1 DP_mult_210_U486 ( .A(DP_b_int_1__8_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n565) );
  OAI22_X1 DP_mult_210_U485 ( .A1(DP_mult_210_n564), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n565), .ZN(DP_mult_210_n621) );
  OR2_X1 DP_mult_210_U484 ( .A1(DP_mult_210_n620), .A2(DP_mult_210_n621), .ZN(
        DP_mult_210_n200) );
  XNOR2_X1 DP_mult_210_U483 ( .A(DP_mult_210_n620), .B(DP_mult_210_n621), .ZN(
        DP_mult_210_n201) );
  OR3_X1 DP_mult_210_U482 ( .A1(DP_mult_210_n600), .A2(DP_b_int_1__0_), .A3(
        DP_mult_210_n524), .ZN(DP_mult_210_n619) );
  OAI21_X1 DP_mult_210_U481 ( .B1(DP_mult_210_n524), .B2(DP_mult_210_n602), 
        .A(DP_mult_210_n619), .ZN(DP_mult_210_n252) );
  OR3_X1 DP_mult_210_U480 ( .A1(DP_mult_210_n585), .A2(DP_b_int_1__0_), .A3(
        DP_mult_210_n522), .ZN(DP_mult_210_n618) );
  OAI21_X1 DP_mult_210_U479 ( .B1(DP_mult_210_n522), .B2(DP_mult_210_n587), 
        .A(DP_mult_210_n618), .ZN(DP_mult_210_n253) );
  OR3_X1 DP_mult_210_U478 ( .A1(DP_mult_210_n570), .A2(DP_b_int_1__0_), .A3(
        DP_mult_210_n520), .ZN(DP_mult_210_n617) );
  OAI21_X1 DP_mult_210_U477 ( .B1(DP_mult_210_n520), .B2(DP_mult_210_n572), 
        .A(DP_mult_210_n617), .ZN(DP_mult_210_n254) );
  OR3_X1 DP_mult_210_U476 ( .A1(DP_mult_210_n555), .A2(DP_b_int_1__0_), .A3(
        DP_mult_210_n518), .ZN(DP_mult_210_n616) );
  OAI21_X1 DP_mult_210_U475 ( .B1(DP_mult_210_n518), .B2(DP_mult_210_n557), 
        .A(DP_mult_210_n616), .ZN(DP_mult_210_n255) );
  OR3_X1 DP_mult_210_U474 ( .A1(DP_mult_210_n540), .A2(DP_b_int_1__0_), .A3(
        DP_mult_210_n516), .ZN(DP_mult_210_n615) );
  OAI21_X1 DP_mult_210_U473 ( .B1(DP_mult_210_n516), .B2(DP_mult_210_n542), 
        .A(DP_mult_210_n615), .ZN(DP_mult_210_n256) );
  INV_X1 DP_mult_210_U472 ( .A(DP_coeff_ret0[1]), .ZN(DP_mult_210_n526) );
  NAND2_X1 DP_mult_210_U471 ( .A1(DP_mult_210_n513), .A2(DP_mult_210_n526), 
        .ZN(DP_mult_210_n527) );
  OAI21_X1 DP_mult_210_U470 ( .B1(DP_b_int_1__0_), .B2(DP_mult_210_n514), .A(
        DP_mult_210_n527), .ZN(DP_mult_210_n257) );
  AOI21_X1 DP_mult_210_U469 ( .B1(DP_mult_210_n602), .B2(DP_mult_210_n600), 
        .A(DP_mult_210_n614), .ZN(DP_mult_210_n613) );
  INV_X1 DP_mult_210_U468 ( .A(DP_mult_210_n613), .ZN(DP_mult_210_n258) );
  XNOR2_X1 DP_mult_210_U467 ( .A(DP_b_int_1__9_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n611) );
  OAI22_X1 DP_mult_210_U466 ( .A1(DP_mult_210_n611), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n612), .ZN(DP_mult_210_n259) );
  XNOR2_X1 DP_mult_210_U465 ( .A(DP_b_int_1__8_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n610) );
  OAI22_X1 DP_mult_210_U464 ( .A1(DP_mult_210_n610), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n611), .ZN(DP_mult_210_n260) );
  XNOR2_X1 DP_mult_210_U463 ( .A(DP_b_int_1__7_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n609) );
  OAI22_X1 DP_mult_210_U462 ( .A1(DP_mult_210_n609), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n610), .ZN(DP_mult_210_n261) );
  XNOR2_X1 DP_mult_210_U461 ( .A(DP_b_int_1__6_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n608) );
  OAI22_X1 DP_mult_210_U460 ( .A1(DP_mult_210_n608), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n609), .ZN(DP_mult_210_n262) );
  XNOR2_X1 DP_mult_210_U459 ( .A(DP_b_int_1__5_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n607) );
  OAI22_X1 DP_mult_210_U458 ( .A1(DP_mult_210_n607), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n608), .ZN(DP_mult_210_n263) );
  XNOR2_X1 DP_mult_210_U457 ( .A(DP_b_int_1__4_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n606) );
  OAI22_X1 DP_mult_210_U456 ( .A1(DP_mult_210_n606), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n607), .ZN(DP_mult_210_n264) );
  XNOR2_X1 DP_mult_210_U455 ( .A(DP_b_int_1__3_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n605) );
  OAI22_X1 DP_mult_210_U454 ( .A1(DP_mult_210_n605), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n606), .ZN(DP_mult_210_n265) );
  XNOR2_X1 DP_mult_210_U453 ( .A(DP_b_int_1__2_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n604) );
  OAI22_X1 DP_mult_210_U452 ( .A1(DP_mult_210_n604), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n605), .ZN(DP_mult_210_n266) );
  XNOR2_X1 DP_mult_210_U451 ( .A(DP_b_int_1__1_), .B(DP_mult_210_n523), .ZN(
        DP_mult_210_n603) );
  OAI22_X1 DP_mult_210_U450 ( .A1(DP_mult_210_n603), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n604), .ZN(DP_mult_210_n267) );
  XNOR2_X1 DP_mult_210_U449 ( .A(DP_mult_210_n523), .B(DP_b_int_1__0_), .ZN(
        DP_mult_210_n601) );
  OAI22_X1 DP_mult_210_U448 ( .A1(DP_mult_210_n601), .A2(DP_mult_210_n602), 
        .B1(DP_mult_210_n600), .B2(DP_mult_210_n603), .ZN(DP_mult_210_n268) );
  INV_X1 DP_mult_210_U447 ( .A(DP_b_int_1__0_), .ZN(DP_mult_210_n525) );
  NOR2_X1 DP_mult_210_U446 ( .A1(DP_mult_210_n525), .A2(DP_mult_210_n600), 
        .ZN(DP_mult_210_n269) );
  AOI21_X1 DP_mult_210_U445 ( .B1(DP_mult_210_n587), .B2(DP_mult_210_n585), 
        .A(DP_mult_210_n599), .ZN(DP_mult_210_n598) );
  INV_X1 DP_mult_210_U444 ( .A(DP_mult_210_n598), .ZN(DP_mult_210_n270) );
  XNOR2_X1 DP_mult_210_U443 ( .A(DP_b_int_1__9_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n596) );
  OAI22_X1 DP_mult_210_U442 ( .A1(DP_mult_210_n596), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n597), .ZN(DP_mult_210_n271) );
  XNOR2_X1 DP_mult_210_U441 ( .A(DP_b_int_1__8_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n595) );
  OAI22_X1 DP_mult_210_U440 ( .A1(DP_mult_210_n595), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n596), .ZN(DP_mult_210_n272) );
  XNOR2_X1 DP_mult_210_U439 ( .A(DP_b_int_1__7_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n594) );
  OAI22_X1 DP_mult_210_U438 ( .A1(DP_mult_210_n594), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n595), .ZN(DP_mult_210_n273) );
  XNOR2_X1 DP_mult_210_U437 ( .A(DP_b_int_1__6_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n593) );
  OAI22_X1 DP_mult_210_U436 ( .A1(DP_mult_210_n593), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n594), .ZN(DP_mult_210_n274) );
  XNOR2_X1 DP_mult_210_U435 ( .A(DP_b_int_1__5_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n592) );
  OAI22_X1 DP_mult_210_U434 ( .A1(DP_mult_210_n592), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n593), .ZN(DP_mult_210_n275) );
  OAI22_X1 DP_mult_210_U433 ( .A1(DP_mult_210_n591), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n592), .ZN(DP_mult_210_n276) );
  XNOR2_X1 DP_mult_210_U432 ( .A(DP_b_int_1__2_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n589) );
  OAI22_X1 DP_mult_210_U431 ( .A1(DP_mult_210_n589), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n590), .ZN(DP_mult_210_n278) );
  XNOR2_X1 DP_mult_210_U430 ( .A(DP_b_int_1__1_), .B(DP_mult_210_n521), .ZN(
        DP_mult_210_n588) );
  OAI22_X1 DP_mult_210_U429 ( .A1(DP_mult_210_n588), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n589), .ZN(DP_mult_210_n279) );
  XNOR2_X1 DP_mult_210_U428 ( .A(DP_mult_210_n521), .B(DP_b_int_1__0_), .ZN(
        DP_mult_210_n586) );
  OAI22_X1 DP_mult_210_U427 ( .A1(DP_mult_210_n586), .A2(DP_mult_210_n587), 
        .B1(DP_mult_210_n585), .B2(DP_mult_210_n588), .ZN(DP_mult_210_n280) );
  NOR2_X1 DP_mult_210_U426 ( .A1(DP_mult_210_n525), .A2(DP_mult_210_n585), 
        .ZN(DP_mult_210_n281) );
  AOI21_X1 DP_mult_210_U425 ( .B1(DP_mult_210_n572), .B2(DP_mult_210_n570), 
        .A(DP_mult_210_n584), .ZN(DP_mult_210_n583) );
  INV_X1 DP_mult_210_U424 ( .A(DP_mult_210_n583), .ZN(DP_mult_210_n282) );
  XNOR2_X1 DP_mult_210_U423 ( .A(DP_b_int_1__9_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n581) );
  OAI22_X1 DP_mult_210_U422 ( .A1(DP_mult_210_n581), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n582), .ZN(DP_mult_210_n283) );
  XNOR2_X1 DP_mult_210_U421 ( .A(DP_b_int_1__8_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n580) );
  OAI22_X1 DP_mult_210_U420 ( .A1(DP_mult_210_n580), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n581), .ZN(DP_mult_210_n284) );
  XNOR2_X1 DP_mult_210_U419 ( .A(DP_b_int_1__7_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n579) );
  OAI22_X1 DP_mult_210_U418 ( .A1(DP_mult_210_n579), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n580), .ZN(DP_mult_210_n285) );
  XNOR2_X1 DP_mult_210_U417 ( .A(DP_b_int_1__6_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n578) );
  OAI22_X1 DP_mult_210_U416 ( .A1(DP_mult_210_n578), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n579), .ZN(DP_mult_210_n286) );
  XNOR2_X1 DP_mult_210_U415 ( .A(DP_b_int_1__5_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n577) );
  OAI22_X1 DP_mult_210_U414 ( .A1(DP_mult_210_n577), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n578), .ZN(DP_mult_210_n287) );
  XNOR2_X1 DP_mult_210_U413 ( .A(DP_b_int_1__4_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n576) );
  OAI22_X1 DP_mult_210_U412 ( .A1(DP_mult_210_n576), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n577), .ZN(DP_mult_210_n288) );
  XNOR2_X1 DP_mult_210_U411 ( .A(DP_b_int_1__3_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n575) );
  OAI22_X1 DP_mult_210_U410 ( .A1(DP_mult_210_n575), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n576), .ZN(DP_mult_210_n289) );
  XNOR2_X1 DP_mult_210_U409 ( .A(DP_b_int_1__2_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n574) );
  OAI22_X1 DP_mult_210_U408 ( .A1(DP_mult_210_n574), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n575), .ZN(DP_mult_210_n290) );
  XNOR2_X1 DP_mult_210_U407 ( .A(DP_b_int_1__1_), .B(DP_mult_210_n519), .ZN(
        DP_mult_210_n573) );
  OAI22_X1 DP_mult_210_U406 ( .A1(DP_mult_210_n573), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n574), .ZN(DP_mult_210_n291) );
  XNOR2_X1 DP_mult_210_U405 ( .A(DP_mult_210_n519), .B(DP_b_int_1__0_), .ZN(
        DP_mult_210_n571) );
  OAI22_X1 DP_mult_210_U404 ( .A1(DP_mult_210_n571), .A2(DP_mult_210_n572), 
        .B1(DP_mult_210_n570), .B2(DP_mult_210_n573), .ZN(DP_mult_210_n292) );
  NOR2_X1 DP_mult_210_U403 ( .A1(DP_mult_210_n525), .A2(DP_mult_210_n570), 
        .ZN(DP_mult_210_n293) );
  AOI21_X1 DP_mult_210_U402 ( .B1(DP_mult_210_n557), .B2(DP_mult_210_n555), 
        .A(DP_mult_210_n569), .ZN(DP_mult_210_n568) );
  INV_X1 DP_mult_210_U401 ( .A(DP_mult_210_n568), .ZN(DP_mult_210_n294) );
  XNOR2_X1 DP_mult_210_U400 ( .A(DP_b_int_1__9_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n566) );
  OAI22_X1 DP_mult_210_U399 ( .A1(DP_mult_210_n566), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n567), .ZN(DP_mult_210_n295) );
  OAI22_X1 DP_mult_210_U398 ( .A1(DP_mult_210_n565), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n566), .ZN(DP_mult_210_n296) );
  XNOR2_X1 DP_mult_210_U397 ( .A(DP_b_int_1__6_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n563) );
  OAI22_X1 DP_mult_210_U396 ( .A1(DP_mult_210_n563), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n564), .ZN(DP_mult_210_n298) );
  XNOR2_X1 DP_mult_210_U395 ( .A(DP_b_int_1__5_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n562) );
  OAI22_X1 DP_mult_210_U394 ( .A1(DP_mult_210_n562), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n563), .ZN(DP_mult_210_n299) );
  XNOR2_X1 DP_mult_210_U393 ( .A(DP_b_int_1__4_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n561) );
  OAI22_X1 DP_mult_210_U392 ( .A1(DP_mult_210_n561), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n562), .ZN(DP_mult_210_n300) );
  XNOR2_X1 DP_mult_210_U391 ( .A(DP_b_int_1__3_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n560) );
  OAI22_X1 DP_mult_210_U390 ( .A1(DP_mult_210_n560), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n561), .ZN(DP_mult_210_n301) );
  XNOR2_X1 DP_mult_210_U389 ( .A(DP_b_int_1__2_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n559) );
  OAI22_X1 DP_mult_210_U388 ( .A1(DP_mult_210_n559), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n560), .ZN(DP_mult_210_n302) );
  XNOR2_X1 DP_mult_210_U387 ( .A(DP_b_int_1__1_), .B(DP_mult_210_n517), .ZN(
        DP_mult_210_n558) );
  OAI22_X1 DP_mult_210_U386 ( .A1(DP_mult_210_n558), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n559), .ZN(DP_mult_210_n303) );
  XNOR2_X1 DP_mult_210_U385 ( .A(DP_mult_210_n517), .B(DP_b_int_1__0_), .ZN(
        DP_mult_210_n556) );
  OAI22_X1 DP_mult_210_U384 ( .A1(DP_mult_210_n556), .A2(DP_mult_210_n557), 
        .B1(DP_mult_210_n555), .B2(DP_mult_210_n558), .ZN(DP_mult_210_n304) );
  NOR2_X1 DP_mult_210_U383 ( .A1(DP_mult_210_n525), .A2(DP_mult_210_n555), 
        .ZN(DP_mult_210_n305) );
  AOI21_X1 DP_mult_210_U382 ( .B1(DP_mult_210_n542), .B2(DP_mult_210_n540), 
        .A(DP_mult_210_n554), .ZN(DP_mult_210_n553) );
  INV_X1 DP_mult_210_U381 ( .A(DP_mult_210_n553), .ZN(DP_mult_210_n306) );
  XNOR2_X1 DP_mult_210_U380 ( .A(DP_b_int_1__9_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n551) );
  OAI22_X1 DP_mult_210_U379 ( .A1(DP_mult_210_n551), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n552), .ZN(DP_mult_210_n307) );
  XNOR2_X1 DP_mult_210_U378 ( .A(DP_b_int_1__8_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n550) );
  OAI22_X1 DP_mult_210_U377 ( .A1(DP_mult_210_n550), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n551), .ZN(DP_mult_210_n308) );
  XNOR2_X1 DP_mult_210_U376 ( .A(DP_b_int_1__7_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n549) );
  OAI22_X1 DP_mult_210_U375 ( .A1(DP_mult_210_n549), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n550), .ZN(DP_mult_210_n309) );
  XNOR2_X1 DP_mult_210_U374 ( .A(DP_b_int_1__6_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n548) );
  OAI22_X1 DP_mult_210_U373 ( .A1(DP_mult_210_n548), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n549), .ZN(DP_mult_210_n310) );
  XNOR2_X1 DP_mult_210_U372 ( .A(DP_b_int_1__5_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n547) );
  OAI22_X1 DP_mult_210_U371 ( .A1(DP_mult_210_n547), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n548), .ZN(DP_mult_210_n311) );
  XNOR2_X1 DP_mult_210_U370 ( .A(DP_b_int_1__4_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n546) );
  OAI22_X1 DP_mult_210_U369 ( .A1(DP_mult_210_n546), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n547), .ZN(DP_mult_210_n312) );
  XNOR2_X1 DP_mult_210_U368 ( .A(DP_b_int_1__3_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n545) );
  OAI22_X1 DP_mult_210_U367 ( .A1(DP_mult_210_n545), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n546), .ZN(DP_mult_210_n313) );
  XNOR2_X1 DP_mult_210_U366 ( .A(DP_b_int_1__2_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n544) );
  OAI22_X1 DP_mult_210_U365 ( .A1(DP_mult_210_n544), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n545), .ZN(DP_mult_210_n314) );
  XNOR2_X1 DP_mult_210_U364 ( .A(DP_b_int_1__1_), .B(DP_mult_210_n515), .ZN(
        DP_mult_210_n543) );
  OAI22_X1 DP_mult_210_U363 ( .A1(DP_mult_210_n543), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n544), .ZN(DP_mult_210_n315) );
  XNOR2_X1 DP_mult_210_U362 ( .A(DP_mult_210_n515), .B(DP_b_int_1__0_), .ZN(
        DP_mult_210_n541) );
  OAI22_X1 DP_mult_210_U361 ( .A1(DP_mult_210_n541), .A2(DP_mult_210_n542), 
        .B1(DP_mult_210_n540), .B2(DP_mult_210_n543), .ZN(DP_mult_210_n316) );
  NOR2_X1 DP_mult_210_U360 ( .A1(DP_mult_210_n525), .A2(DP_mult_210_n540), 
        .ZN(DP_mult_210_n317) );
  XNOR2_X1 DP_mult_210_U359 ( .A(DP_b_int_1__11_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n538) );
  AOI21_X1 DP_mult_210_U358 ( .B1(DP_mult_210_n527), .B2(DP_mult_210_n526), 
        .A(DP_mult_210_n538), .ZN(DP_mult_210_n539) );
  INV_X1 DP_mult_210_U357 ( .A(DP_mult_210_n539), .ZN(DP_mult_210_n318) );
  XNOR2_X1 DP_mult_210_U356 ( .A(DP_b_int_1__10_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n537) );
  OAI22_X1 DP_mult_210_U355 ( .A1(DP_mult_210_n537), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n538), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n319) );
  XNOR2_X1 DP_mult_210_U354 ( .A(DP_b_int_1__9_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n536) );
  OAI22_X1 DP_mult_210_U353 ( .A1(DP_mult_210_n536), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n537), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n320) );
  XNOR2_X1 DP_mult_210_U352 ( .A(DP_b_int_1__8_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n535) );
  OAI22_X1 DP_mult_210_U351 ( .A1(DP_mult_210_n535), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n536), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n321) );
  XNOR2_X1 DP_mult_210_U350 ( .A(DP_b_int_1__7_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n534) );
  OAI22_X1 DP_mult_210_U349 ( .A1(DP_mult_210_n534), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n535), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n322) );
  XNOR2_X1 DP_mult_210_U348 ( .A(DP_b_int_1__6_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n533) );
  OAI22_X1 DP_mult_210_U347 ( .A1(DP_mult_210_n533), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n534), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n323) );
  XNOR2_X1 DP_mult_210_U346 ( .A(DP_b_int_1__5_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n532) );
  OAI22_X1 DP_mult_210_U345 ( .A1(DP_mult_210_n532), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n533), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n324) );
  XNOR2_X1 DP_mult_210_U344 ( .A(DP_b_int_1__4_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n531) );
  OAI22_X1 DP_mult_210_U343 ( .A1(DP_mult_210_n531), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n532), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n325) );
  XNOR2_X1 DP_mult_210_U342 ( .A(DP_b_int_1__3_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n530) );
  OAI22_X1 DP_mult_210_U341 ( .A1(DP_mult_210_n530), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n531), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n326) );
  XNOR2_X1 DP_mult_210_U340 ( .A(DP_b_int_1__2_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n529) );
  OAI22_X1 DP_mult_210_U339 ( .A1(DP_mult_210_n529), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n530), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n327) );
  XNOR2_X1 DP_mult_210_U338 ( .A(DP_b_int_1__1_), .B(DP_mult_210_n513), .ZN(
        DP_mult_210_n528) );
  OAI22_X1 DP_mult_210_U337 ( .A1(DP_mult_210_n528), .A2(DP_mult_210_n527), 
        .B1(DP_mult_210_n529), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n328) );
  OAI22_X1 DP_mult_210_U336 ( .A1(DP_b_int_1__0_), .A2(DP_mult_210_n527), .B1(
        DP_mult_210_n528), .B2(DP_mult_210_n526), .ZN(DP_mult_210_n329) );
  NOR2_X1 DP_mult_210_U335 ( .A1(DP_mult_210_n525), .A2(DP_mult_210_n526), 
        .ZN(DP_coeff_pipe02[0]) );
  INV_X1 DP_mult_210_U334 ( .A(DP_mult_210_n120), .ZN(DP_N121) );
  INV_X1 DP_mult_210_U333 ( .A(DP_a_int_1__1_), .ZN(DP_mult_210_n514) );
  XOR2_X2 DP_mult_210_U332 ( .A(DP_a_int_1__10_), .B(DP_mult_210_n522), .Z(
        DP_mult_210_n600) );
  XOR2_X2 DP_mult_210_U331 ( .A(DP_a_int_1__8_), .B(DP_mult_210_n520), .Z(
        DP_mult_210_n585) );
  XOR2_X2 DP_mult_210_U330 ( .A(DP_a_int_1__6_), .B(DP_mult_210_n518), .Z(
        DP_mult_210_n570) );
  XOR2_X2 DP_mult_210_U329 ( .A(DP_a_int_1__4_), .B(DP_mult_210_n516), .Z(
        DP_mult_210_n555) );
  XOR2_X2 DP_mult_210_U328 ( .A(DP_a_int_1__2_), .B(DP_mult_210_n514), .Z(
        DP_mult_210_n540) );
  INV_X1 DP_mult_210_U327 ( .A(DP_a_int_1__5_), .ZN(DP_mult_210_n518) );
  INV_X1 DP_mult_210_U326 ( .A(DP_a_int_1__3_), .ZN(DP_mult_210_n516) );
  INV_X1 DP_mult_210_U325 ( .A(DP_a_int_1__9_), .ZN(DP_mult_210_n522) );
  INV_X1 DP_mult_210_U324 ( .A(DP_a_int_1__7_), .ZN(DP_mult_210_n520) );
  INV_X1 DP_mult_210_U323 ( .A(DP_a_int_1__11_), .ZN(DP_mult_210_n524) );
  INV_X1 DP_mult_210_U322 ( .A(DP_mult_210_n514), .ZN(DP_mult_210_n513) );
  INV_X1 DP_mult_210_U321 ( .A(DP_mult_210_n522), .ZN(DP_mult_210_n521) );
  INV_X1 DP_mult_210_U320 ( .A(DP_mult_210_n520), .ZN(DP_mult_210_n519) );
  INV_X1 DP_mult_210_U319 ( .A(DP_mult_210_n518), .ZN(DP_mult_210_n517) );
  INV_X1 DP_mult_210_U318 ( .A(DP_mult_210_n516), .ZN(DP_mult_210_n515) );
  INV_X1 DP_mult_210_U317 ( .A(DP_mult_210_n524), .ZN(DP_mult_210_n523) );
  HA_X1 DP_mult_210_U107 ( .A(DP_mult_210_n316), .B(DP_mult_210_n327), .CO(
        DP_mult_210_n250), .S(DP_mult_210_n251) );
  FA_X1 DP_mult_210_U106 ( .A(DP_mult_210_n326), .B(DP_mult_210_n305), .CI(
        DP_mult_210_n315), .CO(DP_mult_210_n248), .S(DP_mult_210_n249) );
  HA_X1 DP_mult_210_U105 ( .A(DP_mult_210_n255), .B(DP_mult_210_n304), .CO(
        DP_mult_210_n246), .S(DP_mult_210_n247) );
  FA_X1 DP_mult_210_U104 ( .A(DP_mult_210_n314), .B(DP_mult_210_n325), .CI(
        DP_mult_210_n247), .CO(DP_mult_210_n244), .S(DP_mult_210_n245) );
  FA_X1 DP_mult_210_U103 ( .A(DP_mult_210_n324), .B(DP_mult_210_n293), .CI(
        DP_mult_210_n313), .CO(DP_mult_210_n242), .S(DP_mult_210_n243) );
  FA_X1 DP_mult_210_U102 ( .A(DP_mult_210_n246), .B(DP_mult_210_n303), .CI(
        DP_mult_210_n243), .CO(DP_mult_210_n240), .S(DP_mult_210_n241) );
  HA_X1 DP_mult_210_U101 ( .A(DP_mult_210_n254), .B(DP_mult_210_n292), .CO(
        DP_mult_210_n238), .S(DP_mult_210_n239) );
  FA_X1 DP_mult_210_U100 ( .A(DP_mult_210_n302), .B(DP_mult_210_n323), .CI(
        DP_mult_210_n312), .CO(DP_mult_210_n236), .S(DP_mult_210_n237) );
  FA_X1 DP_mult_210_U99 ( .A(DP_mult_210_n242), .B(DP_mult_210_n239), .CI(
        DP_mult_210_n237), .CO(DP_mult_210_n234), .S(DP_mult_210_n235) );
  FA_X1 DP_mult_210_U98 ( .A(DP_mult_210_n301), .B(DP_mult_210_n281), .CI(
        DP_mult_210_n322), .CO(DP_mult_210_n232), .S(DP_mult_210_n233) );
  FA_X1 DP_mult_210_U97 ( .A(DP_mult_210_n291), .B(DP_mult_210_n311), .CI(
        DP_mult_210_n238), .CO(DP_mult_210_n230), .S(DP_mult_210_n231) );
  FA_X1 DP_mult_210_U96 ( .A(DP_mult_210_n233), .B(DP_mult_210_n236), .CI(
        DP_mult_210_n231), .CO(DP_mult_210_n228), .S(DP_mult_210_n229) );
  HA_X1 DP_mult_210_U95 ( .A(DP_mult_210_n253), .B(DP_mult_210_n280), .CO(
        DP_mult_210_n226), .S(DP_mult_210_n227) );
  FA_X1 DP_mult_210_U94 ( .A(DP_mult_210_n290), .B(DP_mult_210_n300), .CI(
        DP_mult_210_n310), .CO(DP_mult_210_n224), .S(DP_mult_210_n225) );
  FA_X1 DP_mult_210_U93 ( .A(DP_mult_210_n227), .B(DP_mult_210_n321), .CI(
        DP_mult_210_n232), .CO(DP_mult_210_n222), .S(DP_mult_210_n223) );
  FA_X1 DP_mult_210_U92 ( .A(DP_mult_210_n225), .B(DP_mult_210_n230), .CI(
        DP_mult_210_n223), .CO(DP_mult_210_n220), .S(DP_mult_210_n221) );
  FA_X1 DP_mult_210_U91 ( .A(DP_mult_210_n289), .B(DP_mult_210_n269), .CI(
        DP_mult_210_n320), .CO(DP_mult_210_n218), .S(DP_mult_210_n219) );
  FA_X1 DP_mult_210_U90 ( .A(DP_mult_210_n279), .B(DP_mult_210_n309), .CI(
        DP_mult_210_n299), .CO(DP_mult_210_n216), .S(DP_mult_210_n217) );
  FA_X1 DP_mult_210_U89 ( .A(DP_mult_210_n224), .B(DP_mult_210_n226), .CI(
        DP_mult_210_n219), .CO(DP_mult_210_n214), .S(DP_mult_210_n215) );
  FA_X1 DP_mult_210_U88 ( .A(DP_mult_210_n222), .B(DP_mult_210_n217), .CI(
        DP_mult_210_n215), .CO(DP_mult_210_n212), .S(DP_mult_210_n213) );
  HA_X1 DP_mult_210_U87 ( .A(DP_mult_210_n252), .B(DP_mult_210_n268), .CO(
        DP_mult_210_n210), .S(DP_mult_210_n211) );
  FA_X1 DP_mult_210_U86 ( .A(DP_mult_210_n278), .B(DP_mult_210_n298), .CI(
        DP_mult_210_n319), .CO(DP_mult_210_n208), .S(DP_mult_210_n209) );
  FA_X1 DP_mult_210_U85 ( .A(DP_mult_210_n288), .B(DP_mult_210_n308), .CI(
        DP_mult_210_n211), .CO(DP_mult_210_n206), .S(DP_mult_210_n207) );
  FA_X1 DP_mult_210_U84 ( .A(DP_mult_210_n216), .B(DP_mult_210_n218), .CI(
        DP_mult_210_n209), .CO(DP_mult_210_n204), .S(DP_mult_210_n205) );
  FA_X1 DP_mult_210_U83 ( .A(DP_mult_210_n214), .B(DP_mult_210_n207), .CI(
        DP_mult_210_n205), .CO(DP_mult_210_n202), .S(DP_mult_210_n203) );
  FA_X1 DP_mult_210_U80 ( .A(DP_mult_210_n267), .B(DP_mult_210_n287), .CI(
        DP_mult_210_n318), .CO(DP_mult_210_n198), .S(DP_mult_210_n199) );
  FA_X1 DP_mult_210_U79 ( .A(DP_mult_210_n210), .B(DP_mult_210_n307), .CI(
        DP_mult_210_n201), .CO(DP_mult_210_n196), .S(DP_mult_210_n197) );
  FA_X1 DP_mult_210_U78 ( .A(DP_mult_210_n199), .B(DP_mult_210_n208), .CI(
        DP_mult_210_n206), .CO(DP_mult_210_n194), .S(DP_mult_210_n195) );
  FA_X1 DP_mult_210_U77 ( .A(DP_mult_210_n204), .B(DP_mult_210_n197), .CI(
        DP_mult_210_n195), .CO(DP_mult_210_n192), .S(DP_mult_210_n193) );
  FA_X1 DP_mult_210_U75 ( .A(DP_mult_210_n296), .B(DP_mult_210_n276), .CI(
        DP_mult_210_n191), .CO(DP_mult_210_n188), .S(DP_mult_210_n189) );
  FA_X1 DP_mult_210_U74 ( .A(DP_mult_210_n266), .B(DP_mult_210_n286), .CI(
        DP_mult_210_n200), .CO(DP_mult_210_n186), .S(DP_mult_210_n187) );
  FA_X1 DP_mult_210_U73 ( .A(DP_mult_210_n196), .B(DP_mult_210_n198), .CI(
        DP_mult_210_n189), .CO(DP_mult_210_n184), .S(DP_mult_210_n185) );
  FA_X1 DP_mult_210_U72 ( .A(DP_mult_210_n194), .B(DP_mult_210_n187), .CI(
        DP_mult_210_n185), .CO(DP_mult_210_n182), .S(DP_mult_210_n183) );
  FA_X1 DP_mult_210_U71 ( .A(DP_mult_210_n190), .B(DP_mult_210_n265), .CI(
        DP_mult_210_n306), .CO(DP_mult_210_n180), .S(DP_mult_210_n181) );
  FA_X1 DP_mult_210_U70 ( .A(DP_mult_210_n275), .B(DP_mult_210_n295), .CI(
        DP_mult_210_n285), .CO(DP_mult_210_n178), .S(DP_mult_210_n179) );
  FA_X1 DP_mult_210_U69 ( .A(DP_mult_210_n186), .B(DP_mult_210_n188), .CI(
        DP_mult_210_n179), .CO(DP_mult_210_n176), .S(DP_mult_210_n177) );
  FA_X1 DP_mult_210_U68 ( .A(DP_mult_210_n184), .B(DP_mult_210_n181), .CI(
        DP_mult_210_n177), .CO(DP_mult_210_n174), .S(DP_mult_210_n175) );
  FA_X1 DP_mult_210_U66 ( .A(DP_mult_210_n264), .B(DP_mult_210_n274), .CI(
        DP_mult_210_n173), .CO(DP_mult_210_n170), .S(DP_mult_210_n171) );
  FA_X1 DP_mult_210_U65 ( .A(DP_mult_210_n180), .B(DP_mult_210_n284), .CI(
        DP_mult_210_n178), .CO(DP_mult_210_n168), .S(DP_mult_210_n169) );
  FA_X1 DP_mult_210_U64 ( .A(DP_mult_210_n176), .B(DP_mult_210_n171), .CI(
        DP_mult_210_n169), .CO(DP_mult_210_n166), .S(DP_mult_210_n167) );
  FA_X1 DP_mult_210_U63 ( .A(DP_mult_210_n172), .B(DP_mult_210_n263), .CI(
        DP_mult_210_n294), .CO(DP_mult_210_n164), .S(DP_mult_210_n165) );
  FA_X1 DP_mult_210_U62 ( .A(DP_mult_210_n273), .B(DP_mult_210_n283), .CI(
        DP_mult_210_n170), .CO(DP_mult_210_n162), .S(DP_mult_210_n163) );
  FA_X1 DP_mult_210_U61 ( .A(DP_mult_210_n168), .B(DP_mult_210_n165), .CI(
        DP_mult_210_n163), .CO(DP_mult_210_n160), .S(DP_mult_210_n161) );
  FA_X1 DP_mult_210_U59 ( .A(DP_mult_210_n262), .B(DP_mult_210_n272), .CI(
        DP_mult_210_n159), .CO(DP_mult_210_n156), .S(DP_mult_210_n157) );
  FA_X1 DP_mult_210_U58 ( .A(DP_mult_210_n157), .B(DP_mult_210_n164), .CI(
        DP_mult_210_n162), .CO(DP_mult_210_n154), .S(DP_mult_210_n155) );
  FA_X1 DP_mult_210_U57 ( .A(DP_mult_210_n261), .B(DP_mult_210_n158), .CI(
        DP_mult_210_n282), .CO(DP_mult_210_n152), .S(DP_mult_210_n153) );
  FA_X1 DP_mult_210_U56 ( .A(DP_mult_210_n156), .B(DP_mult_210_n271), .CI(
        DP_mult_210_n153), .CO(DP_mult_210_n150), .S(DP_mult_210_n151) );
  FA_X1 DP_mult_210_U54 ( .A(DP_mult_210_n149), .B(DP_mult_210_n260), .CI(
        DP_mult_210_n152), .CO(DP_mult_210_n146), .S(DP_mult_210_n147) );
  FA_X1 DP_mult_210_U53 ( .A(DP_mult_210_n259), .B(DP_mult_210_n148), .CI(
        DP_mult_210_n270), .CO(DP_mult_210_n144), .S(DP_mult_210_n145) );
  HA_X1 DP_mult_210_U51 ( .A(DP_mult_210_n329), .B(DP_mult_210_n257), .CO(
        DP_mult_210_n141), .S(DP_N99) );
  FA_X1 DP_mult_210_U50 ( .A(DP_mult_210_n328), .B(DP_mult_210_n317), .CI(
        DP_mult_210_n141), .CO(DP_mult_210_n140), .S(DP_N100) );
  FA_X1 DP_mult_210_U49 ( .A(DP_mult_210_n251), .B(DP_mult_210_n256), .CI(
        DP_mult_210_n140), .CO(DP_mult_210_n139), .S(DP_N101) );
  FA_X1 DP_mult_210_U48 ( .A(DP_mult_210_n249), .B(DP_mult_210_n250), .CI(
        DP_mult_210_n139), .CO(DP_mult_210_n138), .S(DP_N102) );
  FA_X1 DP_mult_210_U47 ( .A(DP_mult_210_n245), .B(DP_mult_210_n248), .CI(
        DP_mult_210_n138), .CO(DP_mult_210_n137), .S(DP_N103) );
  FA_X1 DP_mult_210_U46 ( .A(DP_mult_210_n241), .B(DP_mult_210_n244), .CI(
        DP_mult_210_n137), .CO(DP_mult_210_n136), .S(DP_N104) );
  FA_X1 DP_mult_210_U45 ( .A(DP_mult_210_n235), .B(DP_mult_210_n240), .CI(
        DP_mult_210_n136), .CO(DP_mult_210_n135), .S(DP_N105) );
  FA_X1 DP_mult_210_U44 ( .A(DP_mult_210_n229), .B(DP_mult_210_n234), .CI(
        DP_mult_210_n135), .CO(DP_mult_210_n134), .S(DP_N106) );
  FA_X1 DP_mult_210_U43 ( .A(DP_mult_210_n221), .B(DP_mult_210_n228), .CI(
        DP_mult_210_n134), .CO(DP_mult_210_n133), .S(DP_N107) );
  FA_X1 DP_mult_210_U42 ( .A(DP_mult_210_n213), .B(DP_mult_210_n220), .CI(
        DP_mult_210_n133), .CO(DP_mult_210_n132), .S(DP_N108) );
  FA_X1 DP_mult_210_U41 ( .A(DP_mult_210_n203), .B(DP_mult_210_n212), .CI(
        DP_mult_210_n132), .CO(DP_mult_210_n131), .S(DP_N109) );
  FA_X1 DP_mult_210_U40 ( .A(DP_mult_210_n193), .B(DP_mult_210_n202), .CI(
        DP_mult_210_n131), .CO(DP_mult_210_n130), .S(DP_N110) );
  FA_X1 DP_mult_210_U39 ( .A(DP_mult_210_n183), .B(DP_mult_210_n192), .CI(
        DP_mult_210_n130), .CO(DP_mult_210_n129), .S(DP_N111) );
  FA_X1 DP_mult_210_U38 ( .A(DP_mult_210_n175), .B(DP_mult_210_n182), .CI(
        DP_mult_210_n129), .CO(DP_mult_210_n128), .S(DP_N112) );
  FA_X1 DP_mult_210_U37 ( .A(DP_mult_210_n167), .B(DP_mult_210_n174), .CI(
        DP_mult_210_n128), .CO(DP_mult_210_n127), .S(DP_N113) );
  FA_X1 DP_mult_210_U36 ( .A(DP_mult_210_n161), .B(DP_mult_210_n166), .CI(
        DP_mult_210_n127), .CO(DP_mult_210_n126), .S(DP_N114) );
  FA_X1 DP_mult_210_U30 ( .A(DP_mult_210_n160), .B(DP_mult_210_n155), .CI(
        DP_mult_210_n126), .CO(DP_mult_210_n125), .S(DP_N115) );
  FA_X1 DP_mult_210_U20 ( .A(DP_mult_210_n151), .B(DP_mult_210_n154), .CI(
        DP_mult_210_n125), .CO(DP_mult_210_n124), .S(DP_N116) );
  FA_X1 DP_mult_210_U10 ( .A(DP_mult_210_n147), .B(DP_mult_210_n150), .CI(
        DP_mult_210_n124), .CO(DP_mult_210_n123), .S(DP_N117) );
  FA_X1 DP_mult_210_U9 ( .A(DP_mult_210_n146), .B(DP_mult_210_n145), .CI(
        DP_mult_210_n123), .CO(DP_mult_210_n122), .S(DP_N118) );
  FA_X1 DP_mult_210_U8 ( .A(DP_mult_210_n144), .B(DP_mult_210_n143), .CI(
        DP_mult_210_n122), .CO(DP_mult_210_n121), .S(DP_N119) );
  FA_X1 DP_mult_210_U7 ( .A(DP_mult_210_n258), .B(DP_mult_210_n142), .CI(
        DP_mult_210_n121), .CO(DP_mult_210_n120), .S(DP_N120) );
  INV_X1 DP_sub_210_U44 ( .A(DP_N108), .ZN(DP_sub_210_B_not_10_) );
  INV_X1 DP_sub_210_U43 ( .A(DP_N109), .ZN(DP_sub_210_B_not_11_) );
  INV_X1 DP_sub_210_U42 ( .A(DP_N110), .ZN(DP_sub_210_B_not_12_) );
  INV_X1 DP_sub_210_U41 ( .A(DP_N111), .ZN(DP_sub_210_B_not_13_) );
  INV_X1 DP_sub_210_U40 ( .A(DP_N112), .ZN(DP_sub_210_B_not_14_) );
  INV_X1 DP_sub_210_U39 ( .A(DP_N113), .ZN(DP_sub_210_B_not_15_) );
  INV_X1 DP_sub_210_U38 ( .A(DP_N114), .ZN(DP_sub_210_B_not_16_) );
  INV_X1 DP_sub_210_U37 ( .A(DP_N115), .ZN(DP_sub_210_B_not_17_) );
  INV_X1 DP_sub_210_U36 ( .A(DP_N116), .ZN(DP_sub_210_B_not_18_) );
  INV_X1 DP_sub_210_U35 ( .A(DP_N117), .ZN(DP_sub_210_B_not_19_) );
  INV_X1 DP_sub_210_U34 ( .A(DP_N99), .ZN(DP_sub_210_B_not_1_) );
  INV_X1 DP_sub_210_U33 ( .A(DP_N118), .ZN(DP_sub_210_B_not_20_) );
  INV_X1 DP_sub_210_U32 ( .A(DP_N119), .ZN(DP_sub_210_B_not_21_) );
  INV_X1 DP_sub_210_U31 ( .A(DP_N120), .ZN(DP_sub_210_B_not_22_) );
  INV_X1 DP_sub_210_U30 ( .A(DP_N121), .ZN(DP_sub_210_B_not_23_) );
  INV_X1 DP_sub_210_U29 ( .A(DP_N100), .ZN(DP_sub_210_B_not_2_) );
  INV_X1 DP_sub_210_U28 ( .A(DP_N101), .ZN(DP_sub_210_B_not_3_) );
  INV_X1 DP_sub_210_U27 ( .A(DP_N102), .ZN(DP_sub_210_B_not_4_) );
  INV_X1 DP_sub_210_U26 ( .A(DP_N103), .ZN(DP_sub_210_B_not_5_) );
  INV_X1 DP_sub_210_U25 ( .A(DP_N104), .ZN(DP_sub_210_B_not_6_) );
  INV_X1 DP_sub_210_U24 ( .A(DP_N105), .ZN(DP_sub_210_B_not_7_) );
  INV_X1 DP_sub_210_U23 ( .A(DP_N106), .ZN(DP_sub_210_B_not_8_) );
  INV_X1 DP_sub_210_U22 ( .A(DP_N107), .ZN(DP_sub_210_B_not_9_) );
  INV_X1 DP_sub_210_U21 ( .A(DP_coeff_pipe02[0]), .ZN(DP_sub_210_carry_1_) );
  XOR2_X1 DP_sub_210_U20 ( .A(DP_sub_210_B_not_1_), .B(DP_sub_210_carry_1_), 
        .Z(DP_coeff_pipe02[1]) );
  AND2_X1 DP_sub_210_U19 ( .A1(DP_sub_210_carry_1_), .A2(DP_sub_210_B_not_1_), 
        .ZN(DP_sub_210_carry_2_) );
  AND2_X1 DP_sub_210_U18 ( .A1(DP_sub_210_carry_2_), .A2(DP_sub_210_B_not_2_), 
        .ZN(DP_sub_210_carry_3_) );
  XOR2_X1 DP_sub_210_U17 ( .A(DP_sub_210_B_not_3_), .B(DP_sub_210_carry_3_), 
        .Z(DP_coeff_pipe02[3]) );
  AND2_X1 DP_sub_210_U16 ( .A1(DP_sub_210_carry_3_), .A2(DP_sub_210_B_not_3_), 
        .ZN(DP_sub_210_carry_4_) );
  XOR2_X1 DP_sub_210_U15 ( .A(DP_sub_210_B_not_4_), .B(DP_sub_210_carry_4_), 
        .Z(DP_coeff_pipe02[4]) );
  AND2_X1 DP_sub_210_U14 ( .A1(DP_sub_210_carry_4_), .A2(DP_sub_210_B_not_4_), 
        .ZN(DP_sub_210_carry_5_) );
  XOR2_X1 DP_sub_210_U13 ( .A(DP_sub_210_B_not_5_), .B(DP_sub_210_carry_5_), 
        .Z(DP_coeff_pipe02[5]) );
  AND2_X1 DP_sub_210_U12 ( .A1(DP_sub_210_carry_5_), .A2(DP_sub_210_B_not_5_), 
        .ZN(DP_sub_210_carry_6_) );
  XOR2_X1 DP_sub_210_U11 ( .A(DP_sub_210_B_not_6_), .B(DP_sub_210_carry_6_), 
        .Z(DP_coeff_pipe02[6]) );
  AND2_X1 DP_sub_210_U10 ( .A1(DP_sub_210_carry_6_), .A2(DP_sub_210_B_not_6_), 
        .ZN(DP_sub_210_carry_7_) );
  XOR2_X1 DP_sub_210_U9 ( .A(DP_sub_210_B_not_7_), .B(DP_sub_210_carry_7_), 
        .Z(DP_coeff_pipe02[7]) );
  AND2_X1 DP_sub_210_U8 ( .A1(DP_sub_210_carry_7_), .A2(DP_sub_210_B_not_7_), 
        .ZN(DP_sub_210_carry_8_) );
  XOR2_X1 DP_sub_210_U7 ( .A(DP_sub_210_B_not_8_), .B(DP_sub_210_carry_8_), 
        .Z(DP_coeff_pipe02[8]) );
  AND2_X1 DP_sub_210_U6 ( .A1(DP_sub_210_carry_8_), .A2(DP_sub_210_B_not_8_), 
        .ZN(DP_sub_210_carry_9_) );
  XOR2_X1 DP_sub_210_U5 ( .A(DP_sub_210_B_not_9_), .B(DP_sub_210_carry_9_), 
        .Z(DP_coeff_pipe02[9]) );
  AND2_X1 DP_sub_210_U4 ( .A1(DP_sub_210_carry_9_), .A2(DP_sub_210_B_not_9_), 
        .ZN(DP_sub_210_carry_10_) );
  XOR2_X1 DP_sub_210_U3 ( .A(DP_sub_210_B_not_10_), .B(DP_sub_210_carry_10_), 
        .Z(DP_coeff_pipe02[10]) );
  AND2_X1 DP_sub_210_U2 ( .A1(DP_sub_210_carry_10_), .A2(DP_sub_210_B_not_10_), 
        .ZN(DP_sub_210_carry_11_) );
  XOR2_X2 DP_sub_210_U1 ( .A(DP_sub_210_B_not_2_), .B(DP_sub_210_carry_2_), 
        .Z(DP_coeff_pipe02[2]) );
  FA_X1 DP_sub_210_U2_11 ( .A(DP_b_int_2__0_), .B(DP_sub_210_B_not_11_), .CI(
        DP_sub_210_carry_11_), .CO(DP_sub_210_carry_12_), .S(
        DP_coeff_pipe02[11]) );
  FA_X1 DP_sub_210_U2_12 ( .A(DP_b_int_2__1_), .B(DP_sub_210_B_not_12_), .CI(
        DP_sub_210_carry_12_), .CO(DP_sub_210_carry_13_), .S(
        DP_coeff_pipe02[12]) );
  FA_X1 DP_sub_210_U2_13 ( .A(DP_b_int_2__2_), .B(DP_sub_210_B_not_13_), .CI(
        DP_sub_210_carry_13_), .CO(DP_sub_210_carry_14_), .S(
        DP_coeff_pipe02[13]) );
  FA_X1 DP_sub_210_U2_14 ( .A(DP_b_int_2__3_), .B(DP_sub_210_B_not_14_), .CI(
        DP_sub_210_carry_14_), .CO(DP_sub_210_carry_15_), .S(
        DP_coeff_pipe02[14]) );
  FA_X1 DP_sub_210_U2_15 ( .A(DP_b_int_2__4_), .B(DP_sub_210_B_not_15_), .CI(
        DP_sub_210_carry_15_), .CO(DP_sub_210_carry_16_), .S(
        DP_coeff_pipe02[15]) );
  FA_X1 DP_sub_210_U2_16 ( .A(DP_b_int_2__5_), .B(DP_sub_210_B_not_16_), .CI(
        DP_sub_210_carry_16_), .CO(DP_sub_210_carry_17_), .S(
        DP_coeff_pipe02[16]) );
  FA_X1 DP_sub_210_U2_17 ( .A(DP_b_int_2__6_), .B(DP_sub_210_B_not_17_), .CI(
        DP_sub_210_carry_17_), .CO(DP_sub_210_carry_18_), .S(
        DP_coeff_pipe02[17]) );
  FA_X1 DP_sub_210_U2_18 ( .A(DP_b_int_2__7_), .B(DP_sub_210_B_not_18_), .CI(
        DP_sub_210_carry_18_), .CO(DP_sub_210_carry_19_), .S(
        DP_coeff_pipe02[18]) );
  FA_X1 DP_sub_210_U2_19 ( .A(DP_b_int_2__8_), .B(DP_sub_210_B_not_19_), .CI(
        DP_sub_210_carry_19_), .CO(DP_sub_210_carry_20_), .S(
        DP_coeff_pipe02[19]) );
  FA_X1 DP_sub_210_U2_20 ( .A(DP_b_int_2__9_), .B(DP_sub_210_B_not_20_), .CI(
        DP_sub_210_carry_20_), .CO(DP_sub_210_carry_21_), .S(
        DP_coeff_pipe02[20]) );
  FA_X1 DP_sub_210_U2_21 ( .A(DP_b_int_2__10_), .B(DP_sub_210_B_not_21_), .CI(
        DP_sub_210_carry_21_), .CO(DP_sub_210_carry_22_), .S(
        DP_coeff_pipe02[21]) );
  FA_X1 DP_sub_210_U2_22 ( .A(DP_b_int_2__11_), .B(DP_sub_210_B_not_22_), .CI(
        DP_sub_210_carry_22_), .CO(DP_sub_210_carry_23_), .S(
        DP_coeff_pipe02[22]) );
  FA_X1 DP_sub_210_U2_23 ( .A(DP_b_int_2__11_), .B(DP_sub_210_B_not_23_), .CI(
        DP_sub_210_carry_23_), .S(DP_coeff_pipe02[23]) );
  XNOR2_X1 DP_mult_211_U515 ( .A(DP_b_int_2__10_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n607) );
  XNOR2_X1 DP_mult_211_U514 ( .A(DP_mult_211_n519), .B(DP_a_int_1__10_), .ZN(
        DP_mult_211_n621) );
  NAND2_X1 DP_mult_211_U513 ( .A1(DP_mult_211_n595), .A2(DP_mult_211_n621), 
        .ZN(DP_mult_211_n597) );
  XNOR2_X1 DP_mult_211_U512 ( .A(DP_b_int_2__11_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n609) );
  OAI22_X1 DP_mult_211_U511 ( .A1(DP_mult_211_n607), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n609), .ZN(DP_mult_211_n142) );
  INV_X1 DP_mult_211_U510 ( .A(DP_mult_211_n142), .ZN(DP_mult_211_n143) );
  XNOR2_X1 DP_mult_211_U509 ( .A(DP_b_int_2__10_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n592) );
  XNOR2_X1 DP_mult_211_U508 ( .A(DP_mult_211_n517), .B(DP_a_int_1__8_), .ZN(
        DP_mult_211_n620) );
  NAND2_X1 DP_mult_211_U507 ( .A1(DP_mult_211_n580), .A2(DP_mult_211_n620), 
        .ZN(DP_mult_211_n582) );
  XNOR2_X1 DP_mult_211_U506 ( .A(DP_b_int_2__11_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n594) );
  OAI22_X1 DP_mult_211_U505 ( .A1(DP_mult_211_n592), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n594), .ZN(DP_mult_211_n148) );
  INV_X1 DP_mult_211_U504 ( .A(DP_mult_211_n148), .ZN(DP_mult_211_n149) );
  XNOR2_X1 DP_mult_211_U503 ( .A(DP_b_int_2__10_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n577) );
  XNOR2_X1 DP_mult_211_U502 ( .A(DP_mult_211_n516), .B(DP_a_int_1__6_), .ZN(
        DP_mult_211_n619) );
  NAND2_X1 DP_mult_211_U501 ( .A1(DP_mult_211_n565), .A2(DP_mult_211_n619), 
        .ZN(DP_mult_211_n567) );
  XNOR2_X1 DP_mult_211_U500 ( .A(DP_b_int_2__11_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n579) );
  OAI22_X1 DP_mult_211_U499 ( .A1(DP_mult_211_n577), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n579), .ZN(DP_mult_211_n158) );
  INV_X1 DP_mult_211_U498 ( .A(DP_mult_211_n158), .ZN(DP_mult_211_n159) );
  XNOR2_X1 DP_mult_211_U497 ( .A(DP_b_int_2__10_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n562) );
  XNOR2_X1 DP_mult_211_U496 ( .A(DP_mult_211_n515), .B(DP_a_int_1__4_), .ZN(
        DP_mult_211_n618) );
  NAND2_X1 DP_mult_211_U495 ( .A1(DP_mult_211_n550), .A2(DP_mult_211_n618), 
        .ZN(DP_mult_211_n552) );
  XNOR2_X1 DP_mult_211_U494 ( .A(DP_b_int_2__11_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n564) );
  OAI22_X1 DP_mult_211_U493 ( .A1(DP_mult_211_n562), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n564), .ZN(DP_mult_211_n172) );
  INV_X1 DP_mult_211_U492 ( .A(DP_mult_211_n172), .ZN(DP_mult_211_n173) );
  XNOR2_X1 DP_mult_211_U491 ( .A(DP_b_int_2__10_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n547) );
  XNOR2_X1 DP_mult_211_U490 ( .A(DP_mult_211_n514), .B(DP_a_int_1__2_), .ZN(
        DP_mult_211_n617) );
  NAND2_X1 DP_mult_211_U489 ( .A1(DP_mult_211_n535), .A2(DP_mult_211_n617), 
        .ZN(DP_mult_211_n537) );
  XNOR2_X1 DP_mult_211_U488 ( .A(DP_b_int_2__11_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n549) );
  OAI22_X1 DP_mult_211_U487 ( .A1(DP_mult_211_n547), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n549), .ZN(DP_mult_211_n190) );
  INV_X1 DP_mult_211_U486 ( .A(DP_mult_211_n190), .ZN(DP_mult_211_n191) );
  XNOR2_X1 DP_mult_211_U485 ( .A(DP_b_int_2__3_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n585) );
  XNOR2_X1 DP_mult_211_U484 ( .A(DP_b_int_2__4_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n586) );
  OAI22_X1 DP_mult_211_U483 ( .A1(DP_mult_211_n585), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n586), .ZN(DP_mult_211_n615) );
  XNOR2_X1 DP_mult_211_U482 ( .A(DP_b_int_2__7_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n559) );
  XNOR2_X1 DP_mult_211_U481 ( .A(DP_b_int_2__8_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n560) );
  OAI22_X1 DP_mult_211_U480 ( .A1(DP_mult_211_n559), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n560), .ZN(DP_mult_211_n616) );
  OR2_X1 DP_mult_211_U479 ( .A1(DP_mult_211_n615), .A2(DP_mult_211_n616), .ZN(
        DP_mult_211_n200) );
  XNOR2_X1 DP_mult_211_U478 ( .A(DP_mult_211_n615), .B(DP_mult_211_n616), .ZN(
        DP_mult_211_n201) );
  OR3_X1 DP_mult_211_U477 ( .A1(DP_mult_211_n595), .A2(DP_b_int_2__0_), .A3(
        DP_mult_211_n519), .ZN(DP_mult_211_n614) );
  OAI21_X1 DP_mult_211_U476 ( .B1(DP_mult_211_n519), .B2(DP_mult_211_n597), 
        .A(DP_mult_211_n614), .ZN(DP_mult_211_n252) );
  OR3_X1 DP_mult_211_U475 ( .A1(DP_mult_211_n580), .A2(DP_b_int_2__0_), .A3(
        DP_mult_211_n517), .ZN(DP_mult_211_n613) );
  OAI21_X1 DP_mult_211_U474 ( .B1(DP_mult_211_n517), .B2(DP_mult_211_n582), 
        .A(DP_mult_211_n613), .ZN(DP_mult_211_n253) );
  OR3_X1 DP_mult_211_U473 ( .A1(DP_mult_211_n565), .A2(DP_b_int_2__0_), .A3(
        DP_mult_211_n516), .ZN(DP_mult_211_n612) );
  OAI21_X1 DP_mult_211_U472 ( .B1(DP_mult_211_n516), .B2(DP_mult_211_n567), 
        .A(DP_mult_211_n612), .ZN(DP_mult_211_n254) );
  OR3_X1 DP_mult_211_U471 ( .A1(DP_mult_211_n550), .A2(DP_b_int_2__0_), .A3(
        DP_mult_211_n515), .ZN(DP_mult_211_n611) );
  OAI21_X1 DP_mult_211_U470 ( .B1(DP_mult_211_n515), .B2(DP_mult_211_n552), 
        .A(DP_mult_211_n611), .ZN(DP_mult_211_n255) );
  OR3_X1 DP_mult_211_U469 ( .A1(DP_mult_211_n535), .A2(DP_b_int_2__0_), .A3(
        DP_mult_211_n514), .ZN(DP_mult_211_n610) );
  OAI21_X1 DP_mult_211_U468 ( .B1(DP_mult_211_n514), .B2(DP_mult_211_n537), 
        .A(DP_mult_211_n610), .ZN(DP_mult_211_n256) );
  NAND2_X1 DP_mult_211_U467 ( .A1(DP_a_int_1__1_), .A2(DP_mult_211_n521), .ZN(
        DP_mult_211_n522) );
  OAI21_X1 DP_mult_211_U466 ( .B1(DP_b_int_2__0_), .B2(DP_mult_211_n513), .A(
        DP_mult_211_n522), .ZN(DP_mult_211_n257) );
  AOI21_X1 DP_mult_211_U465 ( .B1(DP_mult_211_n597), .B2(DP_mult_211_n595), 
        .A(DP_mult_211_n609), .ZN(DP_mult_211_n608) );
  INV_X1 DP_mult_211_U464 ( .A(DP_mult_211_n608), .ZN(DP_mult_211_n258) );
  XNOR2_X1 DP_mult_211_U463 ( .A(DP_b_int_2__9_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n606) );
  OAI22_X1 DP_mult_211_U462 ( .A1(DP_mult_211_n606), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n607), .ZN(DP_mult_211_n259) );
  XNOR2_X1 DP_mult_211_U461 ( .A(DP_b_int_2__8_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n605) );
  OAI22_X1 DP_mult_211_U460 ( .A1(DP_mult_211_n605), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n606), .ZN(DP_mult_211_n260) );
  XNOR2_X1 DP_mult_211_U459 ( .A(DP_b_int_2__7_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n604) );
  OAI22_X1 DP_mult_211_U458 ( .A1(DP_mult_211_n604), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n605), .ZN(DP_mult_211_n261) );
  XNOR2_X1 DP_mult_211_U457 ( .A(DP_b_int_2__6_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n603) );
  OAI22_X1 DP_mult_211_U456 ( .A1(DP_mult_211_n603), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n604), .ZN(DP_mult_211_n262) );
  XNOR2_X1 DP_mult_211_U455 ( .A(DP_b_int_2__5_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n602) );
  OAI22_X1 DP_mult_211_U454 ( .A1(DP_mult_211_n602), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n603), .ZN(DP_mult_211_n263) );
  XNOR2_X1 DP_mult_211_U453 ( .A(DP_b_int_2__4_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n601) );
  OAI22_X1 DP_mult_211_U452 ( .A1(DP_mult_211_n601), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n602), .ZN(DP_mult_211_n264) );
  XNOR2_X1 DP_mult_211_U451 ( .A(DP_b_int_2__3_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n600) );
  OAI22_X1 DP_mult_211_U450 ( .A1(DP_mult_211_n600), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n601), .ZN(DP_mult_211_n265) );
  XNOR2_X1 DP_mult_211_U449 ( .A(DP_b_int_2__2_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n599) );
  OAI22_X1 DP_mult_211_U448 ( .A1(DP_mult_211_n599), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n600), .ZN(DP_mult_211_n266) );
  XNOR2_X1 DP_mult_211_U447 ( .A(DP_b_int_2__1_), .B(DP_mult_211_n518), .ZN(
        DP_mult_211_n598) );
  OAI22_X1 DP_mult_211_U446 ( .A1(DP_mult_211_n598), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n599), .ZN(DP_mult_211_n267) );
  XNOR2_X1 DP_mult_211_U445 ( .A(DP_mult_211_n518), .B(DP_b_int_2__0_), .ZN(
        DP_mult_211_n596) );
  OAI22_X1 DP_mult_211_U444 ( .A1(DP_mult_211_n596), .A2(DP_mult_211_n597), 
        .B1(DP_mult_211_n595), .B2(DP_mult_211_n598), .ZN(DP_mult_211_n268) );
  INV_X1 DP_mult_211_U443 ( .A(DP_b_int_2__0_), .ZN(DP_mult_211_n520) );
  NOR2_X1 DP_mult_211_U442 ( .A1(DP_mult_211_n520), .A2(DP_mult_211_n595), 
        .ZN(DP_mult_211_n269) );
  AOI21_X1 DP_mult_211_U441 ( .B1(DP_mult_211_n582), .B2(DP_mult_211_n580), 
        .A(DP_mult_211_n594), .ZN(DP_mult_211_n593) );
  INV_X1 DP_mult_211_U440 ( .A(DP_mult_211_n593), .ZN(DP_mult_211_n270) );
  XNOR2_X1 DP_mult_211_U439 ( .A(DP_b_int_2__9_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n591) );
  OAI22_X1 DP_mult_211_U438 ( .A1(DP_mult_211_n591), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n592), .ZN(DP_mult_211_n271) );
  XNOR2_X1 DP_mult_211_U437 ( .A(DP_b_int_2__8_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n590) );
  OAI22_X1 DP_mult_211_U436 ( .A1(DP_mult_211_n590), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n591), .ZN(DP_mult_211_n272) );
  XNOR2_X1 DP_mult_211_U435 ( .A(DP_b_int_2__7_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n589) );
  OAI22_X1 DP_mult_211_U434 ( .A1(DP_mult_211_n589), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n590), .ZN(DP_mult_211_n273) );
  XNOR2_X1 DP_mult_211_U433 ( .A(DP_b_int_2__6_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n588) );
  OAI22_X1 DP_mult_211_U432 ( .A1(DP_mult_211_n588), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n589), .ZN(DP_mult_211_n274) );
  XNOR2_X1 DP_mult_211_U431 ( .A(DP_b_int_2__5_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n587) );
  OAI22_X1 DP_mult_211_U430 ( .A1(DP_mult_211_n587), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n588), .ZN(DP_mult_211_n275) );
  OAI22_X1 DP_mult_211_U429 ( .A1(DP_mult_211_n586), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n587), .ZN(DP_mult_211_n276) );
  XNOR2_X1 DP_mult_211_U428 ( .A(DP_b_int_2__2_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n584) );
  OAI22_X1 DP_mult_211_U427 ( .A1(DP_mult_211_n584), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n585), .ZN(DP_mult_211_n278) );
  XNOR2_X1 DP_mult_211_U426 ( .A(DP_b_int_2__1_), .B(DP_a_int_1__9_), .ZN(
        DP_mult_211_n583) );
  OAI22_X1 DP_mult_211_U425 ( .A1(DP_mult_211_n583), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n584), .ZN(DP_mult_211_n279) );
  XNOR2_X1 DP_mult_211_U424 ( .A(DP_a_int_1__9_), .B(DP_b_int_2__0_), .ZN(
        DP_mult_211_n581) );
  OAI22_X1 DP_mult_211_U423 ( .A1(DP_mult_211_n581), .A2(DP_mult_211_n582), 
        .B1(DP_mult_211_n580), .B2(DP_mult_211_n583), .ZN(DP_mult_211_n280) );
  NOR2_X1 DP_mult_211_U422 ( .A1(DP_mult_211_n520), .A2(DP_mult_211_n580), 
        .ZN(DP_mult_211_n281) );
  AOI21_X1 DP_mult_211_U421 ( .B1(DP_mult_211_n567), .B2(DP_mult_211_n565), 
        .A(DP_mult_211_n579), .ZN(DP_mult_211_n578) );
  INV_X1 DP_mult_211_U420 ( .A(DP_mult_211_n578), .ZN(DP_mult_211_n282) );
  XNOR2_X1 DP_mult_211_U419 ( .A(DP_b_int_2__9_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n576) );
  OAI22_X1 DP_mult_211_U418 ( .A1(DP_mult_211_n576), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n577), .ZN(DP_mult_211_n283) );
  XNOR2_X1 DP_mult_211_U417 ( .A(DP_b_int_2__8_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n575) );
  OAI22_X1 DP_mult_211_U416 ( .A1(DP_mult_211_n575), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n576), .ZN(DP_mult_211_n284) );
  XNOR2_X1 DP_mult_211_U415 ( .A(DP_b_int_2__7_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n574) );
  OAI22_X1 DP_mult_211_U414 ( .A1(DP_mult_211_n574), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n575), .ZN(DP_mult_211_n285) );
  XNOR2_X1 DP_mult_211_U413 ( .A(DP_b_int_2__6_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n573) );
  OAI22_X1 DP_mult_211_U412 ( .A1(DP_mult_211_n573), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n574), .ZN(DP_mult_211_n286) );
  XNOR2_X1 DP_mult_211_U411 ( .A(DP_b_int_2__5_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n572) );
  OAI22_X1 DP_mult_211_U410 ( .A1(DP_mult_211_n572), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n573), .ZN(DP_mult_211_n287) );
  XNOR2_X1 DP_mult_211_U409 ( .A(DP_b_int_2__4_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n571) );
  OAI22_X1 DP_mult_211_U408 ( .A1(DP_mult_211_n571), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n572), .ZN(DP_mult_211_n288) );
  XNOR2_X1 DP_mult_211_U407 ( .A(DP_b_int_2__3_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n570) );
  OAI22_X1 DP_mult_211_U406 ( .A1(DP_mult_211_n570), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n571), .ZN(DP_mult_211_n289) );
  XNOR2_X1 DP_mult_211_U405 ( .A(DP_b_int_2__2_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n569) );
  OAI22_X1 DP_mult_211_U404 ( .A1(DP_mult_211_n569), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n570), .ZN(DP_mult_211_n290) );
  XNOR2_X1 DP_mult_211_U403 ( .A(DP_b_int_2__1_), .B(DP_a_int_1__7_), .ZN(
        DP_mult_211_n568) );
  OAI22_X1 DP_mult_211_U402 ( .A1(DP_mult_211_n568), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n569), .ZN(DP_mult_211_n291) );
  XNOR2_X1 DP_mult_211_U401 ( .A(DP_a_int_1__7_), .B(DP_b_int_2__0_), .ZN(
        DP_mult_211_n566) );
  OAI22_X1 DP_mult_211_U400 ( .A1(DP_mult_211_n566), .A2(DP_mult_211_n567), 
        .B1(DP_mult_211_n565), .B2(DP_mult_211_n568), .ZN(DP_mult_211_n292) );
  NOR2_X1 DP_mult_211_U399 ( .A1(DP_mult_211_n520), .A2(DP_mult_211_n565), 
        .ZN(DP_mult_211_n293) );
  AOI21_X1 DP_mult_211_U398 ( .B1(DP_mult_211_n552), .B2(DP_mult_211_n550), 
        .A(DP_mult_211_n564), .ZN(DP_mult_211_n563) );
  INV_X1 DP_mult_211_U397 ( .A(DP_mult_211_n563), .ZN(DP_mult_211_n294) );
  XNOR2_X1 DP_mult_211_U396 ( .A(DP_b_int_2__9_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n561) );
  OAI22_X1 DP_mult_211_U395 ( .A1(DP_mult_211_n561), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n562), .ZN(DP_mult_211_n295) );
  OAI22_X1 DP_mult_211_U394 ( .A1(DP_mult_211_n560), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n561), .ZN(DP_mult_211_n296) );
  XNOR2_X1 DP_mult_211_U393 ( .A(DP_b_int_2__6_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n558) );
  OAI22_X1 DP_mult_211_U392 ( .A1(DP_mult_211_n558), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n559), .ZN(DP_mult_211_n298) );
  XNOR2_X1 DP_mult_211_U391 ( .A(DP_b_int_2__5_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n557) );
  OAI22_X1 DP_mult_211_U390 ( .A1(DP_mult_211_n557), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n558), .ZN(DP_mult_211_n299) );
  XNOR2_X1 DP_mult_211_U389 ( .A(DP_b_int_2__4_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n556) );
  OAI22_X1 DP_mult_211_U388 ( .A1(DP_mult_211_n556), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n557), .ZN(DP_mult_211_n300) );
  XNOR2_X1 DP_mult_211_U387 ( .A(DP_b_int_2__3_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n555) );
  OAI22_X1 DP_mult_211_U386 ( .A1(DP_mult_211_n555), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n556), .ZN(DP_mult_211_n301) );
  XNOR2_X1 DP_mult_211_U385 ( .A(DP_b_int_2__2_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n554) );
  OAI22_X1 DP_mult_211_U384 ( .A1(DP_mult_211_n554), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n555), .ZN(DP_mult_211_n302) );
  XNOR2_X1 DP_mult_211_U383 ( .A(DP_b_int_2__1_), .B(DP_a_int_1__5_), .ZN(
        DP_mult_211_n553) );
  OAI22_X1 DP_mult_211_U382 ( .A1(DP_mult_211_n553), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n554), .ZN(DP_mult_211_n303) );
  XNOR2_X1 DP_mult_211_U381 ( .A(DP_a_int_1__5_), .B(DP_b_int_2__0_), .ZN(
        DP_mult_211_n551) );
  OAI22_X1 DP_mult_211_U380 ( .A1(DP_mult_211_n551), .A2(DP_mult_211_n552), 
        .B1(DP_mult_211_n550), .B2(DP_mult_211_n553), .ZN(DP_mult_211_n304) );
  NOR2_X1 DP_mult_211_U379 ( .A1(DP_mult_211_n520), .A2(DP_mult_211_n550), 
        .ZN(DP_mult_211_n305) );
  AOI21_X1 DP_mult_211_U378 ( .B1(DP_mult_211_n537), .B2(DP_mult_211_n535), 
        .A(DP_mult_211_n549), .ZN(DP_mult_211_n548) );
  INV_X1 DP_mult_211_U377 ( .A(DP_mult_211_n548), .ZN(DP_mult_211_n306) );
  XNOR2_X1 DP_mult_211_U376 ( .A(DP_b_int_2__9_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n546) );
  OAI22_X1 DP_mult_211_U375 ( .A1(DP_mult_211_n546), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n547), .ZN(DP_mult_211_n307) );
  XNOR2_X1 DP_mult_211_U374 ( .A(DP_b_int_2__8_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n545) );
  OAI22_X1 DP_mult_211_U373 ( .A1(DP_mult_211_n545), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n546), .ZN(DP_mult_211_n308) );
  XNOR2_X1 DP_mult_211_U372 ( .A(DP_b_int_2__7_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n544) );
  OAI22_X1 DP_mult_211_U371 ( .A1(DP_mult_211_n544), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n545), .ZN(DP_mult_211_n309) );
  XNOR2_X1 DP_mult_211_U370 ( .A(DP_b_int_2__6_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n543) );
  OAI22_X1 DP_mult_211_U369 ( .A1(DP_mult_211_n543), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n544), .ZN(DP_mult_211_n310) );
  XNOR2_X1 DP_mult_211_U368 ( .A(DP_b_int_2__5_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n542) );
  OAI22_X1 DP_mult_211_U367 ( .A1(DP_mult_211_n542), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n543), .ZN(DP_mult_211_n311) );
  XNOR2_X1 DP_mult_211_U366 ( .A(DP_b_int_2__4_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n541) );
  OAI22_X1 DP_mult_211_U365 ( .A1(DP_mult_211_n541), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n542), .ZN(DP_mult_211_n312) );
  XNOR2_X1 DP_mult_211_U364 ( .A(DP_b_int_2__3_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n540) );
  OAI22_X1 DP_mult_211_U363 ( .A1(DP_mult_211_n540), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n541), .ZN(DP_mult_211_n313) );
  XNOR2_X1 DP_mult_211_U362 ( .A(DP_b_int_2__2_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n539) );
  OAI22_X1 DP_mult_211_U361 ( .A1(DP_mult_211_n539), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n540), .ZN(DP_mult_211_n314) );
  XNOR2_X1 DP_mult_211_U360 ( .A(DP_b_int_2__1_), .B(DP_a_int_1__3_), .ZN(
        DP_mult_211_n538) );
  OAI22_X1 DP_mult_211_U359 ( .A1(DP_mult_211_n538), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n539), .ZN(DP_mult_211_n315) );
  XNOR2_X1 DP_mult_211_U358 ( .A(DP_a_int_1__3_), .B(DP_b_int_2__0_), .ZN(
        DP_mult_211_n536) );
  OAI22_X1 DP_mult_211_U357 ( .A1(DP_mult_211_n536), .A2(DP_mult_211_n537), 
        .B1(DP_mult_211_n535), .B2(DP_mult_211_n538), .ZN(DP_mult_211_n316) );
  NOR2_X1 DP_mult_211_U356 ( .A1(DP_mult_211_n520), .A2(DP_mult_211_n535), 
        .ZN(DP_mult_211_n317) );
  XNOR2_X1 DP_mult_211_U355 ( .A(DP_b_int_2__11_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n533) );
  AOI21_X1 DP_mult_211_U354 ( .B1(DP_mult_211_n522), .B2(DP_mult_211_n521), 
        .A(DP_mult_211_n533), .ZN(DP_mult_211_n534) );
  INV_X1 DP_mult_211_U353 ( .A(DP_mult_211_n534), .ZN(DP_mult_211_n318) );
  XNOR2_X1 DP_mult_211_U352 ( .A(DP_b_int_2__10_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n532) );
  OAI22_X1 DP_mult_211_U351 ( .A1(DP_mult_211_n532), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n533), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n319) );
  XNOR2_X1 DP_mult_211_U350 ( .A(DP_b_int_2__9_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n531) );
  OAI22_X1 DP_mult_211_U349 ( .A1(DP_mult_211_n531), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n532), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n320) );
  XNOR2_X1 DP_mult_211_U348 ( .A(DP_b_int_2__8_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n530) );
  OAI22_X1 DP_mult_211_U347 ( .A1(DP_mult_211_n530), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n531), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n321) );
  XNOR2_X1 DP_mult_211_U346 ( .A(DP_b_int_2__7_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n529) );
  OAI22_X1 DP_mult_211_U345 ( .A1(DP_mult_211_n529), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n530), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n322) );
  XNOR2_X1 DP_mult_211_U344 ( .A(DP_b_int_2__6_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n528) );
  OAI22_X1 DP_mult_211_U343 ( .A1(DP_mult_211_n528), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n529), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n323) );
  XNOR2_X1 DP_mult_211_U342 ( .A(DP_b_int_2__5_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n527) );
  OAI22_X1 DP_mult_211_U341 ( .A1(DP_mult_211_n527), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n528), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n324) );
  XNOR2_X1 DP_mult_211_U340 ( .A(DP_b_int_2__4_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n526) );
  OAI22_X1 DP_mult_211_U339 ( .A1(DP_mult_211_n526), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n527), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n325) );
  XNOR2_X1 DP_mult_211_U338 ( .A(DP_b_int_2__3_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n525) );
  OAI22_X1 DP_mult_211_U337 ( .A1(DP_mult_211_n525), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n526), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n326) );
  XNOR2_X1 DP_mult_211_U336 ( .A(DP_b_int_2__2_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n524) );
  OAI22_X1 DP_mult_211_U335 ( .A1(DP_mult_211_n524), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n525), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n327) );
  XNOR2_X1 DP_mult_211_U334 ( .A(DP_b_int_2__1_), .B(DP_a_int_1__1_), .ZN(
        DP_mult_211_n523) );
  OAI22_X1 DP_mult_211_U333 ( .A1(DP_mult_211_n523), .A2(DP_mult_211_n522), 
        .B1(DP_mult_211_n524), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n328) );
  OAI22_X1 DP_mult_211_U332 ( .A1(DP_b_int_2__0_), .A2(DP_mult_211_n522), .B1(
        DP_mult_211_n523), .B2(DP_mult_211_n521), .ZN(DP_mult_211_n329) );
  NOR2_X1 DP_mult_211_U331 ( .A1(DP_mult_211_n520), .A2(DP_mult_211_n521), 
        .ZN(DP_coeff_pipe03[0]) );
  INV_X1 DP_mult_211_U330 ( .A(DP_mult_211_n120), .ZN(DP_N145) );
  INV_X1 DP_mult_211_U329 ( .A(DP_a_int_1__1_), .ZN(DP_mult_211_n513) );
  XOR2_X2 DP_mult_211_U328 ( .A(DP_a_int_1__10_), .B(DP_mult_211_n517), .Z(
        DP_mult_211_n595) );
  XOR2_X2 DP_mult_211_U327 ( .A(DP_a_int_1__8_), .B(DP_mult_211_n516), .Z(
        DP_mult_211_n580) );
  XOR2_X2 DP_mult_211_U326 ( .A(DP_a_int_1__6_), .B(DP_mult_211_n515), .Z(
        DP_mult_211_n565) );
  XOR2_X2 DP_mult_211_U325 ( .A(DP_a_int_1__4_), .B(DP_mult_211_n514), .Z(
        DP_mult_211_n550) );
  XOR2_X2 DP_mult_211_U324 ( .A(DP_a_int_1__2_), .B(DP_mult_211_n513), .Z(
        DP_mult_211_n535) );
  INV_X1 DP_mult_211_U323 ( .A(DP_a_int_1__11_), .ZN(DP_mult_211_n519) );
  INV_X1 DP_mult_211_U322 ( .A(DP_a_int_1__5_), .ZN(DP_mult_211_n515) );
  INV_X1 DP_mult_211_U321 ( .A(DP_a_int_1__3_), .ZN(DP_mult_211_n514) );
  INV_X1 DP_mult_211_U320 ( .A(DP_a_int_1__7_), .ZN(DP_mult_211_n516) );
  INV_X1 DP_mult_211_U319 ( .A(DP_a_int_1__9_), .ZN(DP_mult_211_n517) );
  INV_X1 DP_mult_211_U318 ( .A(DP_coeff_ret0[1]), .ZN(DP_mult_211_n521) );
  INV_X1 DP_mult_211_U317 ( .A(DP_mult_211_n519), .ZN(DP_mult_211_n518) );
  HA_X1 DP_mult_211_U107 ( .A(DP_mult_211_n316), .B(DP_mult_211_n327), .CO(
        DP_mult_211_n250), .S(DP_mult_211_n251) );
  FA_X1 DP_mult_211_U106 ( .A(DP_mult_211_n326), .B(DP_mult_211_n305), .CI(
        DP_mult_211_n315), .CO(DP_mult_211_n248), .S(DP_mult_211_n249) );
  HA_X1 DP_mult_211_U105 ( .A(DP_mult_211_n255), .B(DP_mult_211_n304), .CO(
        DP_mult_211_n246), .S(DP_mult_211_n247) );
  FA_X1 DP_mult_211_U104 ( .A(DP_mult_211_n314), .B(DP_mult_211_n325), .CI(
        DP_mult_211_n247), .CO(DP_mult_211_n244), .S(DP_mult_211_n245) );
  FA_X1 DP_mult_211_U103 ( .A(DP_mult_211_n324), .B(DP_mult_211_n293), .CI(
        DP_mult_211_n313), .CO(DP_mult_211_n242), .S(DP_mult_211_n243) );
  FA_X1 DP_mult_211_U102 ( .A(DP_mult_211_n246), .B(DP_mult_211_n303), .CI(
        DP_mult_211_n243), .CO(DP_mult_211_n240), .S(DP_mult_211_n241) );
  HA_X1 DP_mult_211_U101 ( .A(DP_mult_211_n254), .B(DP_mult_211_n292), .CO(
        DP_mult_211_n238), .S(DP_mult_211_n239) );
  FA_X1 DP_mult_211_U100 ( .A(DP_mult_211_n302), .B(DP_mult_211_n323), .CI(
        DP_mult_211_n312), .CO(DP_mult_211_n236), .S(DP_mult_211_n237) );
  FA_X1 DP_mult_211_U99 ( .A(DP_mult_211_n242), .B(DP_mult_211_n239), .CI(
        DP_mult_211_n237), .CO(DP_mult_211_n234), .S(DP_mult_211_n235) );
  FA_X1 DP_mult_211_U98 ( .A(DP_mult_211_n301), .B(DP_mult_211_n281), .CI(
        DP_mult_211_n322), .CO(DP_mult_211_n232), .S(DP_mult_211_n233) );
  FA_X1 DP_mult_211_U97 ( .A(DP_mult_211_n291), .B(DP_mult_211_n311), .CI(
        DP_mult_211_n238), .CO(DP_mult_211_n230), .S(DP_mult_211_n231) );
  FA_X1 DP_mult_211_U96 ( .A(DP_mult_211_n233), .B(DP_mult_211_n236), .CI(
        DP_mult_211_n231), .CO(DP_mult_211_n228), .S(DP_mult_211_n229) );
  HA_X1 DP_mult_211_U95 ( .A(DP_mult_211_n253), .B(DP_mult_211_n280), .CO(
        DP_mult_211_n226), .S(DP_mult_211_n227) );
  FA_X1 DP_mult_211_U94 ( .A(DP_mult_211_n290), .B(DP_mult_211_n300), .CI(
        DP_mult_211_n310), .CO(DP_mult_211_n224), .S(DP_mult_211_n225) );
  FA_X1 DP_mult_211_U93 ( .A(DP_mult_211_n227), .B(DP_mult_211_n321), .CI(
        DP_mult_211_n232), .CO(DP_mult_211_n222), .S(DP_mult_211_n223) );
  FA_X1 DP_mult_211_U92 ( .A(DP_mult_211_n225), .B(DP_mult_211_n230), .CI(
        DP_mult_211_n223), .CO(DP_mult_211_n220), .S(DP_mult_211_n221) );
  FA_X1 DP_mult_211_U91 ( .A(DP_mult_211_n289), .B(DP_mult_211_n269), .CI(
        DP_mult_211_n320), .CO(DP_mult_211_n218), .S(DP_mult_211_n219) );
  FA_X1 DP_mult_211_U90 ( .A(DP_mult_211_n279), .B(DP_mult_211_n309), .CI(
        DP_mult_211_n299), .CO(DP_mult_211_n216), .S(DP_mult_211_n217) );
  FA_X1 DP_mult_211_U89 ( .A(DP_mult_211_n224), .B(DP_mult_211_n226), .CI(
        DP_mult_211_n219), .CO(DP_mult_211_n214), .S(DP_mult_211_n215) );
  FA_X1 DP_mult_211_U88 ( .A(DP_mult_211_n222), .B(DP_mult_211_n217), .CI(
        DP_mult_211_n215), .CO(DP_mult_211_n212), .S(DP_mult_211_n213) );
  HA_X1 DP_mult_211_U87 ( .A(DP_mult_211_n252), .B(DP_mult_211_n268), .CO(
        DP_mult_211_n210), .S(DP_mult_211_n211) );
  FA_X1 DP_mult_211_U86 ( .A(DP_mult_211_n278), .B(DP_mult_211_n298), .CI(
        DP_mult_211_n319), .CO(DP_mult_211_n208), .S(DP_mult_211_n209) );
  FA_X1 DP_mult_211_U85 ( .A(DP_mult_211_n288), .B(DP_mult_211_n308), .CI(
        DP_mult_211_n211), .CO(DP_mult_211_n206), .S(DP_mult_211_n207) );
  FA_X1 DP_mult_211_U84 ( .A(DP_mult_211_n216), .B(DP_mult_211_n218), .CI(
        DP_mult_211_n209), .CO(DP_mult_211_n204), .S(DP_mult_211_n205) );
  FA_X1 DP_mult_211_U83 ( .A(DP_mult_211_n214), .B(DP_mult_211_n207), .CI(
        DP_mult_211_n205), .CO(DP_mult_211_n202), .S(DP_mult_211_n203) );
  FA_X1 DP_mult_211_U80 ( .A(DP_mult_211_n267), .B(DP_mult_211_n287), .CI(
        DP_mult_211_n318), .CO(DP_mult_211_n198), .S(DP_mult_211_n199) );
  FA_X1 DP_mult_211_U79 ( .A(DP_mult_211_n210), .B(DP_mult_211_n307), .CI(
        DP_mult_211_n201), .CO(DP_mult_211_n196), .S(DP_mult_211_n197) );
  FA_X1 DP_mult_211_U78 ( .A(DP_mult_211_n199), .B(DP_mult_211_n208), .CI(
        DP_mult_211_n206), .CO(DP_mult_211_n194), .S(DP_mult_211_n195) );
  FA_X1 DP_mult_211_U77 ( .A(DP_mult_211_n204), .B(DP_mult_211_n197), .CI(
        DP_mult_211_n195), .CO(DP_mult_211_n192), .S(DP_mult_211_n193) );
  FA_X1 DP_mult_211_U75 ( .A(DP_mult_211_n296), .B(DP_mult_211_n276), .CI(
        DP_mult_211_n191), .CO(DP_mult_211_n188), .S(DP_mult_211_n189) );
  FA_X1 DP_mult_211_U74 ( .A(DP_mult_211_n266), .B(DP_mult_211_n286), .CI(
        DP_mult_211_n200), .CO(DP_mult_211_n186), .S(DP_mult_211_n187) );
  FA_X1 DP_mult_211_U73 ( .A(DP_mult_211_n196), .B(DP_mult_211_n198), .CI(
        DP_mult_211_n189), .CO(DP_mult_211_n184), .S(DP_mult_211_n185) );
  FA_X1 DP_mult_211_U72 ( .A(DP_mult_211_n194), .B(DP_mult_211_n187), .CI(
        DP_mult_211_n185), .CO(DP_mult_211_n182), .S(DP_mult_211_n183) );
  FA_X1 DP_mult_211_U71 ( .A(DP_mult_211_n190), .B(DP_mult_211_n265), .CI(
        DP_mult_211_n306), .CO(DP_mult_211_n180), .S(DP_mult_211_n181) );
  FA_X1 DP_mult_211_U70 ( .A(DP_mult_211_n275), .B(DP_mult_211_n295), .CI(
        DP_mult_211_n285), .CO(DP_mult_211_n178), .S(DP_mult_211_n179) );
  FA_X1 DP_mult_211_U69 ( .A(DP_mult_211_n186), .B(DP_mult_211_n188), .CI(
        DP_mult_211_n179), .CO(DP_mult_211_n176), .S(DP_mult_211_n177) );
  FA_X1 DP_mult_211_U68 ( .A(DP_mult_211_n184), .B(DP_mult_211_n181), .CI(
        DP_mult_211_n177), .CO(DP_mult_211_n174), .S(DP_mult_211_n175) );
  FA_X1 DP_mult_211_U66 ( .A(DP_mult_211_n264), .B(DP_mult_211_n274), .CI(
        DP_mult_211_n173), .CO(DP_mult_211_n170), .S(DP_mult_211_n171) );
  FA_X1 DP_mult_211_U65 ( .A(DP_mult_211_n180), .B(DP_mult_211_n284), .CI(
        DP_mult_211_n178), .CO(DP_mult_211_n168), .S(DP_mult_211_n169) );
  FA_X1 DP_mult_211_U64 ( .A(DP_mult_211_n176), .B(DP_mult_211_n171), .CI(
        DP_mult_211_n169), .CO(DP_mult_211_n166), .S(DP_mult_211_n167) );
  FA_X1 DP_mult_211_U63 ( .A(DP_mult_211_n172), .B(DP_mult_211_n263), .CI(
        DP_mult_211_n294), .CO(DP_mult_211_n164), .S(DP_mult_211_n165) );
  FA_X1 DP_mult_211_U62 ( .A(DP_mult_211_n273), .B(DP_mult_211_n283), .CI(
        DP_mult_211_n170), .CO(DP_mult_211_n162), .S(DP_mult_211_n163) );
  FA_X1 DP_mult_211_U61 ( .A(DP_mult_211_n168), .B(DP_mult_211_n165), .CI(
        DP_mult_211_n163), .CO(DP_mult_211_n160), .S(DP_mult_211_n161) );
  FA_X1 DP_mult_211_U59 ( .A(DP_mult_211_n262), .B(DP_mult_211_n272), .CI(
        DP_mult_211_n159), .CO(DP_mult_211_n156), .S(DP_mult_211_n157) );
  FA_X1 DP_mult_211_U58 ( .A(DP_mult_211_n157), .B(DP_mult_211_n164), .CI(
        DP_mult_211_n162), .CO(DP_mult_211_n154), .S(DP_mult_211_n155) );
  FA_X1 DP_mult_211_U57 ( .A(DP_mult_211_n261), .B(DP_mult_211_n158), .CI(
        DP_mult_211_n282), .CO(DP_mult_211_n152), .S(DP_mult_211_n153) );
  FA_X1 DP_mult_211_U56 ( .A(DP_mult_211_n156), .B(DP_mult_211_n271), .CI(
        DP_mult_211_n153), .CO(DP_mult_211_n150), .S(DP_mult_211_n151) );
  FA_X1 DP_mult_211_U54 ( .A(DP_mult_211_n149), .B(DP_mult_211_n260), .CI(
        DP_mult_211_n152), .CO(DP_mult_211_n146), .S(DP_mult_211_n147) );
  FA_X1 DP_mult_211_U53 ( .A(DP_mult_211_n259), .B(DP_mult_211_n148), .CI(
        DP_mult_211_n270), .CO(DP_mult_211_n144), .S(DP_mult_211_n145) );
  HA_X1 DP_mult_211_U51 ( .A(DP_mult_211_n329), .B(DP_mult_211_n257), .CO(
        DP_mult_211_n141), .S(DP_N123) );
  FA_X1 DP_mult_211_U50 ( .A(DP_mult_211_n328), .B(DP_mult_211_n317), .CI(
        DP_mult_211_n141), .CO(DP_mult_211_n140), .S(DP_N124) );
  FA_X1 DP_mult_211_U49 ( .A(DP_mult_211_n251), .B(DP_mult_211_n256), .CI(
        DP_mult_211_n140), .CO(DP_mult_211_n139), .S(DP_N125) );
  FA_X1 DP_mult_211_U48 ( .A(DP_mult_211_n249), .B(DP_mult_211_n250), .CI(
        DP_mult_211_n139), .CO(DP_mult_211_n138), .S(DP_N126) );
  FA_X1 DP_mult_211_U47 ( .A(DP_mult_211_n245), .B(DP_mult_211_n248), .CI(
        DP_mult_211_n138), .CO(DP_mult_211_n137), .S(DP_N127) );
  FA_X1 DP_mult_211_U46 ( .A(DP_mult_211_n241), .B(DP_mult_211_n244), .CI(
        DP_mult_211_n137), .CO(DP_mult_211_n136), .S(DP_N128) );
  FA_X1 DP_mult_211_U45 ( .A(DP_mult_211_n235), .B(DP_mult_211_n240), .CI(
        DP_mult_211_n136), .CO(DP_mult_211_n135), .S(DP_N129) );
  FA_X1 DP_mult_211_U44 ( .A(DP_mult_211_n229), .B(DP_mult_211_n234), .CI(
        DP_mult_211_n135), .CO(DP_mult_211_n134), .S(DP_N130) );
  FA_X1 DP_mult_211_U43 ( .A(DP_mult_211_n221), .B(DP_mult_211_n228), .CI(
        DP_mult_211_n134), .CO(DP_mult_211_n133), .S(DP_N131) );
  FA_X1 DP_mult_211_U42 ( .A(DP_mult_211_n213), .B(DP_mult_211_n220), .CI(
        DP_mult_211_n133), .CO(DP_mult_211_n132), .S(DP_N132) );
  FA_X1 DP_mult_211_U41 ( .A(DP_mult_211_n203), .B(DP_mult_211_n212), .CI(
        DP_mult_211_n132), .CO(DP_mult_211_n131), .S(DP_N133) );
  FA_X1 DP_mult_211_U40 ( .A(DP_mult_211_n193), .B(DP_mult_211_n202), .CI(
        DP_mult_211_n131), .CO(DP_mult_211_n130), .S(DP_N134) );
  FA_X1 DP_mult_211_U39 ( .A(DP_mult_211_n183), .B(DP_mult_211_n192), .CI(
        DP_mult_211_n130), .CO(DP_mult_211_n129), .S(DP_N135) );
  FA_X1 DP_mult_211_U38 ( .A(DP_mult_211_n175), .B(DP_mult_211_n182), .CI(
        DP_mult_211_n129), .CO(DP_mult_211_n128), .S(DP_N136) );
  FA_X1 DP_mult_211_U37 ( .A(DP_mult_211_n167), .B(DP_mult_211_n174), .CI(
        DP_mult_211_n128), .CO(DP_mult_211_n127), .S(DP_N137) );
  FA_X1 DP_mult_211_U36 ( .A(DP_mult_211_n161), .B(DP_mult_211_n166), .CI(
        DP_mult_211_n127), .CO(DP_mult_211_n126), .S(DP_N138) );
  FA_X1 DP_mult_211_U30 ( .A(DP_mult_211_n160), .B(DP_mult_211_n155), .CI(
        DP_mult_211_n126), .CO(DP_mult_211_n125), .S(DP_N139) );
  FA_X1 DP_mult_211_U20 ( .A(DP_mult_211_n151), .B(DP_mult_211_n154), .CI(
        DP_mult_211_n125), .CO(DP_mult_211_n124), .S(DP_N140) );
  FA_X1 DP_mult_211_U10 ( .A(DP_mult_211_n147), .B(DP_mult_211_n150), .CI(
        DP_mult_211_n124), .CO(DP_mult_211_n123), .S(DP_N141) );
  FA_X1 DP_mult_211_U9 ( .A(DP_mult_211_n146), .B(DP_mult_211_n145), .CI(
        DP_mult_211_n123), .CO(DP_mult_211_n122), .S(DP_N142) );
  FA_X1 DP_mult_211_U8 ( .A(DP_mult_211_n144), .B(DP_mult_211_n143), .CI(
        DP_mult_211_n122), .CO(DP_mult_211_n121), .S(DP_N143) );
  FA_X1 DP_mult_211_U7 ( .A(DP_mult_211_n258), .B(DP_mult_211_n142), .CI(
        DP_mult_211_n121), .CO(DP_mult_211_n120), .S(DP_N144) );
  INV_X1 DP_sub_211_U69 ( .A(DP_N132), .ZN(DP_sub_211_B_not_10_) );
  INV_X1 DP_sub_211_U68 ( .A(DP_N133), .ZN(DP_sub_211_B_not_11_) );
  INV_X1 DP_sub_211_U67 ( .A(DP_N134), .ZN(DP_sub_211_B_not_12_) );
  INV_X1 DP_sub_211_U66 ( .A(DP_N135), .ZN(DP_sub_211_B_not_13_) );
  INV_X1 DP_sub_211_U65 ( .A(DP_N136), .ZN(DP_sub_211_B_not_14_) );
  INV_X1 DP_sub_211_U64 ( .A(DP_N137), .ZN(DP_sub_211_B_not_15_) );
  INV_X1 DP_sub_211_U63 ( .A(DP_N138), .ZN(DP_sub_211_B_not_16_) );
  INV_X1 DP_sub_211_U62 ( .A(DP_N139), .ZN(DP_sub_211_B_not_17_) );
  INV_X1 DP_sub_211_U61 ( .A(DP_N140), .ZN(DP_sub_211_B_not_18_) );
  INV_X1 DP_sub_211_U60 ( .A(DP_N141), .ZN(DP_sub_211_B_not_19_) );
  INV_X1 DP_sub_211_U59 ( .A(DP_N123), .ZN(DP_sub_211_B_not_1_) );
  INV_X1 DP_sub_211_U58 ( .A(DP_N142), .ZN(DP_sub_211_B_not_20_) );
  INV_X1 DP_sub_211_U57 ( .A(DP_N143), .ZN(DP_sub_211_B_not_21_) );
  INV_X1 DP_sub_211_U56 ( .A(DP_N144), .ZN(DP_sub_211_B_not_22_) );
  INV_X1 DP_sub_211_U55 ( .A(DP_N145), .ZN(DP_sub_211_B_not_23_) );
  INV_X1 DP_sub_211_U54 ( .A(DP_N124), .ZN(DP_sub_211_B_not_2_) );
  INV_X1 DP_sub_211_U53 ( .A(DP_N125), .ZN(DP_sub_211_B_not_3_) );
  INV_X1 DP_sub_211_U52 ( .A(DP_N126), .ZN(DP_sub_211_B_not_4_) );
  INV_X1 DP_sub_211_U51 ( .A(DP_N127), .ZN(DP_sub_211_B_not_5_) );
  INV_X1 DP_sub_211_U50 ( .A(DP_N128), .ZN(DP_sub_211_B_not_6_) );
  INV_X1 DP_sub_211_U49 ( .A(DP_N129), .ZN(DP_sub_211_B_not_7_) );
  INV_X1 DP_sub_211_U48 ( .A(DP_N130), .ZN(DP_sub_211_B_not_8_) );
  INV_X1 DP_sub_211_U47 ( .A(DP_N131), .ZN(DP_sub_211_B_not_9_) );
  INV_X1 DP_sub_211_U46 ( .A(DP_coeff_pipe03[0]), .ZN(DP_sub_211_carry_1_) );
  XOR2_X1 DP_sub_211_U45 ( .A(DP_sub_211_B_not_1_), .B(DP_sub_211_carry_1_), 
        .Z(DP_coeff_pipe03[1]) );
  AND2_X1 DP_sub_211_U44 ( .A1(DP_sub_211_carry_1_), .A2(DP_sub_211_B_not_1_), 
        .ZN(DP_sub_211_carry_2_) );
  AND2_X1 DP_sub_211_U43 ( .A1(DP_sub_211_carry_2_), .A2(DP_sub_211_B_not_2_), 
        .ZN(DP_sub_211_carry_3_) );
  XOR2_X1 DP_sub_211_U42 ( .A(DP_sub_211_B_not_3_), .B(DP_sub_211_carry_3_), 
        .Z(DP_coeff_pipe03[3]) );
  AND2_X1 DP_sub_211_U41 ( .A1(DP_sub_211_carry_3_), .A2(DP_sub_211_B_not_3_), 
        .ZN(DP_sub_211_carry_4_) );
  XOR2_X1 DP_sub_211_U40 ( .A(DP_sub_211_B_not_4_), .B(DP_sub_211_carry_4_), 
        .Z(DP_coeff_pipe03[4]) );
  AND2_X1 DP_sub_211_U39 ( .A1(DP_sub_211_carry_4_), .A2(DP_sub_211_B_not_4_), 
        .ZN(DP_sub_211_carry_5_) );
  XOR2_X1 DP_sub_211_U38 ( .A(DP_sub_211_B_not_5_), .B(DP_sub_211_carry_5_), 
        .Z(DP_coeff_pipe03[5]) );
  AND2_X1 DP_sub_211_U37 ( .A1(DP_sub_211_carry_5_), .A2(DP_sub_211_B_not_5_), 
        .ZN(DP_sub_211_carry_6_) );
  XOR2_X1 DP_sub_211_U36 ( .A(DP_sub_211_B_not_6_), .B(DP_sub_211_carry_6_), 
        .Z(DP_coeff_pipe03[6]) );
  AND2_X1 DP_sub_211_U35 ( .A1(DP_sub_211_carry_6_), .A2(DP_sub_211_B_not_6_), 
        .ZN(DP_sub_211_carry_7_) );
  XOR2_X1 DP_sub_211_U34 ( .A(DP_sub_211_B_not_7_), .B(DP_sub_211_carry_7_), 
        .Z(DP_coeff_pipe03[7]) );
  AND2_X1 DP_sub_211_U33 ( .A1(DP_sub_211_carry_7_), .A2(DP_sub_211_B_not_7_), 
        .ZN(DP_sub_211_carry_8_) );
  XOR2_X1 DP_sub_211_U32 ( .A(DP_sub_211_B_not_8_), .B(DP_sub_211_carry_8_), 
        .Z(DP_coeff_pipe03[8]) );
  AND2_X1 DP_sub_211_U31 ( .A1(DP_sub_211_carry_8_), .A2(DP_sub_211_B_not_8_), 
        .ZN(DP_sub_211_carry_9_) );
  XOR2_X1 DP_sub_211_U30 ( .A(DP_sub_211_B_not_9_), .B(DP_sub_211_carry_9_), 
        .Z(DP_coeff_pipe03[9]) );
  AND2_X1 DP_sub_211_U29 ( .A1(DP_sub_211_carry_9_), .A2(DP_sub_211_B_not_9_), 
        .ZN(DP_sub_211_carry_10_) );
  XOR2_X1 DP_sub_211_U28 ( .A(DP_sub_211_B_not_10_), .B(DP_sub_211_carry_10_), 
        .Z(DP_coeff_pipe03[10]) );
  AND2_X1 DP_sub_211_U27 ( .A1(DP_sub_211_carry_10_), .A2(DP_sub_211_B_not_10_), .ZN(DP_sub_211_carry_11_) );
  XOR2_X1 DP_sub_211_U26 ( .A(DP_sub_211_B_not_11_), .B(DP_sub_211_carry_11_), 
        .Z(DP_coeff_pipe03[11]) );
  AND2_X1 DP_sub_211_U25 ( .A1(DP_sub_211_carry_11_), .A2(DP_sub_211_B_not_11_), .ZN(DP_sub_211_carry_12_) );
  XOR2_X1 DP_sub_211_U24 ( .A(DP_sub_211_B_not_12_), .B(DP_sub_211_carry_12_), 
        .Z(DP_coeff_pipe03[12]) );
  AND2_X1 DP_sub_211_U23 ( .A1(DP_sub_211_carry_12_), .A2(DP_sub_211_B_not_12_), .ZN(DP_sub_211_carry_13_) );
  XOR2_X1 DP_sub_211_U22 ( .A(DP_sub_211_B_not_13_), .B(DP_sub_211_carry_13_), 
        .Z(DP_coeff_pipe03[13]) );
  AND2_X1 DP_sub_211_U21 ( .A1(DP_sub_211_carry_13_), .A2(DP_sub_211_B_not_13_), .ZN(DP_sub_211_carry_14_) );
  XOR2_X1 DP_sub_211_U20 ( .A(DP_sub_211_B_not_14_), .B(DP_sub_211_carry_14_), 
        .Z(DP_coeff_pipe03[14]) );
  AND2_X1 DP_sub_211_U19 ( .A1(DP_sub_211_carry_14_), .A2(DP_sub_211_B_not_14_), .ZN(DP_sub_211_carry_15_) );
  XOR2_X1 DP_sub_211_U18 ( .A(DP_sub_211_B_not_15_), .B(DP_sub_211_carry_15_), 
        .Z(DP_coeff_pipe03[15]) );
  AND2_X1 DP_sub_211_U17 ( .A1(DP_sub_211_carry_15_), .A2(DP_sub_211_B_not_15_), .ZN(DP_sub_211_carry_16_) );
  XOR2_X1 DP_sub_211_U16 ( .A(DP_sub_211_B_not_16_), .B(DP_sub_211_carry_16_), 
        .Z(DP_coeff_pipe03[16]) );
  AND2_X1 DP_sub_211_U15 ( .A1(DP_sub_211_carry_16_), .A2(DP_sub_211_B_not_16_), .ZN(DP_sub_211_carry_17_) );
  XOR2_X1 DP_sub_211_U14 ( .A(DP_sub_211_B_not_17_), .B(DP_sub_211_carry_17_), 
        .Z(DP_coeff_pipe03[17]) );
  AND2_X1 DP_sub_211_U13 ( .A1(DP_sub_211_carry_17_), .A2(DP_sub_211_B_not_17_), .ZN(DP_sub_211_carry_18_) );
  XOR2_X1 DP_sub_211_U12 ( .A(DP_sub_211_B_not_18_), .B(DP_sub_211_carry_18_), 
        .Z(DP_coeff_pipe03[18]) );
  AND2_X1 DP_sub_211_U11 ( .A1(DP_sub_211_carry_18_), .A2(DP_sub_211_B_not_18_), .ZN(DP_sub_211_carry_19_) );
  XOR2_X1 DP_sub_211_U10 ( .A(DP_sub_211_B_not_19_), .B(DP_sub_211_carry_19_), 
        .Z(DP_coeff_pipe03[19]) );
  AND2_X1 DP_sub_211_U9 ( .A1(DP_sub_211_carry_19_), .A2(DP_sub_211_B_not_19_), 
        .ZN(DP_sub_211_carry_20_) );
  XOR2_X1 DP_sub_211_U8 ( .A(DP_sub_211_B_not_20_), .B(DP_sub_211_carry_20_), 
        .Z(DP_coeff_pipe03[20]) );
  AND2_X1 DP_sub_211_U7 ( .A1(DP_sub_211_carry_20_), .A2(DP_sub_211_B_not_20_), 
        .ZN(DP_sub_211_carry_21_) );
  XOR2_X1 DP_sub_211_U6 ( .A(DP_sub_211_B_not_21_), .B(DP_sub_211_carry_21_), 
        .Z(DP_coeff_pipe03[21]) );
  AND2_X1 DP_sub_211_U5 ( .A1(DP_sub_211_carry_21_), .A2(DP_sub_211_B_not_21_), 
        .ZN(DP_sub_211_carry_22_) );
  XOR2_X1 DP_sub_211_U4 ( .A(DP_sub_211_B_not_22_), .B(DP_sub_211_carry_22_), 
        .Z(DP_coeff_pipe03[22]) );
  AND2_X1 DP_sub_211_U3 ( .A1(DP_sub_211_carry_22_), .A2(DP_sub_211_B_not_22_), 
        .ZN(DP_sub_211_carry_23_) );
  XOR2_X1 DP_sub_211_U2 ( .A(DP_sub_211_B_not_23_), .B(DP_sub_211_carry_23_), 
        .Z(DP_coeff_pipe03[23]) );
  XOR2_X2 DP_sub_211_U1 ( .A(DP_sub_211_B_not_2_), .B(DP_sub_211_carry_2_), 
        .Z(DP_coeff_pipe03[2]) );
  XOR2_X1 DP_add_1_root_sub_0_root_sub_227_U2 ( .A(DP_ret1[0]), .B(DP_ret0[0]), 
        .Z(DP_w_0_) );
  AND2_X1 DP_add_1_root_sub_0_root_sub_227_U1 ( .A1(DP_ret0[0]), .A2(
        DP_ret1[0]), .ZN(DP_add_1_root_sub_0_root_sub_227_carry_1_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_1 ( .A(DP_ret0[1]), .B(DP_ret1[1]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_1_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_2_), .S(DP_fb_1_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_2 ( .A(DP_ret0[2]), .B(DP_ret1[2]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_2_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_3_), .S(DP_fb_2_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_3 ( .A(DP_ret0[3]), .B(DP_ret1[3]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_3_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_4_), .S(DP_fb_3_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_4 ( .A(DP_ret0[4]), .B(DP_ret1[4]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_4_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_5_), .S(DP_fb_4_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_5 ( .A(DP_ret0[5]), .B(DP_ret1[5]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_5_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_6_), .S(DP_fb_5_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_6 ( .A(DP_ret0[6]), .B(DP_ret1[6]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_6_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_7_), .S(DP_fb_6_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_7 ( .A(DP_ret0[7]), .B(DP_ret1[7]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_7_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_8_), .S(DP_fb_7_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_8 ( .A(DP_ret0[8]), .B(DP_ret1[8]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_8_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_9_), .S(DP_fb_8_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_9 ( .A(DP_ret0[9]), .B(DP_ret1[9]), 
        .CI(DP_add_1_root_sub_0_root_sub_227_carry_9_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_10_), .S(DP_fb_9_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_10 ( .A(DP_ret0[10]), .B(
        DP_ret1[10]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_10_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_11_), .S(DP_fb_10_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_11 ( .A(DP_ret0[11]), .B(
        DP_ret1[11]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_11_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_12_), .S(DP_fb_11_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_12 ( .A(DP_ret0[12]), .B(
        DP_ret1[12]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_12_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_13_), .S(DP_fb_12_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_13 ( .A(DP_ret0[13]), .B(
        DP_ret1[13]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_13_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_14_), .S(DP_fb_13_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_14 ( .A(DP_ret0[14]), .B(
        DP_ret1[14]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_14_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_15_), .S(DP_fb_14_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_15 ( .A(DP_ret0[15]), .B(
        DP_ret1[15]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_15_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_16_), .S(DP_fb_15_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_16 ( .A(DP_ret0[16]), .B(
        DP_ret1[16]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_16_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_17_), .S(DP_fb_16_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_17 ( .A(DP_ret0[17]), .B(
        DP_ret1[17]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_17_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_18_), .S(DP_fb_17_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_18 ( .A(DP_ret0[18]), .B(
        DP_ret1[18]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_18_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_19_), .S(DP_fb_18_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_19 ( .A(DP_ret0[19]), .B(
        DP_ret1[19]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_19_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_20_), .S(DP_fb_19_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_20 ( .A(DP_ret0[20]), .B(
        DP_ret1[20]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_20_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_21_), .S(DP_fb_20_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_21 ( .A(DP_ret0[21]), .B(
        DP_ret1[21]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_21_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_22_), .S(DP_fb_21_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_22 ( .A(DP_ret0[22]), .B(
        DP_ret1[22]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_22_), .CO(
        DP_add_1_root_sub_0_root_sub_227_carry_23_), .S(DP_fb_22_) );
  FA_X1 DP_add_1_root_sub_0_root_sub_227_U1_23 ( .A(DP_ret0[23]), .B(
        DP_ret1[23]), .CI(DP_add_1_root_sub_0_root_sub_227_carry_23_), .S(
        DP_fb_23_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U44 ( .A(DP_fb_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_10_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U43 ( .A(DP_fb_11_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_11_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U42 ( .A(DP_fb_12_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_12_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U41 ( .A(DP_fb_13_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_13_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U40 ( .A(DP_fb_14_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_14_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U39 ( .A(DP_fb_15_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_15_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U38 ( .A(DP_fb_16_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_16_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U37 ( .A(DP_fb_17_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_17_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U36 ( .A(DP_fb_18_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_18_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U35 ( .A(DP_fb_19_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_19_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U34 ( .A(DP_fb_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_1_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U33 ( .A(DP_fb_20_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_20_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U32 ( .A(DP_fb_21_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_21_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U31 ( .A(DP_fb_22_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_22_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U30 ( .A(DP_fb_23_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_23_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U29 ( .A(DP_fb_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_2_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U28 ( .A(DP_fb_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_3_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U27 ( .A(DP_fb_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_4_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U26 ( .A(DP_fb_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_5_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U25 ( .A(DP_fb_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_6_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U24 ( .A(DP_fb_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_7_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U23 ( .A(DP_fb_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_8_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U22 ( .A(DP_fb_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_B_not_9_) );
  INV_X1 DP_sub_0_root_sub_0_root_sub_227_U21 ( .A(DP_w_0_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_1_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U20 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_1_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_1_), .Z(DP_w_1_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U19 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_1_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_1_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_2_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U18 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_2_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_2_), .Z(DP_w_2_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U17 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_2_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_2_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_3_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U16 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_3_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_3_), .Z(DP_w_3_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U15 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_3_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_3_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_4_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U14 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_4_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_4_), .Z(DP_w_4_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U13 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_4_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_4_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_5_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U12 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_5_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_5_), .Z(DP_w_5_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U11 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_5_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_5_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_6_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U10 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_6_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_6_), .Z(DP_w_6_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U9 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_6_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_6_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_7_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U8 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_7_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_7_), .Z(DP_w_7_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U7 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_7_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_7_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_8_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U6 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_8_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_8_), .Z(DP_w_8_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U5 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_8_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_8_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_9_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U4 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_9_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_9_), .Z(DP_w_9_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U3 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_9_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_9_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_10_) );
  XOR2_X1 DP_sub_0_root_sub_0_root_sub_227_U2 ( .A(
        DP_sub_0_root_sub_0_root_sub_227_B_not_10_), .B(
        DP_sub_0_root_sub_0_root_sub_227_carry_10_), .Z(DP_w_10_) );
  AND2_X1 DP_sub_0_root_sub_0_root_sub_227_U1 ( .A1(
        DP_sub_0_root_sub_0_root_sub_227_carry_10_), .A2(
        DP_sub_0_root_sub_0_root_sub_227_B_not_10_), .ZN(
        DP_sub_0_root_sub_0_root_sub_227_carry_11_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_11 ( .A(DP_x_0_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_11_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_11_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_12_), .S(DP_w_11_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_12 ( .A(DP_x_1_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_12_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_12_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_13_), .S(DP_w_12_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_13 ( .A(DP_x_2_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_13_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_13_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_14_), .S(DP_w_13_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_14 ( .A(DP_x_3_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_14_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_14_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_15_), .S(DP_w_14_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_15 ( .A(DP_x_4_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_15_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_15_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_16_), .S(DP_w_15_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_16 ( .A(DP_x_5_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_16_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_16_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_17_), .S(DP_w_16_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_17 ( .A(DP_x_6_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_17_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_17_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_18_), .S(DP_w_17_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_18 ( .A(DP_x_7_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_18_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_18_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_19_), .S(DP_w_18_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_19 ( .A(DP_x_8_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_19_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_19_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_20_), .S(DP_w_19_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_20 ( .A(DP_x_9_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_20_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_20_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_21_), .S(DP_w_20_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_21 ( .A(DP_x_10_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_21_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_21_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_22_), .S(DP_w_21_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_22 ( .A(DP_x_11_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_22_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_22_), .CO(
        DP_sub_0_root_sub_0_root_sub_227_carry_23_), .S(DP_w_22_) );
  FA_X1 DP_sub_0_root_sub_0_root_sub_227_U2_23 ( .A(DP_x_11_), .B(
        DP_sub_0_root_sub_0_root_sub_227_B_not_23_), .CI(
        DP_sub_0_root_sub_0_root_sub_227_carry_23_), .S(DP_w_23_) );
  XNOR2_X1 CU_U4 ( .A(CU_n2), .B(CU_presentState_0_), .ZN(sw_regs_en_int) );
  XOR2_X1 CU_U3 ( .A(vIn), .B(sw_regs_en_int), .Z(CU_nextState_0_) );
  DFFR_X1 CU_presentState_reg_1_ ( .D(sw_regs_en_int), .CK(clk), .RN(rst_n), 
        .Q(delayed_controls_0__1_), .QN(CU_n2) );
  DFFR_X1 CU_presentState_reg_0_ ( .D(CU_nextState_0_), .CK(clk), .RN(rst_n), 
        .Q(CU_presentState_0_) );
  NAND2_X1 reg_delay_0_U5 ( .A1(sw_regs_en_int), .A2(1'b1), .ZN(reg_delay_0_n2) );
  OAI21_X1 reg_delay_0_U4 ( .B1(1'b1), .B2(reg_delay_0_n4), .A(reg_delay_0_n2), 
        .ZN(reg_delay_0_n6) );
  NAND2_X1 reg_delay_0_U3 ( .A1(1'b1), .A2(delayed_controls_0__1_), .ZN(
        reg_delay_0_n1) );
  OAI21_X1 reg_delay_0_U2 ( .B1(1'b1), .B2(reg_delay_0_n3), .A(reg_delay_0_n1), 
        .ZN(reg_delay_0_n5) );
  DFFR_X1 reg_delay_0_Q_reg_0_ ( .D(reg_delay_0_n5), .CK(clk), .RN(rst_n), .Q(
        delayed_controls_1__1_), .QN(reg_delay_0_n3) );
  DFFR_X1 reg_delay_0_Q_reg_1_ ( .D(reg_delay_0_n6), .CK(clk), .RN(rst_n), .Q(
        delayed_controls_1__0_), .QN(reg_delay_0_n4) );
  NAND2_X1 reg_delay_1_U5 ( .A1(delayed_controls_1__0_), .A2(1'b1), .ZN(
        reg_delay_1_n11) );
  OAI21_X1 reg_delay_1_U4 ( .B1(1'b1), .B2(reg_delay_1_n9), .A(reg_delay_1_n11), .ZN(reg_delay_1_n7) );
  NAND2_X1 reg_delay_1_U3 ( .A1(1'b1), .A2(delayed_controls_1__1_), .ZN(
        reg_delay_1_n12) );
  OAI21_X1 reg_delay_1_U2 ( .B1(1'b1), .B2(reg_delay_1_n10), .A(
        reg_delay_1_n12), .ZN(reg_delay_1_n8) );
  DFFR_X1 reg_delay_1_Q_reg_0_ ( .D(reg_delay_1_n8), .CK(clk), .RN(rst_n), .Q(
        vOut), .QN(reg_delay_1_n10) );
  DFFR_X1 reg_delay_1_Q_reg_1_ ( .D(reg_delay_1_n7), .CK(clk), .RN(rst_n), .Q(
        delayed_controls_2__0_), .QN(reg_delay_1_n9) );
endmodule

